module real_jpeg_18963_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_550),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_0),
.B(n_551),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_1),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_1),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_1),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_1),
.B(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_1),
.B(n_242),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_2),
.Y(n_168)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_2),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_2),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_2),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_3),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_3),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_3),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_3),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_3),
.B(n_357),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_3),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_3),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_3),
.B(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_4),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_4),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_4),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_4),
.B(n_300),
.Y(n_299)
);

AND2x4_ASAP7_75t_SL g313 ( 
.A(n_4),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g349 ( 
.A(n_4),
.B(n_242),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_5),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_5),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_5),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_5),
.B(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_5),
.A2(n_11),
.B1(n_286),
.B2(n_291),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_5),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_6),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_7),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_7),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_7),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_7),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_7),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_7),
.B(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_8),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_8),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_8),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_8),
.Y(n_355)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_8),
.Y(n_443)
);

BUFx4f_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_9),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g348 ( 
.A(n_9),
.Y(n_348)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_9),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_10),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_10),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_10),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_10),
.B(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_10),
.B(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_10),
.B(n_311),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_10),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_10),
.B(n_288),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_11),
.B(n_205),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_11),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_11),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_11),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_11),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_11),
.B(n_441),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_11),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_11),
.B(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_12),
.Y(n_170)
);

NAND2x1_ASAP7_75t_L g173 ( 
.A(n_12),
.B(n_101),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_12),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g252 ( 
.A(n_12),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_12),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_12),
.B(n_355),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_12),
.B(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_12),
.B(n_458),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_13),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_13),
.Y(n_148)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_13),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_14),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_14),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_14),
.B(n_389),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_14),
.B(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_14),
.B(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_14),
.B(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_14),
.B(n_498),
.Y(n_497)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_15),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_15),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_15),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_15),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_15),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_17),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

XOR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_537),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_118),
.B(n_536),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2x1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_74),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_24),
.B(n_74),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_54),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_41),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_26),
.B(n_41),
.C(n_54),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.C(n_37),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_27),
.A2(n_32),
.B1(n_47),
.B2(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_SL g540 ( 
.A(n_27),
.B(n_43),
.C(n_49),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_30),
.Y(n_317)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_30),
.Y(n_389)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_31),
.Y(n_176)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_67),
.C(n_71),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_32),
.A2(n_58),
.B1(n_71),
.B2(n_72),
.Y(n_112)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_36),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_49),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_43),
.A2(n_48),
.B1(n_542),
.B2(n_547),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_44),
.Y(n_151)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_45),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_108),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_46),
.B(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.C(n_66),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_55),
.A2(n_56),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_59),
.A2(n_60),
.B1(n_66),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_64),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

XOR2x1_ASAP7_75t_L g111 ( 
.A(n_67),
.B(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_70),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_71),
.A2(n_72),
.B1(n_107),
.B2(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_103),
.C(n_107),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_113),
.C(n_114),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_75),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_102),
.C(n_111),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_76),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_86),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_82),
.C(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.C(n_98),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_87),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_163)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_91),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_92),
.Y(n_255)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_98),
.B(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_102),
.B(n_111),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_103),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_107),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_107),
.B(n_126),
.C(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_113),
.B(n_114),
.Y(n_186)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI21x1_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_275),
.B(n_531),
.Y(n_118)
);

NOR3x1_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_187),
.C(n_269),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_120),
.A2(n_532),
.B(n_535),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_185),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_121),
.B(n_185),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_177),
.C(n_182),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_122),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_162),
.C(n_164),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_124),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_135),
.C(n_149),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_125),
.B(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_131),
.A2(n_132),
.B1(n_167),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_167),
.C(n_169),
.Y(n_166)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_133),
.Y(n_498)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_134),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_135),
.B(n_149),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.C(n_145),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_136),
.B(n_145),
.Y(n_209)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_141),
.B(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_144),
.Y(n_250)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_148),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_153),
.C(n_157),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_161),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_162),
.B(n_164),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_173),
.C(n_174),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_166),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_211),
.C(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_167),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_167),
.A2(n_212),
.B1(n_218),
.B2(n_225),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_168),
.Y(n_452)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_168),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_169),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_169),
.A2(n_215),
.B1(n_299),
.B2(n_343),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_171),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_174),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_173),
.B(n_241),
.C(n_246),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_173),
.B(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_174),
.A2(n_204),
.B1(n_206),
.B2(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_177),
.A2(n_182),
.B1(n_183),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_177),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_181),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_178),
.B(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_180),
.B(n_181),
.Y(n_264)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_259),
.Y(n_187)
);

NOR2xp67_ASAP7_75t_SL g533 ( 
.A(n_188),
.B(n_259),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_219),
.C(n_221),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_189),
.B(n_219),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_207),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_191),
.B(n_194),
.C(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_192),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_204),
.C(n_206),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_195),
.B(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_203),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_203),
.Y(n_238)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_238),
.Y(n_237)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_207),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_214),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_208),
.B(n_210),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_214),
.B(n_327),
.Y(n_326)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_215),
.B(n_296),
.C(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_221),
.B(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_239),
.C(n_256),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_222),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.C(n_237),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_223),
.B(n_226),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_227),
.A2(n_232),
.B1(n_233),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_227),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_229),
.B(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_231),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_232),
.B(n_421),
.C(n_422),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_232),
.A2(n_233),
.B1(n_421),
.B2(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_235),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_236),
.Y(n_353)
);

XNOR2x1_ASAP7_75t_SL g335 ( 
.A(n_237),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_239),
.B(n_256),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_249),
.C(n_251),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_240),
.B(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_246),
.Y(n_283)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_245),
.Y(n_458)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_249),
.A2(n_251),
.B1(n_252),
.B2(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_249),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_251),
.A2(n_252),
.B1(n_401),
.B2(n_402),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_252),
.B(n_396),
.C(n_401),
.Y(n_395)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_263),
.C(n_268),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_270),
.A2(n_533),
.B(n_534),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_SL g534 ( 
.A(n_271),
.B(n_274),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_371),
.B(n_528),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_365),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_330),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_278),
.B(n_330),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_323),
.Y(n_278)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_279),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_304),
.C(n_318),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.C(n_295),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_282),
.B(n_406),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_284),
.A2(n_285),
.B1(n_295),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_285),
.A2(n_387),
.B(n_390),
.Y(n_386)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_295),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_299),
.Y(n_343)
);

BUFx2_ASAP7_75t_SL g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_304),
.A2(n_319),
.B1(n_320),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_312),
.C(n_315),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.C(n_310),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_306),
.A2(n_310),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_306),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_306),
.B(n_436),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_308),
.B(n_383),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_310),
.Y(n_385)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_311),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_312),
.A2(n_313),
.B1(n_315),
.B2(n_361),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_315),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_326),
.B1(n_328),
.B2(n_329),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_326),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_326),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_369),
.C(n_370),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.C(n_337),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_331),
.A2(n_332),
.B1(n_335),
.B2(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_338),
.B(n_375),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_359),
.C(n_362),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_380),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_344),
.C(n_350),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_L g426 ( 
.A(n_341),
.B(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_344),
.B(n_350),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_345),
.B(n_349),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_348),
.Y(n_399)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_348),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.C(n_356),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_351),
.A2(n_354),
.B1(n_417),
.B2(n_418),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_354),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_354),
.A2(n_418),
.B1(n_486),
.B2(n_487),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_354),
.B(n_482),
.C(n_486),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_355),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_356),
.B(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_362),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_365),
.A2(n_529),
.B(n_530),
.Y(n_528)
);

AND2x2_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_368),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_366),
.B(n_368),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_428),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_377),
.C(n_408),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_374),
.B(n_378),
.Y(n_527)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_381),
.C(n_404),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_405),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_386),
.C(n_395),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_386),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_384),
.B(n_437),
.C(n_440),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx12f_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_396),
.B(n_514),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_SL g470 ( 
.A(n_397),
.B(n_400),
.Y(n_470)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_397),
.A2(n_477),
.B1(n_478),
.B2(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_409),
.B(n_411),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.C(n_426),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_412),
.B(n_524),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_414),
.B(n_426),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_419),
.C(n_424),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_415),
.B(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_420),
.B(n_425),
.Y(n_519)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_421),
.Y(n_466)
);

XOR2x1_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.C(n_527),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_431),
.A2(n_522),
.B(n_526),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_508),
.B(n_521),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_473),
.B(n_507),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_461),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_434),
.B(n_461),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_444),
.C(n_453),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_435),
.B(n_503),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_440),
.Y(n_436)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_444),
.A2(n_445),
.B1(n_453),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_451),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_446),
.B(n_451),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_453),
.Y(n_504)
);

AO22x1_ASAP7_75t_SL g453 ( 
.A1(n_454),
.A2(n_457),
.B1(n_459),
.B2(n_460),
.Y(n_453)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_454),
.Y(n_459)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_457),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_457),
.B(n_459),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_497),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_467),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_463),
.B(n_464),
.C(n_467),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

MAJx2_ASAP7_75t_L g516 ( 
.A(n_468),
.B(n_470),
.C(n_471),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_501),
.B(n_506),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_475),
.A2(n_489),
.B(n_500),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_481),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_481),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_478),
.Y(n_495)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_482),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_496),
.B(n_499),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_494),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_494),
.Y(n_499)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_505),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_502),
.B(n_505),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_509),
.B(n_520),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_SL g521 ( 
.A(n_509),
.B(n_520),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_511),
.B1(n_517),
.B2(n_518),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_512),
.A2(n_513),
.B1(n_515),
.B2(n_516),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_516),
.C(n_517),
.Y(n_525)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_525),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_525),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_538),
.B(n_549),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_548),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_548),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_541),
.Y(n_539)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_542),
.Y(n_547)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);


endmodule