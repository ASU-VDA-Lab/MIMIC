module fake_jpeg_6525_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx4_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_14),
.B(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_28),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_17),
.B(n_16),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_8),
.B(n_12),
.C(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_8),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_39),
.B(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_23),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

XNOR2x1_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_24),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_27),
.C(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_48),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_43),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

OAI31xp33_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_45),
.A3(n_31),
.B(n_44),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_11),
.B(n_15),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_51),
.B(n_11),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_15),
.Y(n_55)
);


endmodule