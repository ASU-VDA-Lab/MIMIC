module fake_jpeg_17528_n_312 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_21),
.C(n_19),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_52),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_19),
.B1(n_34),
.B2(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_48),
.B1(n_56),
.B2(n_18),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_30),
.B1(n_19),
.B2(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_23),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_34),
.B1(n_18),
.B2(n_30),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_29),
.B1(n_25),
.B2(n_21),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_17),
.B1(n_18),
.B2(n_35),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_27),
.B(n_20),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_57),
.A2(n_25),
.B(n_29),
.C(n_21),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_24),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_66),
.Y(n_70)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_68),
.B(n_11),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_SL g130 ( 
.A1(n_69),
.A2(n_11),
.B(n_5),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_35),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_21),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_0),
.Y(n_116)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_80),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_49),
.B1(n_63),
.B2(n_45),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_81),
.B1(n_83),
.B2(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_33),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_33),
.B1(n_20),
.B2(n_31),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_86),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_32),
.B1(n_31),
.B2(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_0),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_88),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_47),
.B(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_10),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_89),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_93),
.A2(n_103),
.B1(n_104),
.B2(n_3),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_96),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_58),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_51),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_45),
.A2(n_25),
.B1(n_1),
.B2(n_2),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_45),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_82),
.B1(n_77),
.B2(n_71),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_105),
.B(n_5),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_74),
.A2(n_58),
.B(n_61),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_118),
.B(n_79),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_9),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_6),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_129),
.C(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_117),
.B(n_76),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_0),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_79),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_9),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_127),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_130),
.B1(n_79),
.B2(n_3),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_16),
.C(n_5),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_133),
.B1(n_102),
.B2(n_97),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_123),
.B(n_128),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_150),
.B(n_160),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_123),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_138),
.B(n_139),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_155),
.B1(n_163),
.B2(n_131),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_70),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_149),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_144),
.B(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_85),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_84),
.B(n_92),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_156),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_69),
.C(n_98),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_129),
.C(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_102),
.B1(n_101),
.B2(n_99),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_91),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_104),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_157),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_114),
.A2(n_96),
.B(n_94),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_158),
.A2(n_164),
.B(n_119),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_159),
.B(n_105),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_101),
.A3(n_7),
.B1(n_11),
.B2(n_13),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_163),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_110),
.A2(n_90),
.B1(n_103),
.B2(n_13),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_167),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_R g168 ( 
.A(n_140),
.B(n_128),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_179),
.B(n_186),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_173),
.B(n_180),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_127),
.B(n_128),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_143),
.C(n_145),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_113),
.B1(n_112),
.B2(n_121),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_181),
.B(n_193),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_136),
.A2(n_112),
.B1(n_125),
.B2(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_136),
.A2(n_108),
.B1(n_106),
.B2(n_131),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_108),
.B(n_7),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_189),
.B(n_194),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_6),
.B(n_13),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_90),
.B1(n_14),
.B2(n_15),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_6),
.B1(n_15),
.B2(n_16),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_220),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_201),
.B(n_203),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_141),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_209),
.C(n_210),
.Y(n_227)
);

BUFx4f_ASAP7_75t_SL g207 ( 
.A(n_184),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_217),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_138),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_135),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_139),
.C(n_149),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_172),
.C(n_166),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_155),
.Y(n_216)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_142),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_219),
.A2(n_171),
.B(n_192),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_164),
.B(n_162),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_221),
.A2(n_173),
.B(n_168),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_228),
.A2(n_230),
.B(n_239),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_237),
.C(n_238),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_194),
.B1(n_170),
.B2(n_177),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_243),
.B1(n_232),
.B2(n_234),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_189),
.B1(n_171),
.B2(n_177),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_233),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_205),
.B(n_175),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_240),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_166),
.C(n_179),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_165),
.C(n_191),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_205),
.A2(n_182),
.B(n_164),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_190),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_190),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_200),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_182),
.B1(n_187),
.B2(n_184),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_167),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_248),
.Y(n_262)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_241),
.B(n_214),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_197),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_219),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_253),
.A2(n_254),
.B(n_257),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_159),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_216),
.B1(n_222),
.B2(n_198),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_239),
.B1(n_218),
.B2(n_240),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_148),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_211),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_227),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_264),
.B(n_272),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_266),
.A2(n_271),
.B1(n_213),
.B2(n_260),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_229),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_207),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_259),
.A2(n_221),
.B(n_230),
.Y(n_268)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_212),
.B(n_202),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_270),
.A2(n_252),
.B(n_246),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_213),
.B1(n_215),
.B2(n_208),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_212),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_287),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_277),
.B(n_278),
.Y(n_294)
);

OAI221xp5_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_244),
.B1(n_256),
.B2(n_215),
.C(n_249),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_255),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_207),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_251),
.B(n_249),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_280),
.B(n_285),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_284),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_255),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_207),
.B(n_187),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_291),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_296),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_264),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_271),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_270),
.B(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_298),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_299),
.B(n_301),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_282),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_267),
.C(n_272),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_300),
.A2(n_106),
.A3(n_148),
.B1(n_169),
.B2(n_289),
.C1(n_290),
.C2(n_302),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_306),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_302),
.B(n_169),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

OAI31xp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_304),
.A3(n_307),
.B(n_309),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_311),
.Y(n_312)
);


endmodule