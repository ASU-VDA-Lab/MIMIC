module real_aes_6550_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_0), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g452 ( .A(n_0), .Y(n_452) );
INVx1_ASAP7_75t_L g512 ( .A(n_1), .Y(n_512) );
INVx1_ASAP7_75t_L g268 ( .A(n_2), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_3), .A2(n_38), .B1(n_187), .B2(n_540), .Y(n_539) );
AOI21xp33_ASAP7_75t_L g175 ( .A1(n_4), .A2(n_176), .B(n_177), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_5), .B(n_174), .Y(n_489) );
AND2x6_ASAP7_75t_L g149 ( .A(n_6), .B(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_7), .A2(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g110 ( .A(n_8), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_8), .B(n_39), .Y(n_453) );
INVx1_ASAP7_75t_L g184 ( .A(n_9), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_10), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g146 ( .A(n_11), .Y(n_146) );
INVx1_ASAP7_75t_L g508 ( .A(n_12), .Y(n_508) );
INVx1_ASAP7_75t_L g250 ( .A(n_13), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_14), .B(n_152), .Y(n_546) );
AOI222xp33_ASAP7_75t_SL g457 ( .A1(n_15), .A2(n_458), .B1(n_459), .B2(n_468), .C1(n_755), .C2(n_756), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_16), .B(n_142), .Y(n_517) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_17), .B(n_125), .Y(n_124) );
AO32x2_ASAP7_75t_L g537 ( .A1(n_17), .A2(n_141), .A3(n_174), .B1(n_500), .B2(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_18), .B(n_187), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_19), .B(n_195), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_20), .B(n_142), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_21), .A2(n_50), .B1(n_187), .B2(n_540), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_22), .B(n_176), .Y(n_204) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_23), .A2(n_78), .B1(n_152), .B2(n_187), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_24), .B(n_187), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_25), .B(n_172), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g459 ( .A1(n_26), .A2(n_460), .B1(n_461), .B2(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g467 ( .A(n_26), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_27), .A2(n_248), .B(n_249), .C(n_251), .Y(n_247) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_28), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_29), .B(n_189), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_30), .B(n_182), .Y(n_269) );
INVx1_ASAP7_75t_L g160 ( .A(n_31), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_32), .B(n_189), .Y(n_534) );
INVx2_ASAP7_75t_L g154 ( .A(n_33), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_34), .B(n_187), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_35), .B(n_189), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_36), .A2(n_42), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_36), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_37), .A2(n_149), .B(n_161), .C(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g158 ( .A(n_40), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_41), .B(n_182), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_42), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_43), .B(n_187), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_44), .A2(n_88), .B1(n_212), .B2(n_540), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_45), .B(n_187), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_46), .B(n_187), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g164 ( .A(n_47), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_48), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_49), .B(n_176), .Y(n_238) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_51), .A2(n_60), .B1(n_152), .B2(n_187), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_52), .A2(n_152), .B1(n_155), .B2(n_161), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_53), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_54), .B(n_187), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g265 ( .A(n_55), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_56), .B(n_187), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_57), .A2(n_181), .B(n_183), .C(n_186), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_58), .Y(n_225) );
INVx1_ASAP7_75t_L g178 ( .A(n_59), .Y(n_178) );
INVx1_ASAP7_75t_L g150 ( .A(n_61), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_62), .B(n_187), .Y(n_513) );
INVx1_ASAP7_75t_L g145 ( .A(n_63), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_64), .Y(n_122) );
AO32x2_ASAP7_75t_L g557 ( .A1(n_65), .A2(n_174), .A3(n_230), .B1(n_500), .B2(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g497 ( .A(n_66), .Y(n_497) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_67), .A2(n_128), .B1(n_129), .B2(n_132), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_67), .Y(n_132) );
INVx1_ASAP7_75t_L g529 ( .A(n_68), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_SL g194 ( .A1(n_69), .A2(n_186), .B(n_195), .C(n_196), .Y(n_194) );
INVxp67_ASAP7_75t_L g197 ( .A(n_70), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_71), .B(n_152), .Y(n_530) );
INVx1_ASAP7_75t_L g116 ( .A(n_72), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_73), .A2(n_105), .B1(n_117), .B2(n_760), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_74), .Y(n_169) );
INVx1_ASAP7_75t_L g218 ( .A(n_75), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_76), .A2(n_102), .B1(n_465), .B2(n_466), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_76), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_77), .B(n_455), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_79), .A2(n_149), .B(n_161), .C(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_80), .B(n_540), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_81), .B(n_152), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_82), .B(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_84), .B(n_195), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_85), .B(n_152), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_86), .A2(n_149), .B(n_161), .C(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
OR2x2_ASAP7_75t_L g449 ( .A(n_87), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g471 ( .A(n_87), .B(n_451), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_89), .A2(n_103), .B1(n_152), .B2(n_153), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_90), .B(n_189), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_91), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_92), .A2(n_149), .B(n_161), .C(n_233), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_93), .Y(n_240) );
INVx1_ASAP7_75t_L g193 ( .A(n_94), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g246 ( .A(n_95), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_96), .B(n_208), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_97), .A2(n_462), .B1(n_463), .B2(n_464), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_97), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_98), .B(n_152), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_99), .B(n_174), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_100), .B(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_101), .A2(n_176), .B(n_192), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_102), .Y(n_466) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g760 ( .A(n_107), .Y(n_760) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g754 ( .A(n_113), .B(n_451), .Y(n_754) );
NOR2x2_ASAP7_75t_L g755 ( .A(n_113), .B(n_450), .Y(n_755) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_456), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g759 ( .A(n_122), .Y(n_759) );
OAI21x1_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_446), .B(n_454), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_133), .B2(n_134), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g468 ( .A1(n_133), .A2(n_469), .B1(n_472), .B2(n_752), .Y(n_468) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g756 ( .A1(n_134), .A2(n_469), .B1(n_757), .B2(n_758), .Y(n_756) );
AND3x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_371), .C(n_420), .Y(n_134) );
NOR3xp33_ASAP7_75t_SL g135 ( .A(n_136), .B(n_278), .C(n_316), .Y(n_135) );
OAI222xp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_199), .B1(n_253), .B2(n_259), .C1(n_273), .C2(n_276), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_170), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_138), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_138), .B(n_321), .Y(n_412) );
BUFx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g289 ( .A(n_139), .B(n_190), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_139), .B(n_171), .Y(n_297) );
AND2x2_ASAP7_75t_L g332 ( .A(n_139), .B(n_309), .Y(n_332) );
OR2x2_ASAP7_75t_L g356 ( .A(n_139), .B(n_171), .Y(n_356) );
OR2x2_ASAP7_75t_L g364 ( .A(n_139), .B(n_263), .Y(n_364) );
AND2x2_ASAP7_75t_L g367 ( .A(n_139), .B(n_190), .Y(n_367) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g261 ( .A(n_140), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g275 ( .A(n_140), .B(n_190), .Y(n_275) );
AND2x2_ASAP7_75t_L g325 ( .A(n_140), .B(n_263), .Y(n_325) );
AND2x2_ASAP7_75t_L g338 ( .A(n_140), .B(n_171), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_140), .B(n_424), .Y(n_445) );
AO21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_147), .B(n_168), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_141), .B(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g213 ( .A(n_141), .Y(n_213) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_141), .A2(n_264), .B(n_271), .Y(n_263) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_SL g189 ( .A(n_143), .B(n_144), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
OAI22xp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B1(n_164), .B2(n_165), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_148), .A2(n_178), .B(n_179), .C(n_180), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_148), .A2(n_179), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_148), .A2(n_179), .B(n_246), .C(n_247), .Y(n_245) );
INVx4_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
NAND2x1p5_ASAP7_75t_L g165 ( .A(n_149), .B(n_166), .Y(n_165) );
AND2x4_ASAP7_75t_L g176 ( .A(n_149), .B(n_166), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_149), .A2(n_481), .B(n_484), .Y(n_480) );
BUFx3_ASAP7_75t_L g500 ( .A(n_149), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_149), .A2(n_507), .B(n_511), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_149), .A2(n_528), .B(n_531), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_149), .A2(n_544), .B(n_548), .Y(n_543) );
INVx2_ASAP7_75t_L g270 ( .A(n_152), .Y(n_270) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
INVx1_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g155 ( .A1(n_156), .A2(n_158), .B1(n_159), .B2(n_160), .Y(n_155) );
INVx2_ASAP7_75t_L g159 ( .A(n_156), .Y(n_159) );
INVx4_ASAP7_75t_L g248 ( .A(n_156), .Y(n_248) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g163 ( .A(n_157), .Y(n_163) );
AND2x2_ASAP7_75t_L g166 ( .A(n_157), .B(n_167), .Y(n_166) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
INVx3_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
INVx1_ASAP7_75t_L g195 ( .A(n_157), .Y(n_195) );
INVx5_ASAP7_75t_L g179 ( .A(n_161), .Y(n_179) );
AND2x6_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
BUFx3_ASAP7_75t_L g212 ( .A(n_162), .Y(n_212) );
INVx1_ASAP7_75t_L g540 ( .A(n_162), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_165), .A2(n_218), .B(n_219), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_165), .A2(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g487 ( .A(n_167), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g363 ( .A1(n_170), .A2(n_364), .B(n_365), .C(n_368), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_170), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_170), .B(n_308), .Y(n_430) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_190), .Y(n_170) );
AND2x2_ASAP7_75t_SL g274 ( .A(n_171), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g288 ( .A(n_171), .Y(n_288) );
AND2x2_ASAP7_75t_L g315 ( .A(n_171), .B(n_309), .Y(n_315) );
INVx1_ASAP7_75t_SL g323 ( .A(n_171), .Y(n_323) );
AND2x2_ASAP7_75t_L g346 ( .A(n_171), .B(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g424 ( .A(n_171), .Y(n_424) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_188), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_SL g214 ( .A(n_173), .B(n_215), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_173), .B(n_500), .C(n_519), .Y(n_518) );
AO21x1_ASAP7_75t_L g563 ( .A1(n_173), .A2(n_519), .B(n_564), .Y(n_563) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_174), .A2(n_191), .B(n_198), .Y(n_190) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_174), .A2(n_480), .B(n_489), .Y(n_479) );
BUFx2_ASAP7_75t_L g244 ( .A(n_176), .Y(n_244) );
O2A1O1Ixp5_ASAP7_75t_L g496 ( .A1(n_181), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_181), .A2(n_549), .B(n_550), .Y(n_548) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx4_ASAP7_75t_L g236 ( .A(n_182), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_182), .A2(n_488), .B1(n_520), .B2(n_521), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_182), .A2(n_488), .B1(n_539), .B2(n_541), .Y(n_538) );
OAI22xp5_ASAP7_75t_SL g558 ( .A1(n_182), .A2(n_185), .B1(n_559), .B2(n_560), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_185), .B(n_197), .Y(n_196) );
INVx5_ASAP7_75t_L g208 ( .A(n_185), .Y(n_208) );
O2A1O1Ixp5_ASAP7_75t_SL g528 ( .A1(n_186), .A2(n_208), .B(n_529), .C(n_530), .Y(n_528) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_187), .Y(n_237) );
INVx1_ASAP7_75t_L g226 ( .A(n_189), .Y(n_226) );
INVx2_ASAP7_75t_L g230 ( .A(n_189), .Y(n_230) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_189), .A2(n_243), .B(n_252), .Y(n_242) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_189), .A2(n_527), .B(n_534), .Y(n_526) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_189), .A2(n_543), .B(n_551), .Y(n_542) );
BUFx2_ASAP7_75t_L g260 ( .A(n_190), .Y(n_260) );
INVx1_ASAP7_75t_L g322 ( .A(n_190), .Y(n_322) );
INVx3_ASAP7_75t_L g347 ( .A(n_190), .Y(n_347) );
INVx1_ASAP7_75t_L g547 ( .A(n_195), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_199), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_227), .Y(n_199) );
INVx1_ASAP7_75t_L g343 ( .A(n_200), .Y(n_343) );
OAI32xp33_ASAP7_75t_L g349 ( .A1(n_200), .A2(n_288), .A3(n_350), .B1(n_351), .B2(n_352), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_200), .A2(n_354), .B1(n_357), .B2(n_362), .Y(n_353) );
INVx4_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g291 ( .A(n_201), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g369 ( .A(n_201), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g439 ( .A(n_201), .B(n_385), .Y(n_439) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_216), .Y(n_201) );
AND2x2_ASAP7_75t_L g254 ( .A(n_202), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g284 ( .A(n_202), .Y(n_284) );
INVx1_ASAP7_75t_L g303 ( .A(n_202), .Y(n_303) );
OR2x2_ASAP7_75t_L g311 ( .A(n_202), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g318 ( .A(n_202), .B(n_292), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_202), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g339 ( .A(n_202), .B(n_257), .Y(n_339) );
INVx3_ASAP7_75t_L g361 ( .A(n_202), .Y(n_361) );
AND2x2_ASAP7_75t_L g386 ( .A(n_202), .B(n_258), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_202), .B(n_351), .Y(n_434) );
OR2x6_ASAP7_75t_L g202 ( .A(n_203), .B(n_214), .Y(n_202) );
AOI21xp5_ASAP7_75t_SL g203 ( .A1(n_204), .A2(n_205), .B(n_213), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_209), .B(n_210), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_208), .A2(n_268), .B(n_269), .C(n_270), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_208), .A2(n_482), .B(n_483), .Y(n_481) );
INVx2_ASAP7_75t_L g488 ( .A(n_208), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_208), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_210), .A2(n_221), .B(n_222), .Y(n_220) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g251 ( .A(n_212), .Y(n_251) );
INVx1_ASAP7_75t_L g223 ( .A(n_213), .Y(n_223) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_213), .A2(n_492), .B(n_501), .Y(n_491) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_213), .A2(n_506), .B(n_514), .Y(n_505) );
INVx2_ASAP7_75t_L g258 ( .A(n_216), .Y(n_258) );
AND2x2_ASAP7_75t_L g390 ( .A(n_216), .B(n_228), .Y(n_390) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_223), .B(n_224), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_226), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_226), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g432 ( .A(n_227), .Y(n_432) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_241), .Y(n_227) );
INVx1_ASAP7_75t_L g277 ( .A(n_228), .Y(n_277) );
AND2x2_ASAP7_75t_L g304 ( .A(n_228), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_228), .B(n_258), .Y(n_312) );
AND2x2_ASAP7_75t_L g370 ( .A(n_228), .B(n_293), .Y(n_370) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g256 ( .A(n_229), .Y(n_256) );
AND2x2_ASAP7_75t_L g283 ( .A(n_229), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g292 ( .A(n_229), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_229), .B(n_258), .Y(n_358) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_237), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_241), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g305 ( .A(n_241), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_241), .B(n_258), .Y(n_351) );
AND2x2_ASAP7_75t_L g360 ( .A(n_241), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g385 ( .A(n_241), .Y(n_385) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g257 ( .A(n_242), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g293 ( .A(n_242), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_248), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g510 ( .A(n_248), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_248), .A2(n_532), .B(n_533), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_253), .A2(n_263), .B1(n_422), .B2(n_425), .Y(n_421) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OAI21xp5_ASAP7_75t_SL g444 ( .A1(n_255), .A2(n_366), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_256), .B(n_361), .Y(n_378) );
INVx1_ASAP7_75t_L g403 ( .A(n_256), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_257), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g330 ( .A(n_257), .B(n_283), .Y(n_330) );
INVx2_ASAP7_75t_L g286 ( .A(n_258), .Y(n_286) );
INVx1_ASAP7_75t_L g336 ( .A(n_258), .Y(n_336) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_259), .A2(n_411), .B1(n_428), .B2(n_431), .C(n_433), .Y(n_427) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g298 ( .A(n_260), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_260), .B(n_309), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_261), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g352 ( .A(n_261), .B(n_298), .Y(n_352) );
INVx3_ASAP7_75t_SL g393 ( .A(n_261), .Y(n_393) );
AND2x2_ASAP7_75t_L g337 ( .A(n_262), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g366 ( .A(n_262), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_262), .B(n_275), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_262), .B(n_321), .Y(n_407) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g309 ( .A(n_263), .Y(n_309) );
OAI322xp33_ASAP7_75t_L g404 ( .A1(n_263), .A2(n_335), .A3(n_357), .B1(n_405), .B2(n_407), .C1(n_408), .C2(n_409), .Y(n_404) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_270), .A2(n_508), .B(n_509), .C(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_274), .A2(n_277), .B(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_SL g354 ( .A(n_275), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g376 ( .A(n_275), .B(n_288), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_275), .B(n_315), .Y(n_391) );
INVxp67_ASAP7_75t_L g342 ( .A(n_277), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g348 ( .A1(n_277), .A2(n_349), .B(n_353), .C(n_363), .Y(n_348) );
OAI221xp5_ASAP7_75t_SL g278 ( .A1(n_279), .A2(n_287), .B1(n_290), .B2(n_294), .C(n_299), .Y(n_278) );
INVxp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g302 ( .A(n_286), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g419 ( .A(n_286), .Y(n_419) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_287), .A2(n_436), .B1(n_441), .B2(n_442), .C(n_444), .Y(n_435) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_288), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g335 ( .A(n_288), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_288), .B(n_366), .Y(n_373) );
AND2x2_ASAP7_75t_L g415 ( .A(n_288), .B(n_393), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_289), .B(n_314), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_289), .A2(n_301), .B1(n_411), .B2(n_412), .Y(n_410) );
OR2x2_ASAP7_75t_L g441 ( .A(n_289), .B(n_309), .Y(n_441) );
CKINVDCx16_ASAP7_75t_R g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g418 ( .A(n_292), .Y(n_418) );
AND2x2_ASAP7_75t_L g443 ( .A(n_292), .B(n_386), .Y(n_443) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_SL g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g307 ( .A(n_297), .B(n_308), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_306), .B1(n_310), .B2(n_313), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g374 ( .A(n_302), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_302), .B(n_342), .Y(n_409) );
AOI322xp5_ASAP7_75t_L g333 ( .A1(n_304), .A2(n_334), .A3(n_336), .B1(n_337), .B2(n_339), .C1(n_340), .C2(n_344), .Y(n_333) );
INVxp67_ASAP7_75t_L g327 ( .A(n_305), .Y(n_327) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_307), .A2(n_312), .B1(n_329), .B2(n_331), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_308), .B(n_321), .Y(n_408) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_309), .B(n_347), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_309), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g405 ( .A(n_311), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND3xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_333), .C(n_348), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_324), .B2(n_326), .C(n_328), .Y(n_317) );
AND2x2_ASAP7_75t_L g324 ( .A(n_320), .B(n_325), .Y(n_324) );
INVx3_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g334 ( .A(n_325), .B(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_327), .Y(n_406) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_332), .B(n_346), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_335), .B(n_393), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_336), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g411 ( .A(n_339), .Y(n_411) );
AND2x2_ASAP7_75t_L g426 ( .A(n_339), .B(n_403), .Y(n_426) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g420 ( .A1(n_350), .A2(n_421), .B(n_427), .C(n_435), .Y(n_420) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g389 ( .A(n_360), .B(n_390), .Y(n_389) );
NAND2x1_ASAP7_75t_SL g431 ( .A(n_361), .B(n_432), .Y(n_431) );
CKINVDCx16_ASAP7_75t_R g401 ( .A(n_364), .Y(n_401) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g396 ( .A(n_370), .Y(n_396) );
AND2x2_ASAP7_75t_L g400 ( .A(n_370), .B(n_386), .Y(n_400) );
NOR5xp2_ASAP7_75t_L g371 ( .A(n_372), .B(n_387), .C(n_404), .D(n_410), .E(n_413), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B1(n_375), .B2(n_377), .C(n_379), .Y(n_372) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_376), .B(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g402 ( .A(n_386), .B(n_403), .Y(n_402) );
OAI221xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_391), .B1(n_392), .B2(n_394), .C(n_397), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g440 ( .A(n_400), .Y(n_440) );
AOI211xp5_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_416), .B(n_418), .C(n_419), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
CKINVDCx14_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g455 ( .A(n_449), .Y(n_455) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_454), .B(n_457), .C(n_759), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
CKINVDCx14_ASAP7_75t_R g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g757 ( .A(n_472), .Y(n_757) );
NAND2x1p5_ASAP7_75t_L g472 ( .A(n_473), .B(n_676), .Y(n_472) );
AND2x2_ASAP7_75t_SL g473 ( .A(n_474), .B(n_634), .Y(n_473) );
NOR4xp25_ASAP7_75t_L g474 ( .A(n_475), .B(n_574), .C(n_610), .D(n_624), .Y(n_474) );
OAI221xp5_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_522), .B1(n_552), .B2(n_561), .C(n_565), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_476), .B(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_502), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_490), .Y(n_478) );
AND2x2_ASAP7_75t_L g571 ( .A(n_479), .B(n_491), .Y(n_571) );
INVx3_ASAP7_75t_L g579 ( .A(n_479), .Y(n_579) );
AND2x2_ASAP7_75t_L g633 ( .A(n_479), .B(n_505), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_479), .B(n_504), .Y(n_669) );
AND2x2_ASAP7_75t_L g727 ( .A(n_479), .B(n_589), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_488), .Y(n_484) );
INVx2_ASAP7_75t_L g498 ( .A(n_487), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_488), .A2(n_498), .B(n_512), .C(n_513), .Y(n_511) );
AND2x2_ASAP7_75t_L g562 ( .A(n_490), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g576 ( .A(n_490), .B(n_505), .Y(n_576) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_491), .B(n_505), .Y(n_591) );
AND2x2_ASAP7_75t_L g603 ( .A(n_491), .B(n_579), .Y(n_603) );
OR2x2_ASAP7_75t_L g605 ( .A(n_491), .B(n_563), .Y(n_605) );
AND2x2_ASAP7_75t_L g640 ( .A(n_491), .B(n_563), .Y(n_640) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_491), .Y(n_685) );
INVx1_ASAP7_75t_L g693 ( .A(n_491), .Y(n_693) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_496), .B(n_500), .Y(n_492) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_502), .A2(n_611), .B1(n_615), .B2(n_619), .C(n_620), .Y(n_610) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g570 ( .A(n_503), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_515), .Y(n_503) );
INVx2_ASAP7_75t_L g569 ( .A(n_504), .Y(n_569) );
AND2x2_ASAP7_75t_L g622 ( .A(n_504), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g641 ( .A(n_504), .B(n_579), .Y(n_641) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g704 ( .A(n_505), .B(n_579), .Y(n_704) );
AND2x2_ASAP7_75t_L g626 ( .A(n_515), .B(n_571), .Y(n_626) );
OAI322xp33_ASAP7_75t_L g694 ( .A1(n_515), .A2(n_650), .A3(n_695), .B1(n_697), .B2(n_700), .C1(n_702), .C2(n_706), .Y(n_694) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NOR2x1_ASAP7_75t_L g577 ( .A(n_516), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g590 ( .A(n_516), .Y(n_590) );
AND2x2_ASAP7_75t_L g699 ( .A(n_516), .B(n_579), .Y(n_699) );
AND2x2_ASAP7_75t_L g731 ( .A(n_516), .B(n_603), .Y(n_731) );
OR2x2_ASAP7_75t_L g734 ( .A(n_516), .B(n_735), .Y(n_734) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
INVx1_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_535), .Y(n_523) );
INVx1_ASAP7_75t_L g747 ( .A(n_524), .Y(n_747) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g554 ( .A(n_525), .B(n_542), .Y(n_554) );
INVx2_ASAP7_75t_L g587 ( .A(n_525), .Y(n_587) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g609 ( .A(n_526), .Y(n_609) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_526), .Y(n_617) );
OR2x2_ASAP7_75t_L g741 ( .A(n_526), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g566 ( .A(n_535), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g606 ( .A(n_535), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g658 ( .A(n_535), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_542), .Y(n_535) );
AND2x2_ASAP7_75t_L g555 ( .A(n_536), .B(n_556), .Y(n_555) );
NOR2xp67_ASAP7_75t_L g613 ( .A(n_536), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g667 ( .A(n_536), .B(n_557), .Y(n_667) );
OR2x2_ASAP7_75t_L g675 ( .A(n_536), .B(n_609), .Y(n_675) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_L g584 ( .A(n_537), .Y(n_584) );
AND2x2_ASAP7_75t_L g594 ( .A(n_537), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g618 ( .A(n_537), .B(n_542), .Y(n_618) );
AND2x2_ASAP7_75t_L g682 ( .A(n_537), .B(n_557), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_542), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_542), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g595 ( .A(n_542), .Y(n_595) );
INVx1_ASAP7_75t_L g600 ( .A(n_542), .Y(n_600) );
AND2x2_ASAP7_75t_L g612 ( .A(n_542), .B(n_613), .Y(n_612) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_542), .Y(n_690) );
INVx1_ASAP7_75t_L g742 ( .A(n_542), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B(n_547), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_555), .Y(n_552) );
AND2x2_ASAP7_75t_L g719 ( .A(n_553), .B(n_628), .Y(n_719) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g646 ( .A(n_555), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g745 ( .A(n_555), .B(n_680), .Y(n_745) );
INVx1_ASAP7_75t_L g567 ( .A(n_556), .Y(n_567) );
AND2x2_ASAP7_75t_L g593 ( .A(n_556), .B(n_587), .Y(n_593) );
BUFx2_ASAP7_75t_L g652 ( .A(n_556), .Y(n_652) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_557), .Y(n_573) );
INVx1_ASAP7_75t_L g583 ( .A(n_557), .Y(n_583) );
NOR2xp67_ASAP7_75t_L g721 ( .A(n_561), .B(n_568), .Y(n_721) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AOI32xp33_ASAP7_75t_L g565 ( .A1(n_562), .A2(n_566), .A3(n_568), .B1(n_570), .B2(n_572), .Y(n_565) );
AND2x2_ASAP7_75t_L g705 ( .A(n_562), .B(n_578), .Y(n_705) );
AND2x2_ASAP7_75t_L g743 ( .A(n_562), .B(n_641), .Y(n_743) );
INVx1_ASAP7_75t_L g623 ( .A(n_563), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_567), .B(n_629), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_568), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_568), .B(n_571), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_568), .B(n_640), .Y(n_722) );
OR2x2_ASAP7_75t_L g736 ( .A(n_568), .B(n_605), .Y(n_736) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g663 ( .A(n_569), .B(n_571), .Y(n_663) );
OR2x2_ASAP7_75t_L g672 ( .A(n_569), .B(n_659), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_571), .B(n_622), .Y(n_644) );
INVx2_ASAP7_75t_L g659 ( .A(n_573), .Y(n_659) );
OR2x2_ASAP7_75t_L g674 ( .A(n_573), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g689 ( .A(n_573), .B(n_690), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_573), .A2(n_666), .B(n_747), .C(n_748), .Y(n_746) );
OAI321xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_580), .A3(n_585), .B1(n_588), .B2(n_592), .C(n_596), .Y(n_574) );
INVx1_ASAP7_75t_L g687 ( .A(n_575), .Y(n_687) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g698 ( .A(n_576), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g650 ( .A(n_578), .Y(n_650) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_579), .B(n_693), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_580), .A2(n_718), .B1(n_720), .B2(n_722), .C(n_723), .Y(n_717) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
AND2x2_ASAP7_75t_L g655 ( .A(n_582), .B(n_629), .Y(n_655) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_583), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g628 ( .A(n_584), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_585), .A2(n_626), .B(n_671), .C(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g637 ( .A(n_587), .B(n_594), .Y(n_637) );
BUFx2_ASAP7_75t_L g647 ( .A(n_587), .Y(n_647) );
INVx1_ASAP7_75t_L g662 ( .A(n_587), .Y(n_662) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
OR2x2_ASAP7_75t_L g668 ( .A(n_590), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g751 ( .A(n_590), .Y(n_751) );
INVx1_ASAP7_75t_L g744 ( .A(n_591), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g597 ( .A(n_593), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g701 ( .A(n_593), .B(n_618), .Y(n_701) );
INVx1_ASAP7_75t_L g630 ( .A(n_594), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_601), .B1(n_604), .B2(n_606), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_598), .B(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g666 ( .A(n_599), .B(n_667), .Y(n_666) );
BUFx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_600), .B(n_609), .Y(n_629) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g621 ( .A(n_603), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g631 ( .A(n_605), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_608), .A2(n_726), .B1(n_728), .B2(n_729), .C(n_730), .Y(n_725) );
INVx1_ASAP7_75t_L g614 ( .A(n_609), .Y(n_614) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_609), .Y(n_680) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_612), .B(n_731), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_613), .A2(n_618), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_616), .B(n_626), .Y(n_723) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g692 ( .A(n_617), .Y(n_692) );
AND2x2_ASAP7_75t_L g651 ( .A(n_618), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g740 ( .A(n_618), .Y(n_740) );
INVx1_ASAP7_75t_L g656 ( .A(n_621), .Y(n_656) );
INVx1_ASAP7_75t_L g711 ( .A(n_622), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B1(n_630), .B2(n_631), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_628), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g696 ( .A(n_629), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_629), .B(n_667), .Y(n_733) );
OR2x2_ASAP7_75t_L g706 ( .A(n_630), .B(n_659), .Y(n_706) );
INVx1_ASAP7_75t_L g645 ( .A(n_631), .Y(n_645) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_633), .B(n_684), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_653), .C(n_664), .Y(n_634) );
OAI211xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B(n_642), .C(n_648), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_637), .A2(n_708), .B1(n_712), .B2(n_715), .C(n_717), .Y(n_707) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g649 ( .A(n_640), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g703 ( .A(n_640), .B(n_704), .Y(n_703) );
OAI211xp5_ASAP7_75t_L g688 ( .A1(n_641), .A2(n_689), .B(n_691), .C(n_693), .Y(n_688) );
INVx2_ASAP7_75t_L g735 ( .A(n_641), .Y(n_735) );
OAI21xp5_ASAP7_75t_SL g642 ( .A1(n_643), .A2(n_645), .B(n_646), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g714 ( .A(n_647), .B(n_667), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_656), .B(n_657), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_660), .B(n_663), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_658), .B(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_663), .B(n_750), .Y(n_749) );
OAI21xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B(n_670), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g691 ( .A(n_667), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND4x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_707), .C(n_724), .D(n_746), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_694), .Y(n_677) );
OAI211xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_683), .B(n_686), .C(n_688), .Y(n_678) );
OR2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_682), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_693), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g728 ( .A(n_703), .Y(n_728) );
INVx2_ASAP7_75t_SL g716 ( .A(n_704), .Y(n_716) );
OR2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g729 ( .A(n_714), .Y(n_729) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_SL g724 ( .A(n_725), .B(n_732), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
OAI221xp5_ASAP7_75t_SL g732 ( .A1(n_733), .A2(n_734), .B1(n_736), .B2(n_737), .C(n_738), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g758 ( .A(n_753), .Y(n_758) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
endmodule