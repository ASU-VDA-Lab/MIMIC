module fake_ibex_931_n_135 (n_21, n_36, n_14, n_25, n_12, n_13, n_29, n_43, n_5, n_20, n_2, n_9, n_42, n_8, n_37, n_40, n_7, n_28, n_32, n_17, n_10, n_24, n_11, n_18, n_31, n_3, n_1, n_26, n_4, n_35, n_16, n_19, n_44, n_45, n_6, n_27, n_33, n_34, n_39, n_41, n_0, n_23, n_22, n_30, n_38, n_15, n_135);

input n_21;
input n_36;
input n_14;
input n_25;
input n_12;
input n_13;
input n_29;
input n_43;
input n_5;
input n_20;
input n_2;
input n_9;
input n_42;
input n_8;
input n_37;
input n_40;
input n_7;
input n_28;
input n_32;
input n_17;
input n_10;
input n_24;
input n_11;
input n_18;
input n_31;
input n_3;
input n_1;
input n_26;
input n_4;
input n_35;
input n_16;
input n_19;
input n_44;
input n_45;
input n_6;
input n_27;
input n_33;
input n_34;
input n_39;
input n_41;
input n_0;
input n_23;
input n_22;
input n_30;
input n_38;
input n_15;

output n_135;



endmodule