module fake_ariane_1005_n_1779 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1779);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1779;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_37),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_46),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_60),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_15),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_28),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_4),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_17),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_126),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_89),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_12),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_36),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_59),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_106),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_78),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_50),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_46),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_30),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_57),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_8),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_49),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_27),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_114),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_131),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_43),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_29),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_27),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_58),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_32),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_141),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_30),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_61),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_75),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_98),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_37),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_4),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_47),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_67),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_87),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_20),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_51),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_97),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_96),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_133),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_15),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_12),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_77),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_123),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_5),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_41),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_113),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_149),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_116),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_51),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_88),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_44),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_136),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_18),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_1),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_151),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_130),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_99),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_108),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_72),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_16),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_54),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_16),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_148),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_23),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_41),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_156),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_32),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_146),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_39),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_118),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_93),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_52),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_13),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_92),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_25),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_8),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_117),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_22),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_52),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_34),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_45),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_48),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_48),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_56),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_103),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_44),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_56),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_54),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_102),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_143),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_9),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_128),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_110),
.Y(n_271)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_105),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_155),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_63),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_21),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_5),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_104),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_94),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_24),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_64),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_39),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_0),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_120),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_65),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_100),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_74),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_83),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_45),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_157),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_139),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_66),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_14),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_62),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_21),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_43),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_50),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_14),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_38),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_47),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_18),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_17),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_26),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_145),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_152),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_6),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_33),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_31),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_31),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_135),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_26),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_112),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_42),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_2),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_245),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_226),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_245),
.Y(n_318)
);

NOR2xp67_ASAP7_75t_L g319 ( 
.A(n_192),
.B(n_0),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_279),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_286),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_199),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_260),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_216),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_245),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_194),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_245),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_245),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_198),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_257),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_211),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_213),
.B(n_1),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_312),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_257),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_159),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_215),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_201),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_178),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_192),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_160),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_221),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_269),
.B(n_2),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_229),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_178),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_269),
.B(n_3),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_232),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_161),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_260),
.B(n_3),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_162),
.B(n_6),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_178),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_163),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_238),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_239),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_240),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_243),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_257),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_257),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_168),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_247),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_168),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_272),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_272),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_272),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_251),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_289),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_289),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_302),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_278),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_302),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_303),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_164),
.B(n_7),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_278),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_253),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_303),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_173),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_173),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_278),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_296),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_176),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_199),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_297),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_176),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_212),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_298),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_299),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_165),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_316),
.B(n_175),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_316),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_322),
.B(n_244),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_325),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_322),
.B(n_380),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_325),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_326),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_328),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_381),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_323),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_244),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_330),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_330),
.B(n_179),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_336),
.B(n_202),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_349),
.A2(n_260),
.B1(n_210),
.B2(n_166),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_327),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_182),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_384),
.B(n_186),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_362),
.A2(n_237),
.B(n_212),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_362),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_SL g420 ( 
.A(n_353),
.B(n_166),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_334),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_188),
.Y(n_422)
);

AND3x2_ASAP7_75t_L g423 ( 
.A(n_353),
.B(n_174),
.C(n_237),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_197),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_202),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_338),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_343),
.A2(n_315),
.B1(n_314),
.B2(n_258),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_317),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_340),
.B(n_214),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_319),
.B(n_241),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_361),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_345),
.B(n_220),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_363),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_365),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_344),
.B(n_241),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_370),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_335),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_341),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_346),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_371),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_348),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_372),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

OA21x2_ASAP7_75t_L g454 ( 
.A1(n_374),
.A2(n_224),
.B(n_223),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_352),
.B(n_185),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_375),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_356),
.B(n_233),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_339),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_379),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_234),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_351),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_393),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_411),
.B(n_357),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_393),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_420),
.A2(n_354),
.B1(n_376),
.B2(n_347),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_448),
.B(n_358),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_448),
.B(n_359),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_434),
.B(n_360),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_407),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_SL g474 ( 
.A(n_448),
.B(n_355),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_432),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_393),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_448),
.B(n_364),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_397),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_397),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_448),
.B(n_369),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_399),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_434),
.B(n_209),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_432),
.Y(n_484)
);

OAI22xp33_ASAP7_75t_L g485 ( 
.A1(n_429),
.A2(n_389),
.B1(n_386),
.B2(n_378),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_397),
.Y(n_488)
);

INVxp33_ASAP7_75t_L g489 ( 
.A(n_446),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_420),
.A2(n_390),
.B1(n_383),
.B2(n_350),
.Y(n_490)
);

AND2x2_ASAP7_75t_SL g491 ( 
.A(n_444),
.B(n_187),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_401),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_401),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_414),
.B(n_385),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_398),
.B(n_189),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_446),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_444),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_401),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_412),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_412),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_412),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_414),
.B(n_431),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_407),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_431),
.B(n_342),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_444),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_404),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_424),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_L g514 ( 
.A(n_395),
.B(n_204),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_451),
.B(n_320),
.Y(n_515)
);

BUFx4f_ASAP7_75t_L g516 ( 
.A(n_454),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_434),
.B(n_169),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_407),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_423),
.B(n_193),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_424),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_424),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_440),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_434),
.B(n_394),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_404),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_440),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_459),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_404),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_421),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_451),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_451),
.B(n_167),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_430),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_415),
.B(n_196),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_430),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_434),
.B(n_366),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_441),
.A2(n_264),
.B1(n_315),
.B2(n_314),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_399),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_399),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_421),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_L g542 ( 
.A(n_395),
.B(n_204),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_434),
.B(n_236),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_430),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_435),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_413),
.A2(n_280),
.B1(n_265),
.B2(n_283),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_413),
.B(n_172),
.C(n_171),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_394),
.B(n_248),
.Y(n_548)
);

AND2x2_ASAP7_75t_SL g549 ( 
.A(n_405),
.B(n_203),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_395),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_394),
.B(n_271),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_400),
.B(n_167),
.Y(n_552)
);

OR2x6_ASAP7_75t_L g553 ( 
.A(n_455),
.B(n_205),
.Y(n_553)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_429),
.Y(n_554)
);

NAND2x1p5_ASAP7_75t_L g555 ( 
.A(n_454),
.B(n_418),
.Y(n_555)
);

OAI22xp33_ASAP7_75t_SL g556 ( 
.A1(n_441),
.A2(n_462),
.B1(n_458),
.B2(n_437),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_396),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_396),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_400),
.B(n_367),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_427),
.B(n_209),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_396),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_441),
.B(n_170),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_441),
.A2(n_171),
.B1(n_310),
.B2(n_172),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_415),
.B(n_206),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_436),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_441),
.B(n_170),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_402),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_402),
.B(n_406),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_436),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_436),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_423),
.B(n_217),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_402),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_436),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_406),
.B(n_368),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_441),
.B(n_180),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_406),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_403),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_416),
.B(n_180),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_416),
.B(n_373),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_455),
.A2(n_231),
.B1(n_242),
.B2(n_222),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_427),
.B(n_209),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_452),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_405),
.B(n_459),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_440),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_403),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_403),
.Y(n_586)
);

NOR3xp33_ASAP7_75t_L g587 ( 
.A(n_462),
.B(n_275),
.C(n_290),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_416),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_403),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_403),
.B(n_377),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_409),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_426),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_409),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_455),
.A2(n_308),
.B1(n_227),
.B2(n_250),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_409),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_409),
.B(n_427),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_427),
.B(n_181),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_426),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_435),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_409),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_440),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_427),
.B(n_181),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_427),
.B(n_190),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_415),
.B(n_256),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_455),
.B(n_190),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_408),
.B(n_191),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_440),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_408),
.B(n_392),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_SL g609 ( 
.A(n_408),
.B(n_382),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_455),
.B(n_209),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_454),
.Y(n_611)
);

INVxp33_ASAP7_75t_L g612 ( 
.A(n_437),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_455),
.A2(n_337),
.B1(n_331),
.B2(n_324),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_592),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_592),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_491),
.A2(n_410),
.B1(n_392),
.B2(n_458),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_473),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_612),
.B(n_410),
.Y(n_618)
);

AOI22x1_ASAP7_75t_L g619 ( 
.A1(n_577),
.A2(n_438),
.B1(n_460),
.B2(n_443),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_472),
.B(n_204),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_556),
.B(n_449),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_598),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_464),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_491),
.B(n_438),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_598),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_482),
.B(n_449),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_466),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_482),
.B(n_449),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_553),
.B(n_452),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_482),
.B(n_449),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_608),
.B(n_438),
.Y(n_631)
);

OAI221xp5_ASAP7_75t_L g632 ( 
.A1(n_467),
.A2(n_546),
.B1(n_594),
.B2(n_580),
.C(n_547),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_466),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_463),
.B(n_321),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_499),
.B(n_417),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_473),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_487),
.B(n_449),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_511),
.B(n_443),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_468),
.B(n_443),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_470),
.Y(n_641)
);

OAI22x1_ASAP7_75t_SL g642 ( 
.A1(n_475),
.A2(n_276),
.B1(n_275),
.B2(n_184),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_506),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_470),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_476),
.Y(n_645)
);

O2A1O1Ixp5_ASAP7_75t_L g646 ( 
.A1(n_596),
.A2(n_595),
.B(n_487),
.C(n_519),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_512),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_487),
.B(n_595),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_481),
.B(n_445),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_509),
.Y(n_650)
);

A2O1A1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_554),
.A2(n_460),
.B(n_445),
.C(n_457),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_465),
.B(n_417),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_512),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_530),
.B(n_489),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_521),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_574),
.B(n_422),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_530),
.B(n_422),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_476),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_579),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_595),
.B(n_449),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_516),
.B(n_449),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_516),
.B(n_449),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_520),
.A2(n_454),
.B1(n_445),
.B2(n_460),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_524),
.B(n_425),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_525),
.B(n_425),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_528),
.B(n_439),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_516),
.B(n_450),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_521),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_498),
.B(n_439),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_522),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_498),
.B(n_439),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_559),
.B(n_177),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_498),
.B(n_439),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_506),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_480),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_548),
.B(n_442),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_480),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_532),
.B(n_450),
.Y(n_678)
);

NOR3xp33_ASAP7_75t_L g679 ( 
.A(n_485),
.B(n_261),
.C(n_309),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_609),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_532),
.B(n_450),
.Y(n_681)
);

NOR2xp67_ASAP7_75t_SL g682 ( 
.A(n_469),
.B(n_177),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_553),
.B(n_442),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_522),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_486),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_590),
.B(n_183),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_551),
.B(n_442),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_532),
.B(n_450),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_472),
.B(n_204),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_533),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_606),
.B(n_442),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_472),
.B(n_204),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_513),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_486),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_533),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_535),
.Y(n_696)
);

INVxp67_ASAP7_75t_SL g697 ( 
.A(n_513),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_610),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_472),
.B(n_204),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_475),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_539),
.B(n_450),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_505),
.B(n_183),
.Y(n_702)
);

AND2x4_ASAP7_75t_SL g703 ( 
.A(n_553),
.B(n_447),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_471),
.B(n_184),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_520),
.A2(n_454),
.B1(n_453),
.B2(n_461),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_550),
.A2(n_457),
.B(n_456),
.C(n_447),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_518),
.B(n_447),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_610),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_543),
.B(n_447),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_582),
.B(n_456),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_539),
.B(n_456),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_553),
.A2(n_282),
.B1(n_254),
.B2(n_277),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_488),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_539),
.B(n_456),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_513),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_540),
.B(n_457),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_535),
.Y(n_717)
);

AND2x6_ASAP7_75t_L g718 ( 
.A(n_550),
.B(n_209),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_540),
.B(n_477),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_540),
.B(n_457),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_536),
.B(n_254),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_508),
.B(n_450),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_552),
.B(n_450),
.Y(n_723)
);

O2A1O1Ixp5_ASAP7_75t_L g724 ( 
.A1(n_519),
.A2(n_433),
.B(n_428),
.C(n_246),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_544),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_488),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_492),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_531),
.B(n_258),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_492),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_544),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_490),
.A2(n_282),
.B1(n_290),
.B2(n_277),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_502),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_611),
.B(n_450),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_578),
.B(n_453),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_507),
.B(n_276),
.C(n_266),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_611),
.B(n_453),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_519),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_557),
.A2(n_572),
.B(n_588),
.C(n_558),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_557),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_558),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_611),
.B(n_453),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_534),
.B(n_453),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_534),
.B(n_564),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_502),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_520),
.A2(n_454),
.B1(n_461),
.B2(n_453),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_561),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_503),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_503),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_564),
.B(n_453),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_610),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_561),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_610),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_567),
.Y(n_753)
);

AOI221xp5_ASAP7_75t_L g754 ( 
.A1(n_538),
.A2(n_262),
.B1(n_266),
.B2(n_259),
.C(n_264),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_567),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_478),
.B(n_259),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_517),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_571),
.B(n_453),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_517),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_604),
.B(n_461),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_572),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_583),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_604),
.B(n_461),
.Y(n_763)
);

INVx5_ASAP7_75t_L g764 ( 
.A(n_472),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_529),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_529),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_494),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_555),
.A2(n_418),
.B(n_433),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_610),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_576),
.B(n_461),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_576),
.Y(n_771)
);

AO22x2_ASAP7_75t_L g772 ( 
.A1(n_571),
.A2(n_428),
.B1(n_235),
.B2(n_281),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_588),
.Y(n_773)
);

INVx8_ASAP7_75t_L g774 ( 
.A(n_483),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_577),
.B(n_461),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_494),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_585),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_585),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_586),
.B(n_461),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_586),
.B(n_461),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_589),
.B(n_191),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_496),
.B(n_562),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_589),
.B(n_255),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_537),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_591),
.B(n_255),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_591),
.B(n_593),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_648),
.A2(n_568),
.B(n_593),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_614),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_656),
.A2(n_652),
.B1(n_659),
.B2(n_649),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_648),
.A2(n_600),
.B(n_493),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_637),
.Y(n_791)
);

AOI33xp33_ASAP7_75t_L g792 ( 
.A1(n_754),
.A2(n_497),
.A3(n_571),
.B1(n_495),
.B2(n_493),
.B3(n_500),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_664),
.B(n_479),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_623),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_637),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_615),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_622),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_629),
.B(n_497),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_768),
.A2(n_555),
.B(n_600),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_654),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_635),
.B(n_549),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_733),
.A2(n_504),
.B(n_479),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_629),
.B(n_484),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_733),
.A2(n_504),
.B(n_500),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_616),
.B(n_495),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_774),
.B(n_583),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_640),
.A2(n_602),
.B1(n_605),
.B2(n_484),
.Y(n_807)
);

NOR2x1_ASAP7_75t_L g808 ( 
.A(n_657),
.B(n_515),
.Y(n_808)
);

O2A1O1Ixp5_ASAP7_75t_L g809 ( 
.A1(n_686),
.A2(n_603),
.B(n_597),
.C(n_575),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_629),
.B(n_566),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_618),
.B(n_501),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_736),
.A2(n_501),
.B(n_514),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_647),
.A2(n_601),
.B1(n_563),
.B2(n_555),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_736),
.A2(n_542),
.B(n_514),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_625),
.B(n_537),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_634),
.B(n_549),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_653),
.B(n_541),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_655),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_624),
.B(n_474),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_741),
.A2(n_542),
.B(n_601),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_636),
.B(n_650),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_741),
.A2(n_601),
.B(n_494),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_668),
.B(n_541),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_670),
.B(n_565),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_700),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_646),
.A2(n_565),
.B(n_569),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_684),
.B(n_569),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_624),
.B(n_474),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_690),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_724),
.A2(n_570),
.B(n_573),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_743),
.B(n_527),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_695),
.A2(n_587),
.B1(n_607),
.B2(n_494),
.Y(n_832)
);

AOI33xp33_ASAP7_75t_L g833 ( 
.A1(n_731),
.A2(n_310),
.A3(n_262),
.B1(n_573),
.B2(n_570),
.B3(n_300),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_661),
.A2(n_584),
.B(n_494),
.Y(n_834)
);

AOI21x1_ASAP7_75t_L g835 ( 
.A1(n_661),
.A2(n_418),
.B(n_419),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_762),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_696),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_717),
.B(n_510),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_672),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_662),
.A2(n_510),
.B(n_607),
.Y(n_840)
);

INVx4_ASAP7_75t_L g841 ( 
.A(n_774),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_662),
.A2(n_667),
.B(n_628),
.Y(n_842)
);

O2A1O1Ixp5_ASAP7_75t_L g843 ( 
.A1(n_682),
.A2(n_249),
.B(n_263),
.C(n_267),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_758),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_706),
.A2(n_545),
.B(n_599),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_667),
.A2(n_510),
.B(n_607),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_725),
.A2(n_523),
.B1(n_607),
.B2(n_510),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_721),
.B(n_527),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_706),
.A2(n_545),
.B(n_599),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_683),
.B(n_510),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_627),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_730),
.A2(n_740),
.B1(n_746),
.B2(n_739),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_680),
.B(n_613),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_712),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_637),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_751),
.B(n_523),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_704),
.A2(n_523),
.B(n_607),
.C(n_526),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_633),
.Y(n_858)
);

AOI21x1_ASAP7_75t_L g859 ( 
.A1(n_626),
.A2(n_419),
.B(n_292),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_782),
.B(n_523),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_641),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_683),
.B(n_523),
.Y(n_862)
);

AOI33xp33_ASAP7_75t_L g863 ( 
.A1(n_639),
.A2(n_755),
.A3(n_753),
.B1(n_761),
.B2(n_773),
.B3(n_771),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_756),
.A2(n_632),
.B(n_728),
.C(n_738),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_738),
.A2(n_526),
.B(n_584),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_651),
.A2(n_526),
.B(n_584),
.C(n_311),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_758),
.B(n_483),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_626),
.A2(n_584),
.B(n_526),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_639),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_666),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_786),
.A2(n_599),
.B(n_545),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_683),
.B(n_669),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_631),
.B(n_526),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_641),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_628),
.A2(n_584),
.B(n_545),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_651),
.A2(n_288),
.B(n_285),
.C(n_268),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_786),
.A2(n_545),
.B(n_599),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_758),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_676),
.B(n_483),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_774),
.Y(n_880)
);

A2O1A1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_702),
.A2(n_273),
.B(n_306),
.C(n_304),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_644),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_630),
.A2(n_599),
.B(n_581),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_687),
.B(n_483),
.Y(n_884)
);

OA21x2_ASAP7_75t_L g885 ( 
.A1(n_621),
.A2(n_419),
.B(n_270),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_671),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_722),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_679),
.A2(n_301),
.B(n_307),
.C(n_274),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_665),
.B(n_483),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_673),
.B(n_483),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_691),
.B(n_560),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_630),
.A2(n_274),
.B(n_270),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_637),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_707),
.B(n_560),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_638),
.A2(n_581),
.B(n_560),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_643),
.Y(n_896)
);

AOI21x1_ASAP7_75t_L g897 ( 
.A1(n_638),
.A2(n_419),
.B(n_581),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_703),
.A2(n_284),
.B(n_287),
.C(n_291),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_660),
.A2(n_284),
.B(n_287),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_660),
.A2(n_581),
.B(n_560),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_703),
.A2(n_581),
.B1(n_560),
.B2(n_610),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_709),
.B(n_560),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_734),
.A2(n_291),
.B(n_293),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_775),
.A2(n_780),
.B(n_779),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_643),
.B(n_293),
.Y(n_905)
);

NOR2x1_ASAP7_75t_L g906 ( 
.A(n_735),
.B(n_435),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_678),
.A2(n_581),
.B(n_313),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_619),
.A2(n_204),
.B(n_435),
.Y(n_908)
);

OR2x2_ASAP7_75t_SL g909 ( 
.A(n_642),
.B(n_228),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_723),
.A2(n_313),
.B(n_225),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_719),
.B(n_195),
.Y(n_911)
);

BUFx4f_ASAP7_75t_L g912 ( 
.A(n_774),
.Y(n_912)
);

AO21x1_ASAP7_75t_L g913 ( 
.A1(n_621),
.A2(n_204),
.B(n_435),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_742),
.A2(n_7),
.B(n_10),
.C(n_11),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_674),
.A2(n_200),
.B1(n_305),
.B2(n_295),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_711),
.A2(n_219),
.B(n_252),
.Y(n_916)
);

O2A1O1Ixp5_ASAP7_75t_L g917 ( 
.A1(n_749),
.A2(n_435),
.B(n_11),
.C(n_13),
.Y(n_917)
);

BUFx4f_ASAP7_75t_L g918 ( 
.A(n_643),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_772),
.B(n_435),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_714),
.A2(n_230),
.B(n_218),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_772),
.B(n_435),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_760),
.B(n_208),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_643),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_772),
.A2(n_663),
.B1(n_705),
.B2(n_745),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_644),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_763),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_778),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_777),
.B(n_207),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_678),
.A2(n_228),
.B(n_73),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_777),
.B(n_693),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_710),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_716),
.A2(n_228),
.B(n_71),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_674),
.A2(n_228),
.B1(n_19),
.B2(n_20),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_720),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_698),
.B(n_10),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_781),
.A2(n_19),
.B(n_22),
.C(n_23),
.Y(n_936)
);

INVx4_ASAP7_75t_L g937 ( 
.A(n_764),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_617),
.B(n_228),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_617),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_617),
.A2(n_29),
.B1(n_33),
.B2(n_35),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_770),
.A2(n_35),
.B(n_36),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_693),
.B(n_38),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_693),
.B(n_737),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_681),
.A2(n_40),
.B(n_42),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_737),
.B(n_40),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_697),
.A2(n_90),
.B(n_154),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_767),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_767),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_698),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_949)
);

NOR2x1p5_ASAP7_75t_SL g950 ( 
.A(n_645),
.B(n_85),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_777),
.B(n_53),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_715),
.B(n_737),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_776),
.A2(n_91),
.B(n_68),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_767),
.Y(n_954)
);

NAND2xp33_ASAP7_75t_L g955 ( 
.A(n_767),
.B(n_55),
.Y(n_955)
);

O2A1O1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_783),
.A2(n_785),
.B(n_681),
.C(n_688),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_645),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_688),
.A2(n_69),
.B(n_70),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_764),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_701),
.A2(n_76),
.B(n_79),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_715),
.B(n_80),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_701),
.A2(n_81),
.B(n_82),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_708),
.B(n_84),
.Y(n_963)
);

AOI21x1_ASAP7_75t_L g964 ( 
.A1(n_658),
.A2(n_784),
.B(n_766),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_658),
.B(n_95),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_784),
.A2(n_101),
.B(n_109),
.C(n_111),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_675),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_675),
.A2(n_732),
.B(n_766),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_677),
.A2(n_115),
.B(n_119),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_764),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_677),
.B(n_122),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_769),
.Y(n_972)
);

NOR2x1_ASAP7_75t_L g973 ( 
.A(n_685),
.B(n_132),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_764),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_789),
.A2(n_764),
.B1(n_765),
.B2(n_727),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_839),
.B(n_727),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_848),
.A2(n_699),
.B(n_692),
.C(n_620),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_798),
.B(n_825),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_816),
.B(n_726),
.Y(n_979)
);

BUFx4f_ASAP7_75t_L g980 ( 
.A(n_806),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_805),
.A2(n_699),
.B(n_692),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_870),
.B(n_793),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_793),
.A2(n_689),
.B(n_620),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_836),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_811),
.B(n_732),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_835),
.A2(n_729),
.B(n_765),
.Y(n_986)
);

NAND2xp33_ASAP7_75t_SL g987 ( 
.A(n_798),
.B(n_769),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_854),
.A2(n_752),
.B1(n_750),
.B2(n_708),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_918),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_806),
.B(n_752),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_912),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_873),
.A2(n_689),
.B(n_759),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_909),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_864),
.A2(n_729),
.B(n_757),
.C(n_685),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_869),
.B(n_744),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_821),
.B(n_750),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_800),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_873),
.A2(n_726),
.B(n_757),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_801),
.B(n_759),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_794),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_805),
.A2(n_748),
.B1(n_747),
.B2(n_694),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_807),
.A2(n_881),
.B(n_888),
.C(n_831),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_806),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_886),
.B(n_748),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_867),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_809),
.A2(n_694),
.B(n_713),
.C(n_744),
.Y(n_1006)
);

INVx3_ASAP7_75t_SL g1007 ( 
.A(n_803),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_811),
.B(n_713),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_931),
.B(n_747),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_860),
.A2(n_718),
.B(n_144),
.C(n_158),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_814),
.A2(n_718),
.B(n_904),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_819),
.B(n_718),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_867),
.B(n_718),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_788),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_792),
.A2(n_718),
.B(n_863),
.C(n_942),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_904),
.A2(n_718),
.B(n_799),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_818),
.A2(n_829),
.B1(n_837),
.B2(n_924),
.Y(n_1017)
);

CKINVDCx10_ASAP7_75t_R g1018 ( 
.A(n_808),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_955),
.A2(n_936),
.B(n_828),
.C(n_914),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_865),
.A2(n_964),
.B(n_847),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_842),
.A2(n_787),
.B(n_834),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_840),
.A2(n_846),
.B(n_956),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_SL g1023 ( 
.A(n_898),
.B(n_944),
.C(n_941),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_878),
.B(n_810),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_810),
.B(n_844),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_796),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_797),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_926),
.B(n_872),
.Y(n_1028)
);

O2A1O1Ixp5_ASAP7_75t_L g1029 ( 
.A1(n_857),
.A2(n_865),
.B(n_832),
.C(n_905),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_853),
.B(n_935),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_852),
.A2(n_945),
.B1(n_815),
.B2(n_887),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_876),
.A2(n_929),
.B(n_961),
.C(n_911),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_812),
.A2(n_822),
.B(n_820),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_812),
.A2(n_802),
.B(n_826),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_890),
.A2(n_927),
.B1(n_874),
.B2(n_851),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_918),
.Y(n_1036)
);

AOI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_890),
.A2(n_862),
.B1(n_850),
.B2(n_935),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_934),
.B(n_967),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_833),
.B(n_919),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_951),
.A2(n_944),
.B(n_941),
.C(n_813),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_815),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_947),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_868),
.A2(n_804),
.B(n_790),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_951),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_915),
.A2(n_889),
.B1(n_963),
.B2(n_933),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_817),
.B(n_823),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_SL g1047 ( 
.A(n_912),
.B(n_841),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_841),
.B(n_880),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_804),
.A2(n_856),
.B(n_838),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_889),
.A2(n_866),
.B(n_843),
.C(n_943),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_817),
.B(n_823),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_939),
.B(n_940),
.C(n_949),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_974),
.B(n_795),
.Y(n_1053)
);

O2A1O1Ixp5_ASAP7_75t_L g1054 ( 
.A1(n_938),
.A2(n_849),
.B(n_845),
.C(n_830),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_824),
.B(n_827),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_922),
.A2(n_952),
.B(n_928),
.C(n_930),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_791),
.B(n_893),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_974),
.B(n_795),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_838),
.A2(n_856),
.B(n_824),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_921),
.B(n_858),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_827),
.B(n_861),
.Y(n_1061)
);

BUFx8_ASAP7_75t_L g1062 ( 
.A(n_795),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_922),
.A2(n_928),
.B(n_930),
.C(n_917),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_875),
.A2(n_891),
.B(n_871),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_906),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_882),
.B(n_957),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_880),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_SL g1068 ( 
.A1(n_963),
.A2(n_907),
.B1(n_972),
.B2(n_960),
.Y(n_1068)
);

BUFx4f_ASAP7_75t_L g1069 ( 
.A(n_855),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_947),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_925),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_791),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_903),
.A2(n_962),
.B(n_891),
.C(n_910),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_855),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_877),
.A2(n_968),
.B(n_894),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_SL g1076 ( 
.A(n_937),
.B(n_970),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_908),
.A2(n_971),
.B(n_965),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_947),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_894),
.A2(n_902),
.B(n_971),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_902),
.A2(n_879),
.B(n_884),
.C(n_966),
.Y(n_1080)
);

OAI22x1_ASAP7_75t_L g1081 ( 
.A1(n_901),
.A2(n_923),
.B1(n_885),
.B2(n_959),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_879),
.B(n_884),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_948),
.A2(n_954),
.B1(n_895),
.B2(n_900),
.Y(n_1083)
);

BUFx4f_ASAP7_75t_L g1084 ( 
.A(n_855),
.Y(n_1084)
);

OAI22x1_ASAP7_75t_L g1085 ( 
.A1(n_923),
.A2(n_885),
.B1(n_973),
.B2(n_897),
.Y(n_1085)
);

INVx8_ASAP7_75t_L g1086 ( 
.A(n_974),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_896),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_896),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_948),
.B(n_954),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_948),
.Y(n_1090)
);

OA21x2_ASAP7_75t_L g1091 ( 
.A1(n_913),
.A2(n_965),
.B(n_932),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_883),
.A2(n_920),
.B(n_916),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_SL g1093 ( 
.A(n_937),
.B(n_970),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_950),
.Y(n_1094)
);

AND2x2_ASAP7_75t_SL g1095 ( 
.A(n_946),
.B(n_953),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_859),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_892),
.B(n_899),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_958),
.A2(n_864),
.B(n_656),
.C(n_652),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_969),
.B(n_789),
.Y(n_1099)
);

AOI21x1_ASAP7_75t_L g1100 ( 
.A1(n_865),
.A2(n_964),
.B(n_835),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_L g1101 ( 
.A(n_848),
.B(n_672),
.C(n_789),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_788),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_789),
.B(n_499),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_801),
.B(n_816),
.Y(n_1104)
);

AOI21x1_ASAP7_75t_L g1105 ( 
.A1(n_865),
.A2(n_964),
.B(n_835),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_789),
.B(n_656),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_789),
.A2(n_839),
.B(n_659),
.C(n_672),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_912),
.B(n_918),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_789),
.A2(n_864),
.B1(n_616),
.B2(n_656),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_R g1110 ( 
.A(n_825),
.B(n_475),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_789),
.A2(n_864),
.B1(n_616),
.B2(n_656),
.Y(n_1111)
);

CKINVDCx14_ASAP7_75t_R g1112 ( 
.A(n_836),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_835),
.A2(n_865),
.B(n_908),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_SL g1114 ( 
.A1(n_789),
.A2(n_864),
.B(n_839),
.C(n_793),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_788),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_789),
.B(n_652),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_793),
.A2(n_789),
.B(n_873),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_801),
.B(n_816),
.Y(n_1118)
);

OR2x2_ASAP7_75t_L g1119 ( 
.A(n_1104),
.B(n_1118),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1120)
);

NOR2x1_ASAP7_75t_L g1121 ( 
.A(n_1036),
.B(n_1074),
.Y(n_1121)
);

AOI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1109),
.A2(n_1111),
.B1(n_1116),
.B2(n_1101),
.C(n_1107),
.Y(n_1122)
);

AND2x6_ASAP7_75t_L g1123 ( 
.A(n_990),
.B(n_989),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1000),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1032),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1103),
.A2(n_1117),
.B(n_976),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_1099),
.A2(n_982),
.B(n_1015),
.C(n_1031),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1014),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1099),
.A2(n_1095),
.B(n_1114),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1085),
.A2(n_1079),
.A3(n_1080),
.B(n_1094),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_982),
.A2(n_1031),
.B1(n_1045),
.B2(n_1068),
.Y(n_1131)
);

INVx5_ASAP7_75t_L g1132 ( 
.A(n_989),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1100),
.A2(n_1105),
.B(n_1113),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1062),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1062),
.Y(n_1135)
);

BUFx4f_ASAP7_75t_L g1136 ( 
.A(n_989),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1051),
.A2(n_1055),
.B1(n_984),
.B2(n_1046),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_1016),
.A2(n_1096),
.A3(n_1001),
.B(n_975),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1026),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_997),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1027),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1054),
.A2(n_1063),
.B(n_1050),
.Y(n_1142)
);

AO32x2_ASAP7_75t_L g1143 ( 
.A1(n_1017),
.A2(n_975),
.A3(n_1001),
.B1(n_1083),
.B2(n_1003),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1002),
.A2(n_1052),
.B(n_1019),
.C(n_1040),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_SL g1145 ( 
.A1(n_1051),
.A2(n_1055),
.B(n_1044),
.C(n_977),
.Y(n_1145)
);

OA21x2_ASAP7_75t_L g1146 ( 
.A1(n_1022),
.A2(n_1077),
.B(n_1021),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1059),
.A2(n_983),
.B(n_1011),
.Y(n_1147)
);

BUFx2_ASAP7_75t_R g1148 ( 
.A(n_1007),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1023),
.A2(n_1056),
.B(n_978),
.C(n_1029),
.Y(n_1149)
);

OAI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1024),
.A2(n_979),
.B1(n_1017),
.B2(n_1037),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_999),
.A2(n_1073),
.B(n_1012),
.C(n_1041),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_1033),
.A2(n_1034),
.B(n_1043),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1061),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_SL g1154 ( 
.A1(n_1010),
.A2(n_1053),
.B(n_1058),
.C(n_1067),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1030),
.B(n_1038),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1049),
.A2(n_1082),
.B(n_992),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1005),
.B(n_1025),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1064),
.A2(n_1092),
.B(n_985),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_981),
.A2(n_1081),
.A3(n_1075),
.B(n_994),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_1004),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_1039),
.A2(n_1006),
.B(n_985),
.C(n_988),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1008),
.A2(n_1082),
.B(n_1083),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1025),
.B(n_1028),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_1036),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1102),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_1110),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1115),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_SL g1168 ( 
.A1(n_1048),
.A2(n_1061),
.B(n_1009),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1069),
.Y(n_1169)
);

OA21x2_ASAP7_75t_L g1170 ( 
.A1(n_1020),
.A2(n_986),
.B(n_998),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1091),
.A2(n_1093),
.B(n_1076),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1018),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1091),
.A2(n_1076),
.B(n_1047),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1071),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1047),
.A2(n_1048),
.B(n_995),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1097),
.A2(n_996),
.B(n_1060),
.Y(n_1176)
);

NOR3xp33_ASAP7_75t_L g1177 ( 
.A(n_1112),
.B(n_1057),
.C(n_991),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1024),
.B(n_1088),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1048),
.A2(n_987),
.B(n_1067),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1065),
.A2(n_1089),
.B(n_1035),
.C(n_1072),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1066),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1087),
.Y(n_1182)
);

BUFx2_ASAP7_75t_R g1183 ( 
.A(n_1013),
.Y(n_1183)
);

NOR2xp67_ASAP7_75t_L g1184 ( 
.A(n_1042),
.B(n_1078),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1042),
.B(n_1078),
.C(n_1070),
.Y(n_1185)
);

AOI31xp67_ASAP7_75t_L g1186 ( 
.A1(n_990),
.A2(n_1078),
.A3(n_1090),
.B(n_1042),
.Y(n_1186)
);

INVxp67_ASAP7_75t_SL g1187 ( 
.A(n_980),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1070),
.B(n_1090),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1069),
.A2(n_1084),
.B(n_1108),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_980),
.B(n_1084),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1086),
.A2(n_1070),
.B(n_1090),
.C(n_993),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1086),
.A2(n_1106),
.B(n_1101),
.Y(n_1192)
);

BUFx12f_ASAP7_75t_L g1193 ( 
.A(n_1086),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_L g1194 ( 
.A(n_1036),
.B(n_825),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1014),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1014),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1197)
);

AO32x2_ASAP7_75t_L g1198 ( 
.A1(n_1109),
.A2(n_1111),
.A3(n_1031),
.B1(n_1017),
.B2(n_975),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1085),
.A2(n_1079),
.A3(n_913),
.B(n_1080),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_SL g1200 ( 
.A(n_1036),
.B(n_475),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_984),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1106),
.A2(n_1101),
.B(n_839),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1014),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_SL g1206 ( 
.A(n_1036),
.B(n_475),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1106),
.A2(n_1101),
.B(n_839),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1106),
.B(n_1116),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1061),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_989),
.Y(n_1210)
);

AOI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1020),
.A2(n_1011),
.B(n_1100),
.Y(n_1211)
);

INVx8_ASAP7_75t_L g1212 ( 
.A(n_1086),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1106),
.B(n_1116),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1062),
.Y(n_1214)
);

AO31x2_ASAP7_75t_L g1215 ( 
.A1(n_1085),
.A2(n_1079),
.A3(n_913),
.B(n_1080),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_SL g1216 ( 
.A1(n_1032),
.A2(n_1116),
.B(n_1098),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1085),
.A2(n_1079),
.A3(n_913),
.B(n_1080),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1020),
.A2(n_1011),
.B(n_1100),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_989),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1100),
.A2(n_1105),
.B(n_1113),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1104),
.B(n_801),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1110),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1061),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1101),
.C(n_656),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1101),
.C(n_656),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1014),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_SL g1228 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1098),
.C(n_1111),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1014),
.Y(n_1229)
);

NAND3x1_ASAP7_75t_L g1230 ( 
.A(n_1101),
.B(n_816),
.C(n_1106),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1014),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1110),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_989),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_L g1235 ( 
.A(n_1062),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1085),
.A2(n_1079),
.A3(n_913),
.B(n_1080),
.Y(n_1237)
);

AND2x6_ASAP7_75t_L g1238 ( 
.A(n_990),
.B(n_935),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1062),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1062),
.Y(n_1240)
);

NAND3xp33_ASAP7_75t_L g1241 ( 
.A(n_1101),
.B(n_1106),
.C(n_672),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_989),
.Y(n_1242)
);

INVx5_ASAP7_75t_L g1243 ( 
.A(n_989),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_989),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1100),
.A2(n_1105),
.B(n_1113),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1247)
);

CKINVDCx11_ASAP7_75t_R g1248 ( 
.A(n_1007),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1062),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1101),
.A2(n_848),
.B(n_672),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1106),
.B(n_1116),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1101),
.C(n_656),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1032),
.A2(n_1116),
.B(n_1098),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1085),
.A2(n_1079),
.A3(n_913),
.B(n_1080),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1116),
.A2(n_1106),
.B(n_1098),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1110),
.Y(n_1256)
);

AO31x2_ASAP7_75t_L g1257 ( 
.A1(n_1085),
.A2(n_1079),
.A3(n_913),
.B(n_1080),
.Y(n_1257)
);

CKINVDCx16_ASAP7_75t_R g1258 ( 
.A(n_1110),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1100),
.A2(n_1105),
.B(n_1113),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1106),
.A2(n_1116),
.B(n_1101),
.C(n_656),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1106),
.B(n_1116),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1100),
.A2(n_1105),
.B(n_1113),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1106),
.A2(n_1101),
.B(n_839),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1128),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1208),
.B(n_1213),
.Y(n_1265)
);

CKINVDCx6p67_ASAP7_75t_R g1266 ( 
.A(n_1235),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1258),
.A2(n_1166),
.B1(n_1241),
.B2(n_1263),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1131),
.A2(n_1250),
.B1(n_1125),
.B2(n_1261),
.Y(n_1268)
);

INVx6_ASAP7_75t_L g1269 ( 
.A(n_1132),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1248),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1212),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1251),
.A2(n_1119),
.B1(n_1122),
.B2(n_1207),
.Y(n_1272)
);

INVx6_ASAP7_75t_L g1273 ( 
.A(n_1132),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1222),
.A2(n_1150),
.B1(n_1203),
.B2(n_1137),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1155),
.A2(n_1120),
.B1(n_1197),
.B2(n_1255),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1134),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1212),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1238),
.A2(n_1126),
.B1(n_1142),
.B2(n_1247),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1139),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1141),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1165),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_SL g1282 ( 
.A1(n_1223),
.A2(n_1232),
.B1(n_1256),
.B2(n_1135),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1167),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1169),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1249),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1172),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1195),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1169),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1196),
.Y(n_1289)
);

BUFx8_ASAP7_75t_L g1290 ( 
.A(n_1214),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1238),
.A2(n_1244),
.B1(n_1201),
.B2(n_1217),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1204),
.A2(n_1236),
.B1(n_1234),
.B2(n_1238),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1239),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1205),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1225),
.B(n_1226),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1238),
.A2(n_1160),
.B1(n_1224),
.B2(n_1153),
.Y(n_1296)
);

BUFx8_ASAP7_75t_L g1297 ( 
.A(n_1240),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1230),
.A2(n_1252),
.B1(n_1260),
.B2(n_1216),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1202),
.B(n_1163),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1227),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1198),
.A2(n_1192),
.B1(n_1129),
.B2(n_1209),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1153),
.A2(n_1209),
.B1(n_1224),
.B2(n_1229),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1193),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1140),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1231),
.A2(n_1174),
.B1(n_1157),
.B2(n_1181),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1169),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1200),
.A2(n_1206),
.B1(n_1198),
.B2(n_1162),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1253),
.A2(n_1144),
.B1(n_1151),
.B2(n_1149),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1188),
.Y(n_1309)
);

OAI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1187),
.A2(n_1190),
.B1(n_1157),
.B2(n_1178),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1164),
.A2(n_1194),
.B1(n_1161),
.B2(n_1177),
.Y(n_1311)
);

CKINVDCx11_ASAP7_75t_R g1312 ( 
.A(n_1210),
.Y(n_1312)
);

INVx2_ASAP7_75t_R g1313 ( 
.A(n_1186),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1182),
.Y(n_1314)
);

BUFx8_ASAP7_75t_L g1315 ( 
.A(n_1210),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1148),
.Y(n_1316)
);

BUFx2_ASAP7_75t_SL g1317 ( 
.A(n_1243),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1198),
.A2(n_1143),
.B1(n_1123),
.B2(n_1173),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1188),
.Y(n_1319)
);

BUFx10_ASAP7_75t_L g1320 ( 
.A(n_1220),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1176),
.A2(n_1175),
.B1(n_1136),
.B2(n_1243),
.Y(n_1321)
);

BUFx2_ASAP7_75t_SL g1322 ( 
.A(n_1243),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1164),
.A2(n_1245),
.B1(n_1179),
.B2(n_1189),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_1220),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1123),
.A2(n_1242),
.B1(n_1233),
.B2(n_1121),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1123),
.A2(n_1242),
.B1(n_1233),
.B2(n_1245),
.Y(n_1326)
);

BUFx8_ASAP7_75t_SL g1327 ( 
.A(n_1242),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1123),
.A2(n_1156),
.B1(n_1228),
.B2(n_1185),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1127),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1184),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1145),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1180),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1191),
.A2(n_1183),
.B1(n_1168),
.B2(n_1147),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1143),
.A2(n_1171),
.B1(n_1158),
.B2(n_1152),
.Y(n_1334)
);

INVx5_ASAP7_75t_L g1335 ( 
.A(n_1154),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1143),
.Y(n_1336)
);

INVx6_ASAP7_75t_L g1337 ( 
.A(n_1130),
.Y(n_1337)
);

INVx8_ASAP7_75t_L g1338 ( 
.A(n_1130),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1138),
.A2(n_1257),
.B1(n_1237),
.B2(n_1218),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1159),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1138),
.A2(n_1257),
.B1(n_1237),
.B2(n_1218),
.Y(n_1341)
);

NAND2x1p5_ASAP7_75t_L g1342 ( 
.A(n_1170),
.B(n_1146),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1159),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1133),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1170),
.A2(n_1146),
.B1(n_1138),
.B2(n_1259),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1199),
.B(n_1237),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1211),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1219),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1199),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1262),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1221),
.A2(n_1246),
.B1(n_1218),
.B2(n_1215),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1215),
.A2(n_816),
.B1(n_1131),
.B2(n_491),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1215),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1254),
.A2(n_1106),
.B1(n_1116),
.B2(n_1250),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1254),
.B(n_1257),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1254),
.A2(n_816),
.B1(n_1131),
.B2(n_1101),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1131),
.A2(n_816),
.B1(n_1101),
.B2(n_1106),
.Y(n_1357)
);

BUFx10_ASAP7_75t_L g1358 ( 
.A(n_1223),
.Y(n_1358)
);

INVx4_ASAP7_75t_L g1359 ( 
.A(n_1212),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1212),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1193),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1212),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1250),
.A2(n_1106),
.B1(n_1116),
.B2(n_1241),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1128),
.Y(n_1364)
);

BUFx3_ASAP7_75t_L g1365 ( 
.A(n_1193),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1188),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1131),
.A2(n_816),
.B1(n_491),
.B2(n_1109),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1148),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1128),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1140),
.Y(n_1370)
);

BUFx8_ASAP7_75t_SL g1371 ( 
.A(n_1235),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1235),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1193),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1131),
.A2(n_816),
.B1(n_1101),
.B2(n_1106),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1235),
.Y(n_1375)
);

CKINVDCx11_ASAP7_75t_R g1376 ( 
.A(n_1235),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1250),
.A2(n_1106),
.B1(n_1116),
.B2(n_1241),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1128),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1128),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1124),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1131),
.A2(n_816),
.B1(n_1101),
.B2(n_1106),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1188),
.Y(n_1382)
);

BUFx10_ASAP7_75t_L g1383 ( 
.A(n_1223),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1235),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1208),
.B(n_1213),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1370),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1338),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1335),
.Y(n_1388)
);

AOI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1298),
.A2(n_1354),
.B(n_1308),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1338),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1346),
.A2(n_1355),
.B(n_1345),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1348),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1367),
.A2(n_1374),
.B1(n_1357),
.B2(n_1381),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1342),
.A2(n_1345),
.B(n_1351),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1299),
.Y(n_1395)
);

INVx6_ASAP7_75t_L g1396 ( 
.A(n_1315),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1336),
.Y(n_1397)
);

AOI21xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1268),
.A2(n_1377),
.B(n_1363),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1351),
.A2(n_1292),
.B(n_1275),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1264),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1292),
.A2(n_1275),
.B(n_1331),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1279),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1280),
.Y(n_1403)
);

AOI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1295),
.A2(n_1311),
.B(n_1340),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1281),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1283),
.Y(n_1406)
);

BUFx8_ASAP7_75t_L g1407 ( 
.A(n_1375),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1265),
.B(n_1385),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1287),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1338),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1337),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1343),
.B(n_1335),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1289),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1356),
.A2(n_1349),
.B(n_1302),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1294),
.Y(n_1415)
);

AOI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1333),
.A2(n_1329),
.B(n_1332),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1300),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1328),
.A2(n_1356),
.B(n_1296),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1364),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1369),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1268),
.B(n_1302),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1378),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1350),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1379),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1296),
.A2(n_1328),
.B(n_1374),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1353),
.Y(n_1426)
);

BUFx8_ASAP7_75t_SL g1427 ( 
.A(n_1371),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1272),
.B(n_1357),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1334),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1272),
.A2(n_1367),
.B1(n_1307),
.B2(n_1368),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1301),
.B(n_1318),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1301),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1318),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1319),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1344),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1339),
.B(n_1341),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1339),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1341),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1334),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1309),
.B(n_1366),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1305),
.A2(n_1382),
.B(n_1381),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1307),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1278),
.B(n_1352),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1347),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1313),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1269),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1274),
.A2(n_1380),
.B(n_1291),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1278),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1352),
.A2(n_1274),
.B1(n_1267),
.B2(n_1291),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1321),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1323),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1323),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1310),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1273),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1314),
.B(n_1304),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1304),
.B(n_1312),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1325),
.A2(n_1326),
.B(n_1276),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1361),
.A2(n_1373),
.B1(n_1365),
.B2(n_1316),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1312),
.B(n_1320),
.Y(n_1459)
);

AO32x2_ASAP7_75t_L g1460 ( 
.A1(n_1393),
.A2(n_1411),
.A3(n_1390),
.B1(n_1387),
.B2(n_1410),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1395),
.B(n_1315),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1396),
.Y(n_1462)
);

AO32x2_ASAP7_75t_L g1463 ( 
.A1(n_1411),
.A2(n_1282),
.A3(n_1360),
.B1(n_1359),
.B2(n_1327),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1412),
.B(n_1361),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1405),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1386),
.B(n_1373),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1430),
.A2(n_1293),
.B1(n_1285),
.B2(n_1306),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1398),
.B(n_1288),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1428),
.A2(n_1398),
.B(n_1449),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1386),
.B(n_1372),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1388),
.Y(n_1471)
);

OAI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1389),
.A2(n_1360),
.B(n_1359),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_SL g1473 ( 
.A1(n_1421),
.A2(n_1270),
.B(n_1317),
.C(n_1322),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1417),
.B(n_1266),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1400),
.B(n_1402),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1443),
.A2(n_1284),
.B(n_1288),
.C(n_1330),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1434),
.B(n_1444),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1443),
.A2(n_1432),
.B1(n_1431),
.B2(n_1442),
.C(n_1429),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1444),
.Y(n_1479)
);

A2O1A1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1421),
.A2(n_1288),
.B(n_1330),
.C(n_1277),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1444),
.B(n_1306),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1423),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1425),
.A2(n_1376),
.B1(n_1384),
.B2(n_1303),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1391),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1400),
.B(n_1402),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1442),
.A2(n_1271),
.B(n_1277),
.C(n_1362),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1423),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1444),
.B(n_1383),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1425),
.A2(n_1376),
.B1(n_1297),
.B2(n_1290),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1456),
.B(n_1358),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1448),
.A2(n_1271),
.B1(n_1277),
.B2(n_1290),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1456),
.B(n_1358),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1394),
.A2(n_1324),
.B(n_1297),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1408),
.B(n_1324),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1459),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1389),
.A2(n_1383),
.B(n_1270),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1403),
.B(n_1286),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1425),
.A2(n_1286),
.B1(n_1431),
.B2(n_1432),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1403),
.B(n_1406),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1425),
.A2(n_1399),
.B(n_1418),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1406),
.Y(n_1501)
);

NAND2xp33_ASAP7_75t_R g1502 ( 
.A(n_1457),
.B(n_1447),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1440),
.B(n_1409),
.Y(n_1503)
);

AO32x2_ASAP7_75t_L g1504 ( 
.A1(n_1387),
.A2(n_1390),
.A3(n_1410),
.B1(n_1446),
.B2(n_1458),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1413),
.Y(n_1505)
);

OA21x2_ASAP7_75t_L g1506 ( 
.A1(n_1394),
.A2(n_1399),
.B(n_1418),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1440),
.B(n_1415),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1454),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1445),
.Y(n_1509)
);

AOI221xp5_ASAP7_75t_L g1510 ( 
.A1(n_1439),
.A2(n_1433),
.B1(n_1437),
.B2(n_1438),
.C(n_1436),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1404),
.A2(n_1401),
.B(n_1416),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1433),
.A2(n_1437),
.B1(n_1438),
.B2(n_1436),
.Y(n_1512)
);

A2O1A1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1439),
.A2(n_1441),
.B(n_1451),
.C(n_1452),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1453),
.A2(n_1447),
.B1(n_1452),
.B2(n_1451),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1419),
.B(n_1420),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1501),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1505),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1509),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1484),
.B(n_1392),
.Y(n_1519)
);

INVxp67_ASAP7_75t_SL g1520 ( 
.A(n_1484),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1469),
.A2(n_1447),
.B1(n_1414),
.B2(n_1453),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1477),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1475),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1503),
.B(n_1507),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1485),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1465),
.B(n_1397),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1499),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1515),
.B(n_1513),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1506),
.B(n_1391),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1482),
.B(n_1391),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1482),
.B(n_1423),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1487),
.B(n_1391),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1500),
.B(n_1397),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1487),
.B(n_1460),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1460),
.B(n_1435),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1508),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1460),
.B(n_1435),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1467),
.A2(n_1447),
.B1(n_1404),
.B2(n_1414),
.Y(n_1538)
);

AOI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1478),
.A2(n_1414),
.B1(n_1441),
.B2(n_1457),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1513),
.B(n_1422),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1479),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1518),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1538),
.B(n_1511),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1534),
.B(n_1460),
.Y(n_1544)
);

NAND5xp2_ASAP7_75t_L g1545 ( 
.A(n_1521),
.B(n_1496),
.C(n_1489),
.D(n_1472),
.E(n_1473),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1519),
.Y(n_1546)
);

AOI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1528),
.A2(n_1510),
.B1(n_1512),
.B2(n_1498),
.C(n_1514),
.Y(n_1547)
);

INVxp67_ASAP7_75t_L g1548 ( 
.A(n_1536),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1531),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1521),
.A2(n_1512),
.B1(n_1414),
.B2(n_1450),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1519),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1518),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1534),
.B(n_1504),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1534),
.B(n_1504),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1516),
.Y(n_1555)
);

NAND4xp25_ASAP7_75t_L g1556 ( 
.A(n_1538),
.B(n_1497),
.C(n_1468),
.D(n_1474),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1504),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1539),
.A2(n_1483),
.B1(n_1426),
.B2(n_1468),
.Y(n_1558)
);

AOI211xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1539),
.A2(n_1473),
.B(n_1480),
.C(n_1476),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1528),
.A2(n_1476),
.B1(n_1480),
.B2(n_1486),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1520),
.Y(n_1561)
);

AND2x4_ASAP7_75t_SL g1562 ( 
.A(n_1536),
.B(n_1464),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1530),
.B(n_1504),
.Y(n_1563)
);

OAI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1540),
.A2(n_1502),
.B1(n_1486),
.B2(n_1491),
.C(n_1416),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1540),
.A2(n_1495),
.B1(n_1494),
.B2(n_1462),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1532),
.B(n_1535),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1532),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1535),
.A2(n_1502),
.B1(n_1493),
.B2(n_1457),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1529),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1529),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1424),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1531),
.B(n_1471),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1547),
.A2(n_1529),
.B1(n_1537),
.B2(n_1533),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1569),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_SL g1577 ( 
.A(n_1559),
.B(n_1537),
.C(n_1461),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1553),
.B(n_1524),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1571),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1542),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1554),
.B(n_1537),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1544),
.B(n_1546),
.Y(n_1582)
);

INVxp33_ASAP7_75t_L g1583 ( 
.A(n_1564),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1554),
.B(n_1522),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1554),
.B(n_1522),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1571),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1571),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1544),
.B(n_1526),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1557),
.B(n_1541),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1547),
.A2(n_1462),
.B1(n_1527),
.B2(n_1525),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1542),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1569),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1551),
.B(n_1517),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1551),
.B(n_1517),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1544),
.B(n_1526),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1555),
.Y(n_1596)
);

AND2x4_ASAP7_75t_SL g1597 ( 
.A(n_1543),
.B(n_1572),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1549),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1569),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1557),
.B(n_1523),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1563),
.B(n_1523),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1563),
.B(n_1527),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1555),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1562),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1583),
.B(n_1556),
.Y(n_1605)
);

NOR2x1_ASAP7_75t_L g1606 ( 
.A(n_1577),
.B(n_1556),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1596),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1573),
.B(n_1561),
.Y(n_1608)
);

NOR2x1p5_ASAP7_75t_L g1609 ( 
.A(n_1577),
.B(n_1549),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1596),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1575),
.B(n_1566),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1583),
.A2(n_1559),
.B1(n_1543),
.B2(n_1564),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1582),
.B(n_1552),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1596),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1573),
.A2(n_1543),
.B1(n_1560),
.B2(n_1558),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1603),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1574),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1590),
.B(n_1565),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1603),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1575),
.B(n_1566),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1575),
.B(n_1566),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1590),
.B(n_1561),
.Y(n_1622)
);

INVxp67_ASAP7_75t_L g1623 ( 
.A(n_1580),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1597),
.B(n_1543),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1574),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1582),
.B(n_1552),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1603),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1574),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1593),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1576),
.B(n_1562),
.Y(n_1630)
);

INVxp67_ASAP7_75t_L g1631 ( 
.A(n_1580),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1574),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1588),
.B(n_1543),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1593),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1594),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

NAND2x1_ASAP7_75t_L g1637 ( 
.A(n_1604),
.B(n_1561),
.Y(n_1637)
);

NAND2x2_ASAP7_75t_L g1638 ( 
.A(n_1604),
.B(n_1427),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1592),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1576),
.B(n_1548),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1582),
.B(n_1588),
.Y(n_1641)
);

NAND2x1p5_ASAP7_75t_L g1642 ( 
.A(n_1604),
.B(n_1464),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1597),
.B(n_1543),
.Y(n_1643)
);

OAI21xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1581),
.A2(n_1543),
.B(n_1567),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1597),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1584),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1576),
.B(n_1562),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1607),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1609),
.B(n_1646),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1645),
.B(n_1597),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1605),
.B(n_1612),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1641),
.B(n_1588),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1610),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1605),
.B(n_1578),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1645),
.B(n_1578),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1606),
.B(n_1578),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1629),
.B(n_1634),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1635),
.B(n_1600),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1617),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1630),
.B(n_1581),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1614),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1618),
.B(n_1407),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1630),
.B(n_1581),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1647),
.B(n_1589),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1608),
.A2(n_1545),
.B1(n_1570),
.B2(n_1579),
.C(n_1558),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1647),
.B(n_1589),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1616),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1636),
.B(n_1600),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1615),
.B(n_1623),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1631),
.B(n_1600),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1611),
.B(n_1598),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1619),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1618),
.B(n_1601),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1627),
.B(n_1601),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1622),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1641),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1617),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1613),
.Y(n_1678)
);

BUFx3_ASAP7_75t_L g1679 ( 
.A(n_1637),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1611),
.B(n_1598),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1613),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1624),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1626),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1682),
.Y(n_1684)
);

AOI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1651),
.A2(n_1644),
.B(n_1633),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1650),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1662),
.A2(n_1643),
.B1(n_1624),
.B2(n_1642),
.Y(n_1687)
);

OA21x2_ASAP7_75t_L g1688 ( 
.A1(n_1665),
.A2(n_1628),
.B(n_1625),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1667),
.Y(n_1689)
);

NAND2xp33_ASAP7_75t_SL g1690 ( 
.A(n_1656),
.B(n_1626),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1667),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1665),
.A2(n_1560),
.B1(n_1568),
.B2(n_1550),
.Y(n_1692)
);

AOI32xp33_ASAP7_75t_L g1693 ( 
.A1(n_1656),
.A2(n_1643),
.A3(n_1624),
.B1(n_1585),
.B2(n_1584),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1648),
.Y(n_1694)
);

OAI322xp33_ASAP7_75t_L g1695 ( 
.A1(n_1675),
.A2(n_1640),
.A3(n_1595),
.B1(n_1579),
.B2(n_1586),
.C1(n_1587),
.C2(n_1565),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1669),
.A2(n_1568),
.B1(n_1550),
.B2(n_1639),
.C(n_1632),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1648),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1682),
.Y(n_1698)
);

AO22x1_ASAP7_75t_L g1699 ( 
.A1(n_1679),
.A2(n_1643),
.B1(n_1407),
.B2(n_1598),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1653),
.Y(n_1700)
);

AOI21xp33_ASAP7_75t_L g1701 ( 
.A1(n_1675),
.A2(n_1628),
.B(n_1625),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1669),
.A2(n_1585),
.B(n_1584),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1654),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1673),
.A2(n_1585),
.B(n_1591),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1673),
.A2(n_1545),
.B(n_1591),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1653),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_SL g1707 ( 
.A(n_1649),
.B(n_1407),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1679),
.B(n_1481),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1684),
.B(n_1654),
.Y(n_1709)
);

AOI222xp33_ASAP7_75t_L g1710 ( 
.A1(n_1696),
.A2(n_1690),
.B1(n_1702),
.B2(n_1704),
.C1(n_1703),
.C2(n_1688),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1694),
.Y(n_1711)
);

AOI21xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1688),
.A2(n_1708),
.B(n_1699),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1689),
.B(n_1678),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1697),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1700),
.Y(n_1715)
);

OAI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1692),
.A2(n_1649),
.B1(n_1679),
.B2(n_1676),
.C(n_1652),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1698),
.B(n_1676),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1706),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1691),
.B(n_1678),
.Y(n_1719)
);

O2A1O1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1705),
.A2(n_1683),
.B(n_1681),
.C(n_1670),
.Y(n_1720)
);

AOI21xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1708),
.A2(n_1683),
.B(n_1681),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_SL g1722 ( 
.A1(n_1704),
.A2(n_1670),
.B(n_1652),
.C(n_1657),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1686),
.B(n_1663),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1702),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1701),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1693),
.B(n_1663),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1695),
.A2(n_1657),
.B1(n_1661),
.B2(n_1672),
.C(n_1677),
.Y(n_1727)
);

OAI21xp33_ASAP7_75t_L g1728 ( 
.A1(n_1707),
.A2(n_1650),
.B(n_1655),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1717),
.Y(n_1729)
);

AOI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1725),
.A2(n_1677),
.B(n_1659),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1713),
.Y(n_1731)
);

INVxp67_ASAP7_75t_L g1732 ( 
.A(n_1724),
.Y(n_1732)
);

NAND2x1_ASAP7_75t_L g1733 ( 
.A(n_1723),
.B(n_1655),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1709),
.B(n_1663),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1713),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1719),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1710),
.B(n_1701),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1719),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1734),
.B(n_1721),
.Y(n_1739)
);

NAND4xp25_ASAP7_75t_SL g1740 ( 
.A(n_1737),
.B(n_1720),
.C(n_1716),
.D(n_1726),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_L g1741 ( 
.A(n_1737),
.B(n_1712),
.C(n_1722),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1732),
.A2(n_1727),
.B1(n_1685),
.B2(n_1718),
.C(n_1715),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1738),
.B(n_1711),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1729),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1730),
.Y(n_1745)
);

AND4x1_ASAP7_75t_L g1746 ( 
.A(n_1731),
.B(n_1728),
.C(n_1714),
.D(n_1407),
.Y(n_1746)
);

NOR3xp33_ASAP7_75t_L g1747 ( 
.A(n_1738),
.B(n_1687),
.C(n_1677),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1741),
.A2(n_1736),
.B(n_1735),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1745),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1740),
.A2(n_1733),
.B1(n_1659),
.B2(n_1661),
.C(n_1672),
.Y(n_1750)
);

AO22x2_ASAP7_75t_L g1751 ( 
.A1(n_1739),
.A2(n_1659),
.B1(n_1660),
.B2(n_1680),
.Y(n_1751)
);

OAI211xp5_ASAP7_75t_L g1752 ( 
.A1(n_1742),
.A2(n_1680),
.B(n_1671),
.C(n_1658),
.Y(n_1752)
);

AOI221xp5_ASAP7_75t_L g1753 ( 
.A1(n_1749),
.A2(n_1744),
.B1(n_1747),
.B2(n_1743),
.C(n_1746),
.Y(n_1753)
);

NAND4xp25_ASAP7_75t_SL g1754 ( 
.A(n_1750),
.B(n_1680),
.C(n_1671),
.D(n_1660),
.Y(n_1754)
);

AOI211xp5_ASAP7_75t_L g1755 ( 
.A1(n_1748),
.A2(n_1658),
.B(n_1668),
.C(n_1671),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1751),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1752),
.A2(n_1666),
.B1(n_1664),
.B2(n_1668),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1751),
.B(n_1664),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1756),
.Y(n_1759)
);

XOR2xp5_ASAP7_75t_L g1760 ( 
.A(n_1758),
.B(n_1455),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1757),
.Y(n_1761)
);

NOR2xp67_ASAP7_75t_L g1762 ( 
.A(n_1754),
.B(n_1674),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1755),
.B(n_1666),
.Y(n_1763)
);

NOR2x1_ASAP7_75t_L g1764 ( 
.A(n_1759),
.B(n_1753),
.Y(n_1764)
);

A2O1A1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1759),
.A2(n_1632),
.B(n_1639),
.C(n_1674),
.Y(n_1765)
);

NOR3xp33_ASAP7_75t_L g1766 ( 
.A(n_1761),
.B(n_1492),
.C(n_1490),
.Y(n_1766)
);

XNOR2xp5_ASAP7_75t_L g1767 ( 
.A(n_1764),
.B(n_1760),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1767),
.A2(n_1763),
.B1(n_1762),
.B2(n_1766),
.Y(n_1768)
);

AOI22x1_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1765),
.B1(n_1598),
.B2(n_1620),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1768),
.A2(n_1638),
.B1(n_1595),
.B2(n_1621),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1769),
.A2(n_1638),
.B1(n_1621),
.B2(n_1620),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1770),
.A2(n_1396),
.B1(n_1599),
.B2(n_1592),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1592),
.B1(n_1599),
.B2(n_1579),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1771),
.A2(n_1592),
.B(n_1599),
.Y(n_1774)
);

AOI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1595),
.B(n_1599),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1773),
.B(n_1602),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1396),
.B1(n_1586),
.B2(n_1587),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_R g1778 ( 
.A1(n_1777),
.A2(n_1598),
.B1(n_1642),
.B2(n_1548),
.C(n_1463),
.Y(n_1778)
);

AOI211xp5_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1488),
.B(n_1470),
.C(n_1466),
.Y(n_1779)
);


endmodule