module fake_jpeg_28782_n_530 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_530);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_53),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_82),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_81),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_23),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_37),
.B(n_16),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_32),
.B(n_14),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_23),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_23),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_96),
.Y(n_144)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_97),
.B(n_98),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_23),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_32),
.B(n_14),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_106),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_66),
.A2(n_31),
.B(n_32),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_156),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_68),
.B(n_51),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_161),
.Y(n_173)
);

INVx6_ASAP7_75t_SL g134 ( 
.A(n_55),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_134),
.B(n_139),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_75),
.B(n_53),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_141),
.B(n_169),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_86),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_87),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_66),
.B(n_30),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_42),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_61),
.B(n_0),
.Y(n_161)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_59),
.Y(n_167)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_76),
.B(n_19),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_171),
.B(n_211),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_179),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_47),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_192),
.Y(n_225)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_117),
.B(n_18),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_31),
.B(n_47),
.C(n_23),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_180),
.B(n_222),
.Y(n_259)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_110),
.A2(n_51),
.B1(n_70),
.B2(n_100),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_182),
.A2(n_190),
.B1(n_197),
.B2(n_202),
.Y(n_233)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_131),
.A2(n_95),
.B(n_102),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_184),
.A2(n_107),
.B(n_84),
.Y(n_238)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_107),
.B(n_50),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_189),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_128),
.A2(n_51),
.B1(n_83),
.B2(n_50),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_35),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_137),
.Y(n_193)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_109),
.A2(n_65),
.B1(n_99),
.B2(n_104),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_200),
.B1(n_145),
.B2(n_152),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_64),
.B1(n_69),
.B2(n_85),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_195),
.A2(n_203),
.B1(n_152),
.B2(n_145),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_117),
.B(n_18),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_198),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_129),
.A2(n_50),
.B1(n_52),
.B2(n_20),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_114),
.B(n_18),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_114),
.A2(n_74),
.B1(n_77),
.B2(n_80),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_124),
.A2(n_50),
.B1(n_45),
.B2(n_52),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_115),
.A2(n_20),
.B1(n_45),
.B2(n_52),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_133),
.A2(n_20),
.B1(n_45),
.B2(n_40),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_144),
.B(n_19),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_167),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_140),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_210),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_146),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_111),
.A2(n_40),
.B1(n_30),
.B2(n_42),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_148),
.Y(n_215)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_160),
.B(n_105),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_157),
.C(n_108),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_130),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_221),
.Y(n_252)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_146),
.B(n_35),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_108),
.B(n_18),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_175),
.A2(n_214),
.B1(n_176),
.B2(n_173),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_226),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_173),
.A2(n_126),
.B1(n_162),
.B2(n_154),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_173),
.A2(n_126),
.B1(n_162),
.B2(n_154),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_241),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_262),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_246),
.B(n_209),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_188),
.A2(n_165),
.B1(n_135),
.B2(n_150),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_248),
.A2(n_127),
.B1(n_201),
.B2(n_191),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_249),
.B(n_170),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_216),
.B(n_136),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_260),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_172),
.B(n_132),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_180),
.A2(n_168),
.B1(n_140),
.B2(n_112),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_166),
.B1(n_143),
.B2(n_142),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_263),
.A2(n_127),
.B1(n_205),
.B2(n_178),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_184),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_266),
.A2(n_274),
.B(n_282),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_225),
.B(n_192),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_271),
.Y(n_302)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_270),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_292),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_232),
.A2(n_187),
.B1(n_194),
.B2(n_181),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_170),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_238),
.B(n_186),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_277),
.B(n_288),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_221),
.B1(n_207),
.B2(n_183),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_287),
.B1(n_294),
.B2(n_300),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_228),
.A2(n_206),
.B1(n_210),
.B2(n_177),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_225),
.B(n_185),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_284),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_215),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_285),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_286),
.A2(n_261),
.B1(n_236),
.B2(n_255),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_240),
.A2(n_193),
.B1(n_218),
.B2(n_174),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_259),
.B(n_201),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_178),
.C(n_204),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_293),
.Y(n_305)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_230),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_291),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_247),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_224),
.B(n_219),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_243),
.A2(n_217),
.B1(n_213),
.B2(n_199),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_245),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_296),
.Y(n_308)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_171),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_248),
.Y(n_306)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_265),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_299),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_253),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_268),
.A2(n_272),
.B1(n_273),
.B2(n_277),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_303),
.A2(n_310),
.B1(n_314),
.B2(n_319),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_SL g363 ( 
.A1(n_306),
.A2(n_229),
.B(n_250),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_268),
.A2(n_277),
.B1(n_266),
.B2(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_224),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_316),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_278),
.A2(n_233),
.B1(n_246),
.B2(n_234),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_237),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_259),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_320),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_278),
.A2(n_274),
.B1(n_284),
.B2(n_283),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_269),
.B(n_237),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_276),
.A2(n_258),
.B(n_242),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_322),
.A2(n_298),
.B(n_296),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_231),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_327),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_276),
.A2(n_258),
.B(n_254),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_325),
.A2(n_253),
.B(n_279),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_329),
.Y(n_336)
);

AOI32xp33_ASAP7_75t_L g330 ( 
.A1(n_276),
.A2(n_289),
.A3(n_297),
.B1(n_294),
.B2(n_275),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_261),
.Y(n_345)
);

NOR2x1_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_256),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_301),
.Y(n_361)
);

O2A1O1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_306),
.A2(n_300),
.B(n_286),
.C(n_254),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_349),
.Y(n_368)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_337),
.B(n_340),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_338),
.A2(n_343),
.B(n_345),
.Y(n_391)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_332),
.Y(n_339)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

NOR3xp33_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_292),
.C(n_290),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_285),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_302),
.Y(n_383)
);

INVx13_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_344),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_305),
.B(n_325),
.C(n_320),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_353),
.C(n_325),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_324),
.A2(n_239),
.B1(n_255),
.B2(n_236),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_347),
.A2(n_363),
.B1(n_329),
.B2(n_321),
.Y(n_387)
);

AOI21xp33_ASAP7_75t_SL g348 ( 
.A1(n_323),
.A2(n_291),
.B(n_230),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_348),
.A2(n_350),
.B(n_354),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_270),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_310),
.A2(n_291),
.B(n_204),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_308),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_352),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_308),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_305),
.B(n_247),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_331),
.A2(n_230),
.B(n_251),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_331),
.A2(n_227),
.B(n_251),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_360),
.Y(n_369)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_333),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_362),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_312),
.B(n_229),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_261),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_311),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_319),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_373),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_319),
.Y(n_373)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_356),
.B(n_326),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_375),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_304),
.Y(n_376)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_383),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_352),
.B(n_304),
.Y(n_379)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_379),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_327),
.Y(n_382)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_342),
.B(n_310),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_317),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_328),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_386),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_336),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_328),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_389),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_311),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_330),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_390),
.B(n_395),
.C(n_309),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_345),
.A2(n_317),
.B1(n_313),
.B2(n_309),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g418 ( 
.A1(n_392),
.A2(n_397),
.B1(n_372),
.B2(n_387),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_303),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_393),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_361),
.B(n_322),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_394),
.B(n_396),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_322),
.C(n_303),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_419),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_390),
.A2(n_336),
.B1(n_350),
.B2(n_343),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_405),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_404),
.A2(n_420),
.B1(n_370),
.B2(n_394),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_391),
.A2(n_338),
.B(n_354),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_381),
.B(n_365),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_408),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_396),
.A2(n_336),
.B1(n_314),
.B2(n_347),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_359),
.Y(n_409)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_409),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_SL g411 ( 
.A(n_391),
.B(n_314),
.C(n_334),
.Y(n_411)
);

AOI21xp33_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_371),
.B(n_369),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_367),
.B(n_362),
.C(n_355),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_416),
.C(n_373),
.Y(n_426)
);

AO21x2_ASAP7_75t_L g415 ( 
.A1(n_368),
.A2(n_334),
.B(n_344),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_415),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_378),
.B(n_360),
.C(n_335),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_421),
.Y(n_438)
);

A2O1A1Ixp33_ASAP7_75t_SL g420 ( 
.A1(n_397),
.A2(n_317),
.B(n_344),
.C(n_321),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_389),
.B(n_357),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_383),
.B(n_315),
.Y(n_424)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_424),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_370),
.A2(n_339),
.B1(n_358),
.B2(n_315),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_369),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_433),
.C(n_440),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_427),
.A2(n_429),
.B1(n_442),
.B2(n_399),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_419),
.A2(n_384),
.B1(n_395),
.B2(n_368),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_413),
.B(n_393),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_432),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_382),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_416),
.B(n_374),
.C(n_379),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_412),
.Y(n_435)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_422),
.Y(n_436)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_436),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_376),
.C(n_371),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_401),
.Y(n_441)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_441),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_411),
.A2(n_377),
.B1(n_380),
.B2(n_385),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_443),
.A2(n_415),
.B(n_420),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_444),
.A2(n_400),
.B1(n_410),
.B2(n_423),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_414),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_366),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_401),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_447),
.B(n_403),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_402),
.B(n_385),
.C(n_380),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_405),
.C(n_425),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_450),
.Y(n_479)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_452),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_430),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_465),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_444),
.B1(n_446),
.B2(n_420),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_456),
.A2(n_27),
.B1(n_41),
.B2(n_33),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_442),
.A2(n_427),
.B1(n_428),
.B2(n_408),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_457),
.A2(n_464),
.B1(n_467),
.B2(n_431),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_459),
.B(n_460),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_426),
.B(n_398),
.C(n_417),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_448),
.C(n_432),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_466),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_439),
.A2(n_366),
.B1(n_377),
.B2(n_420),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_415),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_429),
.A2(n_415),
.B(n_321),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_440),
.A2(n_415),
.B1(n_307),
.B2(n_239),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_445),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_468),
.B(n_482),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_469),
.B(n_473),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_484),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_437),
.C(n_434),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_471),
.B(n_474),
.C(n_480),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_457),
.A2(n_437),
.B1(n_250),
.B2(n_40),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_472),
.A2(n_453),
.B1(n_463),
.B2(n_458),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_451),
.B(n_250),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_40),
.C(n_171),
.Y(n_474)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_476),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_113),
.C(n_41),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_18),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_1),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_483),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_27),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_478),
.A2(n_460),
.B(n_465),
.Y(n_485)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_485),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_456),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_493),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_477),
.A2(n_466),
.B(n_467),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_488),
.A2(n_474),
.B(n_483),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_489),
.A2(n_490),
.B1(n_3),
.B2(n_4),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_479),
.A2(n_453),
.B1(n_455),
.B2(n_27),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_479),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_469),
.B(n_113),
.C(n_41),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_499),
.C(n_491),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_33),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_495),
.B(n_1),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_33),
.C(n_26),
.Y(n_499)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_501),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_509),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_487),
.A2(n_480),
.B(n_26),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_503),
.B(n_506),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_510),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_498),
.B(n_3),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_26),
.B(n_4),
.Y(n_507)
);

AOI221xp5_ASAP7_75t_L g515 ( 
.A1(n_507),
.A2(n_508),
.B1(n_488),
.B2(n_496),
.C(n_6),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_3),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_3),
.Y(n_509)
);

OAI21x1_ASAP7_75t_SL g521 ( 
.A1(n_515),
.A2(n_516),
.B(n_513),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g516 ( 
.A(n_500),
.B(n_497),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_505),
.A2(n_494),
.B1(n_499),
.B2(n_492),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_517),
.A2(n_510),
.B(n_508),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_518),
.B(n_519),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_512),
.A2(n_492),
.B(n_5),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_SL g520 ( 
.A(n_516),
.B(n_4),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_520),
.B(n_5),
.Y(n_524)
);

AOI322xp5_ASAP7_75t_L g523 ( 
.A1(n_521),
.A2(n_514),
.A3(n_511),
.B1(n_7),
.B2(n_8),
.C1(n_5),
.C2(n_12),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_523),
.A2(n_13),
.B(n_7),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_5),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_L g527 ( 
.A1(n_525),
.A2(n_526),
.B(n_522),
.C(n_8),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_6),
.B1(n_11),
.B2(n_13),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_L g529 ( 
.A1(n_528),
.A2(n_6),
.B(n_11),
.C(n_13),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_13),
.Y(n_530)
);


endmodule