module fake_netlist_1_8911_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_25;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_6), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_7), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_9), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_4), .B(n_3), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_8), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_2), .Y(n_18) );
O2A1O1Ixp33_ASAP7_75t_L g19 ( .A1(n_11), .A2(n_0), .B(n_1), .C(n_2), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_12), .B(n_0), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_11), .A2(n_1), .B(n_3), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_15), .A2(n_5), .B(n_7), .Y(n_22) );
NAND2xp5_ASAP7_75t_SL g23 ( .A(n_14), .B(n_5), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_16), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_15), .B1(n_18), .B2(n_13), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_13), .Y(n_26) );
BUFx3_ASAP7_75t_L g27 ( .A(n_22), .Y(n_27) );
BUFx3_ASAP7_75t_L g28 ( .A(n_21), .Y(n_28) );
INVx2_ASAP7_75t_SL g29 ( .A(n_28), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_26), .B(n_23), .Y(n_30) );
OR2x2_ASAP7_75t_L g31 ( .A(n_26), .B(n_8), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AOI222xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_30), .B1(n_25), .B2(n_17), .C1(n_27), .C2(n_28), .Y(n_34) );
NOR2xp33_ASAP7_75t_R g35 ( .A(n_32), .B(n_31), .Y(n_35) );
AOI322xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_25), .A3(n_30), .B1(n_27), .B2(n_28), .C1(n_19), .C2(n_29), .Y(n_36) );
INVx1_ASAP7_75t_SL g37 ( .A(n_35), .Y(n_37) );
OAI22xp5_ASAP7_75t_SL g38 ( .A1(n_37), .A2(n_27), .B1(n_32), .B2(n_9), .Y(n_38) );
NAND2xp5_ASAP7_75t_SL g39 ( .A(n_36), .B(n_10), .Y(n_39) );
AOI22xp5_ASAP7_75t_L g40 ( .A1(n_38), .A2(n_10), .B1(n_36), .B2(n_39), .Y(n_40) );
endmodule