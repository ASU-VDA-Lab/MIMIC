module fake_jpeg_1534_n_338 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_41),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_42),
.B(n_38),
.Y(n_104)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_17),
.B(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_54),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_17),
.B(n_13),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_12),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_65),
.Y(n_93)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_15),
.B(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_11),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_11),
.Y(n_101)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_30),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_75),
.B(n_101),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_30),
.B1(n_32),
.B2(n_15),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_77),
.A2(n_85),
.B1(n_0),
.B2(n_1),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_40),
.A2(n_23),
.B1(n_38),
.B2(n_32),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_80),
.A2(n_96),
.B1(n_99),
.B2(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_41),
.A2(n_18),
.B1(n_31),
.B2(n_35),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_117),
.B1(n_71),
.B2(n_69),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_23),
.B1(n_36),
.B2(n_35),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_48),
.A2(n_31),
.B1(n_23),
.B2(n_34),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_38),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_97),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_34),
.B1(n_28),
.B2(n_20),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_106),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_45),
.B(n_18),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_28),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_110),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_36),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_58),
.A2(n_33),
.B1(n_24),
.B2(n_20),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_27),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_8),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_64),
.A2(n_33),
.B1(n_24),
.B2(n_9),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_61),
.B1(n_72),
.B2(n_53),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_52),
.B1(n_46),
.B2(n_66),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_145),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_124),
.B(n_143),
.Y(n_196)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_103),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_27),
.B1(n_26),
.B2(n_21),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_76),
.A2(n_26),
.B1(n_21),
.B2(n_2),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_128),
.A2(n_138),
.B1(n_149),
.B2(n_160),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_134),
.B1(n_136),
.B2(n_140),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_131),
.Y(n_175)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_133),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_74),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_151),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_8),
.Y(n_145)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_150),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_158),
.Y(n_181)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_159),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_119),
.C(n_88),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_114),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_80),
.B1(n_116),
.B2(n_82),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_131),
.B1(n_160),
.B2(n_151),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_88),
.B1(n_119),
.B2(n_87),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_166),
.A2(n_169),
.B1(n_182),
.B2(n_186),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_83),
.B1(n_87),
.B2(n_86),
.Y(n_169)
);

AO22x1_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_79),
.B1(n_82),
.B2(n_116),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_173),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_130),
.A2(n_114),
.B1(n_115),
.B2(n_86),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_173),
.A2(n_166),
.B1(n_190),
.B2(n_174),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_131),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_134),
.A2(n_115),
.B1(n_79),
.B2(n_82),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_79),
.B(n_145),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_155),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_146),
.B(n_123),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_184),
.B(n_126),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_129),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_188),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_129),
.A2(n_144),
.B1(n_156),
.B2(n_152),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_139),
.B(n_147),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_187),
.A2(n_192),
.B(n_171),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_135),
.B(n_141),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_126),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_210),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_132),
.C(n_137),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_201),
.Y(n_240)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_159),
.C(n_150),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_203),
.B(n_204),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_184),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_205),
.B(n_212),
.Y(n_241)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_226),
.Y(n_233)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_209),
.Y(n_239)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_158),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_149),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_213),
.B(n_214),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_165),
.B(n_133),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_218),
.Y(n_245)
);

AO21x1_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_187),
.B(n_167),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_162),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_219),
.B(n_206),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_180),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_221),
.Y(n_247)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_228),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_164),
.A2(n_167),
.B1(n_163),
.B2(n_196),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_163),
.B(n_192),
.C(n_172),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_SL g248 ( 
.A(n_225),
.B(n_227),
.C(n_223),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_189),
.C(n_172),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_170),
.A2(n_189),
.B1(n_168),
.B2(n_180),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_175),
.B1(n_191),
.B2(n_216),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_231),
.A2(n_211),
.B1(n_200),
.B2(n_221),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_175),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_242),
.C(n_243),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_198),
.B(n_199),
.Y(n_242)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_210),
.C(n_212),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_205),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_244),
.B(n_251),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_202),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_227),
.B(n_223),
.Y(n_262)
);

XOR2x2_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_201),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_218),
.Y(n_256)
);

AND2x6_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_225),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_253),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_268),
.Y(n_279)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_258),
.Y(n_290)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_254),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_263),
.Y(n_277)
);

AO21x2_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_216),
.B(n_222),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_264),
.B1(n_270),
.B2(n_248),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_262),
.A2(n_250),
.B(n_237),
.Y(n_286)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_230),
.A2(n_202),
.B1(n_209),
.B2(n_215),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_269),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_229),
.A2(n_208),
.B1(n_245),
.B2(n_231),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_246),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_272),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_240),
.C(n_242),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_233),
.C(n_249),
.Y(n_287)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_236),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_243),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_240),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_281),
.A2(n_283),
.B(n_286),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_266),
.B1(n_271),
.B2(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_260),
.C(n_256),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_267),
.B(n_234),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_236),
.Y(n_291)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_273),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_303),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_299),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_286),
.A2(n_262),
.B(n_270),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_298),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_260),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_268),
.C(n_265),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_264),
.C(n_269),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_301),
.B(n_305),
.Y(n_316)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_261),
.B(n_235),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_261),
.C(n_235),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_R g307 ( 
.A(n_293),
.B(n_296),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_304),
.B(n_305),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_303),
.A2(n_261),
.B1(n_282),
.B2(n_283),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_309),
.A2(n_311),
.B1(n_314),
.B2(n_315),
.Y(n_323)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_288),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_298),
.Y(n_318)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_300),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_295),
.A2(n_284),
.B1(n_277),
.B2(n_276),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_310),
.A2(n_284),
.B1(n_304),
.B2(n_301),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_320),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_306),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_312),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_308),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_315),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_308),
.Y(n_328)
);

OAI321xp33_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_285),
.A3(n_276),
.B1(n_280),
.B2(n_299),
.C(n_294),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_322),
.A2(n_313),
.B(n_312),
.Y(n_324)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_328),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.C(n_330),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_331),
.A2(n_323),
.B1(n_327),
.B2(n_324),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_309),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_335),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_280),
.B(n_306),
.C(n_318),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_235),
.Y(n_338)
);


endmodule