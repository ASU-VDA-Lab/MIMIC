module real_jpeg_1251_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_10;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_0),
.B(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_0),
.B(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

AO21x2_ASAP7_75t_L g11 ( 
.A1(n_3),
.A2(n_12),
.B(n_13),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_5),
.B(n_24),
.Y(n_23)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_5),
.B(n_24),
.Y(n_25)
);

A2O1A1O1Ixp25_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_9),
.B(n_17),
.C(n_18),
.D(n_27),
.Y(n_6)
);

O2A1O1Ixp33_ASAP7_75t_SL g27 ( 
.A1(n_7),
.A2(n_9),
.B(n_18),
.C(n_28),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_15),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_14),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);


endmodule