module real_jpeg_24638_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_48),
.B1(n_62),
.B2(n_63),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_247)
);

INVx8_ASAP7_75t_SL g61 ( 
.A(n_4),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_5),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_5),
.A2(n_28),
.B(n_43),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_5),
.B(n_91),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_5),
.A2(n_25),
.B1(n_180),
.B2(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_5),
.A2(n_62),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_5),
.B(n_78),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_154),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_154),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_6),
.A2(n_67),
.B1(n_70),
.B2(n_154),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_7),
.A2(n_52),
.B1(n_67),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_7),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_8),
.Y(n_88)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_10),
.A2(n_67),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_114),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_114),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_114),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_163),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_163),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_11),
.A2(n_77),
.B1(n_163),
.B2(n_275),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_85),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_13),
.A2(n_68),
.B1(n_85),
.B2(n_125),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_85),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_35),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_14),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_14),
.A2(n_35),
.B1(n_62),
.B2(n_63),
.Y(n_271)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_15),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_140),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_20),
.B(n_119),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.C(n_100),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_21),
.A2(n_80),
.B1(n_81),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_21),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_53),
.B2(n_79),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_22),
.A2(n_54),
.B(n_56),
.Y(n_138)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_24),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_24),
.A2(n_36),
.B1(n_54),
.B2(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_25),
.A2(n_106),
.B(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_25),
.A2(n_108),
.B1(n_171),
.B2(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_33),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_25),
.A2(n_211),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_26),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_26),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_26),
.A2(n_107),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_27),
.B(n_187),
.Y(n_186)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_31),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_31),
.A2(n_104),
.B(n_228),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_34),
.B(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_36),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_47),
.B(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_37),
.A2(n_46),
.B1(n_47),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_37),
.A2(n_46),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_37),
.A2(n_94),
.B(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_38),
.A2(n_95),
.B(n_96),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_38),
.A2(n_96),
.B1(n_153),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_38),
.A2(n_96),
.B1(n_162),
.B2(n_204),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_38),
.A2(n_50),
.B(n_95),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_46),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_40),
.A2(n_41),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_40),
.B(n_89),
.Y(n_209)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_SL g155 ( 
.A1(n_41),
.A2(n_45),
.B(n_151),
.C(n_156),
.Y(n_155)
);

OAI32xp33_ASAP7_75t_L g208 ( 
.A1(n_41),
.A2(n_62),
.A3(n_88),
.B1(n_200),
.B2(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_46),
.B(n_151),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_46),
.A2(n_97),
.B(n_110),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_51),
.Y(n_98)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_71),
.B(n_75),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_57),
.A2(n_112),
.B(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_57),
.A2(n_58),
.B1(n_112),
.B2(n_274),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_66),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_58),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_60),
.B1(n_67),
.B2(n_70),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_59),
.A2(n_63),
.A3(n_125),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_60),
.B(n_62),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_63),
.B1(n_88),
.B2(n_89),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_63),
.B(n_151),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_70),
.A2(n_151),
.B(n_243),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_72),
.B(n_78),
.Y(n_115)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_73),
.B(n_151),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_77),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_78),
.A2(n_127),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_78),
.A2(n_127),
.B1(n_260),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_93),
.B(n_99),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_93),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_87),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_86),
.A2(n_92),
.B(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_86),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_86),
.A2(n_91),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_86),
.A2(n_91),
.B1(n_222),
.B2(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_86),
.A2(n_256),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_87),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_87),
.B(n_271),
.Y(n_270)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_118),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_121),
.B1(n_136),
.B2(n_137),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_100),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.C(n_116),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_101),
.A2(n_102),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_103),
.B(n_109),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_105),
.B(n_173),
.Y(n_211)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_111),
.B(n_116),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_138),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_128),
.B2(n_135),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_134),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_131),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_133),
.A2(n_201),
.B(n_271),
.Y(n_287)
);

AOI311xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_296),
.A3(n_308),
.B(n_311),
.C(n_312),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_262),
.C(n_291),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_237),
.B(n_261),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_215),
.B(n_236),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_193),
.B(n_214),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_167),
.B(n_192),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_157),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_147),
.B(n_157),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_155),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_148),
.A2(n_149),
.B1(n_155),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_188),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_165),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_164),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_164),
.C(n_165),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_166),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_176),
.B(n_191),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_174),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_181),
.B(n_190),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_194),
.B(n_195),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_207),
.B1(n_212),
.B2(n_213),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_196)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_206),
.C(n_212),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_210),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_217),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_229),
.B2(n_230),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_232),
.C(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_225),
.C(n_226),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_239),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_253),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_240)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_241),
.B(n_252),
.C(n_253),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_242),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_248),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_245),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_247),
.Y(n_279)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_257),
.C(n_258),
.Y(n_276)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_263),
.A2(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_281),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_264),
.B(n_281),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_276),
.C(n_277),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_266),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_269),
.C(n_272),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_276),
.B(n_277),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_280),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_281),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_289),
.CI(n_290),
.CON(n_281),
.SN(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_288),
.Y(n_282)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_283),
.Y(n_288)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_293),
.Y(n_314)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

O2A1O1Ixp33_ASAP7_75t_SL g312 ( 
.A1(n_297),
.A2(n_309),
.B(n_313),
.C(n_316),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_305),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_305),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_298),
.B(n_310),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_301),
.CI(n_304),
.CON(n_298),
.SN(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);


endmodule