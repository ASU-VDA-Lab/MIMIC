module real_jpeg_16616_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_586;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_591),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_0),
.B(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_1),
.Y(n_437)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_2),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_2),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_185),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_3),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_3),
.A2(n_189),
.B1(n_245),
.B2(n_254),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_3),
.A2(n_189),
.B1(n_448),
.B2(n_451),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_3),
.A2(n_189),
.B1(n_507),
.B2(n_509),
.Y(n_506)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_196),
.A3(n_199),
.B1(n_202),
.B2(n_206),
.Y(n_195)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_4),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_4),
.A2(n_205),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

OAI32xp33_ASAP7_75t_L g342 ( 
.A1(n_4),
.A2(n_196),
.A3(n_199),
.B1(n_202),
.B2(n_206),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_4),
.B(n_24),
.Y(n_351)
);

OAI32xp33_ASAP7_75t_L g417 ( 
.A1(n_4),
.A2(n_418),
.A3(n_422),
.B1(n_426),
.B2(n_429),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_4),
.A2(n_196),
.B1(n_205),
.B2(n_456),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_4),
.B(n_70),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_4),
.B(n_544),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_4),
.B(n_318),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_5),
.A2(n_112),
.B1(n_113),
.B2(n_115),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_5),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_5),
.A2(n_115),
.B1(n_166),
.B2(n_169),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_5),
.A2(n_115),
.B1(n_237),
.B2(n_241),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_5),
.A2(n_115),
.B1(n_280),
.B2(n_307),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_6),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_6),
.A2(n_109),
.B1(n_225),
.B2(n_230),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_6),
.A2(n_109),
.B1(n_274),
.B2(n_279),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_6),
.A2(n_109),
.B1(n_374),
.B2(n_376),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_44),
.B1(n_62),
.B2(n_65),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_7),
.A2(n_44),
.B1(n_226),
.B2(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_7),
.A2(n_44),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_8),
.A2(n_34),
.B1(n_97),
.B2(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_8),
.A2(n_34),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_8),
.A2(n_34),
.B1(n_241),
.B2(n_300),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_9),
.Y(n_223)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_9),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_9),
.Y(n_298)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_10),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_10),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_11),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_11),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_11),
.A2(n_246),
.B1(n_346),
.B2(n_349),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_11),
.A2(n_246),
.B1(n_496),
.B2(n_501),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_11),
.A2(n_246),
.B1(n_535),
.B2(n_539),
.Y(n_534)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_12),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_15),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_15),
.Y(n_127)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_15),
.Y(n_219)
);

BUFx4f_ASAP7_75t_L g229 ( 
.A(n_15),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_16),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_17),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_156),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_154),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_22),
.B(n_57),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_23),
.A2(n_48),
.B(n_291),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

OR2x6_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_24),
.B(n_40),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_24),
.A2(n_47),
.B1(n_243),
.B2(n_248),
.Y(n_242)
);

AO22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_28),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_28),
.Y(n_193)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_28),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_30),
.Y(n_172)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_30),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_30),
.Y(n_432)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_33),
.Y(n_401)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_35),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_36),
.Y(n_254)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g247 ( 
.A(n_38),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_39),
.A2(n_105),
.B(n_110),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_47),
.Y(n_39)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_41),
.Y(n_245)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_42),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_48),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_48),
.A2(n_111),
.B(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_48),
.A2(n_110),
.B1(n_249),
.B2(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_48),
.A2(n_110),
.B1(n_244),
.B2(n_320),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_48),
.A2(n_151),
.B(n_401),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_51),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_52),
.Y(n_325)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_150),
.C(n_152),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_58),
.B(n_150),
.CI(n_152),
.CON(n_175),
.SN(n_175)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_103),
.C(n_116),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_59),
.A2(n_60),
.B1(n_116),
.B2(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AO21x1_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_68),
.B(n_94),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_61),
.B(n_70),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_61),
.Y(n_372)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_64),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_66),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_67),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_68),
.A2(n_70),
.B(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_68),
.A2(n_165),
.B(n_173),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_68),
.A2(n_94),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_68),
.A2(n_70),
.B1(n_165),
.B2(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_69),
.A2(n_96),
.B(n_174),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_69),
.A2(n_95),
.B1(n_184),
.B2(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_69),
.A2(n_95),
.B1(n_327),
.B2(n_345),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_69),
.A2(n_95),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_69),
.A2(n_95),
.B1(n_345),
.B2(n_455),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_81),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

AO22x2_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_76),
.Y(n_288)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_78),
.Y(n_285)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_89),
.B2(n_92),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_99),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_102),
.Y(n_377)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_162),
.C(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_117),
.B(n_164),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_129),
.B(n_141),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_118),
.B(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_118),
.A2(n_129),
.B1(n_492),
.B2(n_495),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_118),
.A2(n_129),
.B1(n_442),
.B2(n_495),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_119),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_119),
.B(n_142),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_120),
.Y(n_318)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_126),
.B2(n_128),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_123),
.Y(n_477)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_127),
.Y(n_241)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_127),
.Y(n_270)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_127),
.Y(n_542)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_128),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_129),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_129),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_129),
.A2(n_394),
.B(n_463),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_139),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_139),
.Y(n_452)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_140),
.Y(n_428)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_140),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_142),
.A2(n_305),
.B(n_317),
.Y(n_316)
);

OAI32xp33_ASAP7_75t_L g472 ( 
.A1(n_143),
.A2(n_473),
.A3(n_478),
.B1(n_482),
.B2(n_485),
.Y(n_472)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_148),
.Y(n_450)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21x1_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_176),
.B(n_589),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_175),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_159),
.B(n_175),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_160),
.A2(n_162),
.B1(n_569),
.B2(n_570),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_160),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_162),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_162),
.A2(n_570),
.B1(n_574),
.B2(n_575),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_163),
.B(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g593 ( 
.A(n_175),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_565),
.B(n_586),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_406),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_356),
.B(n_381),
.C(n_382),
.D(n_405),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_312),
.C(n_336),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_180),
.B(n_312),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_256),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_181),
.B(n_257),
.C(n_311),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_194),
.C(n_242),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_182),
.B(n_242),
.Y(n_314)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_188),
.Y(n_375)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_194),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_213),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_205),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_205),
.B(n_483),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_SL g492 ( 
.A1(n_205),
.A2(n_482),
.B(n_493),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_205),
.A2(n_215),
.B1(n_533),
.B2(n_534),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_213),
.B(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_224),
.B1(n_233),
.B2(n_236),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_214),
.A2(n_236),
.B(n_261),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_214),
.A2(n_261),
.B(n_439),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_214),
.A2(n_233),
.B1(n_520),
.B2(n_527),
.Y(n_519)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_215),
.B(n_267),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_215),
.A2(n_299),
.B(n_362),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_215),
.A2(n_506),
.B(n_513),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_215),
.A2(n_521),
.B1(n_534),
.B2(n_547),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_217),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_220),
.Y(n_533)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_222),
.Y(n_544)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_224),
.A2(n_302),
.B(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_229),
.Y(n_524)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_229),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_231),
.Y(n_539)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_232),
.Y(n_489)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_232),
.Y(n_512)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_255),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_251),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_251),
.A2(n_255),
.B1(n_328),
.B2(n_332),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_251),
.A2(n_255),
.B1(n_443),
.B2(n_445),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_251),
.A2(n_255),
.B1(n_522),
.B2(n_525),
.Y(n_521)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_293),
.B2(n_311),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_289),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_259),
.B(n_290),
.C(n_292),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_271),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_260),
.B(n_271),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_267),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_SL g353 ( 
.A(n_265),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_266),
.Y(n_365)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_283),
.Y(n_271)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_277),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_277),
.Y(n_503)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_278),
.Y(n_500)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g395 ( 
.A(n_283),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_303),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_294),
.B(n_303),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_302),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_295),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_299),
.Y(n_439)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g367 ( 
.A1(n_305),
.A2(n_306),
.B(n_317),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_305),
.A2(n_441),
.B1(n_447),
.B2(n_453),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_309),
.Y(n_444)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_310),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.C(n_335),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_335),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.C(n_326),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_326),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_318),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_319),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_330),
.Y(n_348)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_354),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_337),
.B(n_354),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.C(n_343),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_338),
.B(n_561),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_340),
.A2(n_341),
.B1(n_343),
.B2(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_343),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_350),
.C(n_352),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_344),
.B(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_351),
.B(n_352),
.Y(n_466)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_356),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_358),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_380),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_369),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_360),
.B(n_369),
.C(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_360)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_361),
.Y(n_368)
);

NOR2x1_ASAP7_75t_R g398 ( 
.A(n_361),
.B(n_367),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_361),
.A2(n_368),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

AOI21xp33_ASAP7_75t_L g578 ( 
.A1(n_368),
.A2(n_402),
.B(n_579),
.Y(n_578)
);

XNOR2x1_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_379),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_378),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_371),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_373),
.Y(n_392)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_378),
.B(n_379),
.C(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_380),
.Y(n_385)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR3xp33_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_408),
.C(n_411),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_386),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_387),
.B(n_397),
.C(n_404),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_390),
.A2(n_397),
.B1(n_403),
.B2(n_404),
.Y(n_389)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_390),
.Y(n_404)
);

OAI21xp33_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_393),
.B(n_396),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_391),
.B(n_393),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_396),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_396),
.A2(n_573),
.B1(n_576),
.B2(n_585),
.Y(n_584)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_397),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_398),
.Y(n_579)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_400),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_412),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_559),
.B(n_564),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_468),
.B(n_558),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_459),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_415),
.B(n_459),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_440),
.C(n_454),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_416),
.B(n_555),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_438),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_417),
.B(n_438),
.Y(n_461)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_440),
.B(n_454),
.Y(n_555)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_447),
.Y(n_463)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx8_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_464),
.B1(n_465),
.B2(n_467),
.Y(n_459)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_460),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_461),
.B(n_462),
.C(n_464),
.Y(n_563)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_469),
.A2(n_553),
.B(n_557),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_470),
.A2(n_517),
.B(n_552),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_504),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_471),
.B(n_504),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_490),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_472),
.A2(n_490),
.B1(n_491),
.B2(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_472),
.Y(n_529)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx8_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_514),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_505),
.B(n_515),
.C(n_516),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_506),
.Y(n_527)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_518),
.A2(n_530),
.B(n_551),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_528),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_519),
.B(n_528),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_524),
.Y(n_526)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_531),
.A2(n_545),
.B(n_550),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_540),
.Y(n_531)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_541),
.B(n_543),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_544),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_546),
.B(n_549),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_546),
.B(n_549),
.Y(n_550)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

NOR2xp67_ASAP7_75t_SL g553 ( 
.A(n_554),
.B(n_556),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_554),
.B(n_556),
.Y(n_557)
);

NOR2xp67_ASAP7_75t_SL g559 ( 
.A(n_560),
.B(n_563),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_560),
.B(n_563),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_566),
.B(n_580),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g586 ( 
.A1(n_566),
.A2(n_587),
.B(n_588),
.Y(n_586)
);

NOR2xp67_ASAP7_75t_SL g566 ( 
.A(n_567),
.B(n_571),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_567),
.B(n_571),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_576),
.C(n_577),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_573),
.Y(n_585)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_574),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_577),
.A2(n_578),
.B1(n_583),
.B2(n_584),
.Y(n_582)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_581),
.B(n_582),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_581),
.B(n_582),
.Y(n_587)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);


endmodule