module fake_jpeg_5927_n_50 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_50);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_50;

wire n_33;
wire n_45;
wire n_27;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_22),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_36),
.B1(n_37),
.B2(n_6),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

CKINVDCx11_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_17),
.B1(n_4),
.B2(n_5),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_1),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_28),
.B(n_1),
.C(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_31),
.C(n_10),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_11),
.B2(n_16),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_40),
.B(n_19),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_44),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

MAJx2_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_18),
.C(n_20),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_49),
.A2(n_21),
.B(n_24),
.Y(n_50)
);


endmodule