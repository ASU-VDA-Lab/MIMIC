module real_jpeg_20348_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_346, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_346;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_0),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_0),
.A2(n_23),
.B1(n_70),
.B2(n_71),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_0),
.A2(n_23),
.B1(n_52),
.B2(n_54),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_1),
.A2(n_52),
.B1(n_54),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_1),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_1),
.A2(n_70),
.B1(n_71),
.B2(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_94),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_1),
.A2(n_24),
.B1(n_26),
.B2(n_94),
.Y(n_212)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

A2O1A1O1Ixp25_ASAP7_75t_L g90 ( 
.A1(n_3),
.A2(n_54),
.B(n_66),
.C(n_91),
.D(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_3),
.B(n_51),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_3),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_3),
.A2(n_112),
.B(n_114),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_3),
.A2(n_32),
.B(n_48),
.C(n_148),
.D(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_32),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_3),
.B(n_36),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_33),
.B(n_192),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_129),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_4),
.A2(n_52),
.B1(n_54),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_4),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_4),
.A2(n_70),
.B1(n_71),
.B2(n_106),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_106),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_106),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_5),
.A2(n_70),
.B1(n_71),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_5),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_5),
.A2(n_52),
.B1(n_54),
.B2(n_160),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_160),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_5),
.A2(n_24),
.B1(n_26),
.B2(n_160),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_6),
.B(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_6),
.B(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_6),
.Y(n_123)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_6),
.A2(n_113),
.B1(n_159),
.B2(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_24),
.B1(n_26),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_7),
.A2(n_61),
.B1(n_70),
.B2(n_71),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_7),
.A2(n_52),
.B1(n_54),
.B2(n_61),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_61),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_9),
.A2(n_24),
.B1(n_26),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_9),
.A2(n_63),
.B1(n_70),
.B2(n_71),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_9),
.A2(n_52),
.B1(n_54),
.B2(n_63),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_63),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_10),
.A2(n_70),
.B1(n_71),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_10),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_52),
.B1(n_54),
.B2(n_111),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_111),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_111),
.Y(n_249)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_12),
.A2(n_24),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_12),
.A2(n_35),
.B1(n_52),
.B2(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_12),
.A2(n_35),
.B1(n_70),
.B2(n_71),
.Y(n_238)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_40),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_21),
.B(n_42),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_34),
.B2(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_22),
.A2(n_27),
.B1(n_36),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_24),
.A2(n_29),
.B(n_129),
.C(n_191),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_34),
.B(n_36),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_27),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_27),
.B(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_28),
.A2(n_31),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_28),
.A2(n_31),
.B1(n_220),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_28),
.A2(n_211),
.B(n_249),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_28),
.A2(n_31),
.B1(n_60),
.B2(n_293),
.Y(n_313)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_29),
.Y(n_192)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_31),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_31),
.A2(n_221),
.B(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_36),
.B(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_80),
.B(n_343),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_75),
.C(n_77),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_43),
.A2(n_44),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_58),
.C(n_64),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_45),
.A2(n_46),
.B1(n_64),
.B2(n_318),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_47),
.A2(n_56),
.B1(n_169),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_47),
.A2(n_206),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_51),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_48),
.B(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_48),
.A2(n_51),
.B1(n_246),
.B2(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_48),
.A2(n_51),
.B1(n_265),
.B2(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_49),
.B(n_54),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_50),
.A2(n_52),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_56),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_56),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_56),
.A2(n_170),
.B(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_58),
.A2(n_59),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_64),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_64),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_73),
.B(n_74),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_65),
.A2(n_73),
.B1(n_105),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_65),
.A2(n_146),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_65),
.A2(n_73),
.B1(n_203),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_65),
.A2(n_73),
.B1(n_231),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_65),
.A2(n_73),
.B1(n_240),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_66),
.A2(n_69),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_67),
.B(n_71),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_70),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_73),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_73),
.A2(n_107),
.B(n_203),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_74),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_339),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_75),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_336),
.B(n_342),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_309),
.A3(n_329),
.B1(n_334),
.B2(n_335),
.C(n_345),
.Y(n_81)
);

AOI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_257),
.A3(n_297),
.B1(n_303),
.B2(n_308),
.C(n_346),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_214),
.C(n_253),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_184),
.B(n_213),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_163),
.B(n_183),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_140),
.B(n_162),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_116),
.B(n_139),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_89),
.B(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_95),
.B1(n_96),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_92),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_104),
.C(n_109),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_112),
.B(n_114),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_112),
.A2(n_123),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_112),
.A2(n_123),
.B1(n_196),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_112),
.A2(n_123),
.B1(n_229),
.B2(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_112),
.A2(n_131),
.B(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_113),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_115),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_126),
.B(n_138),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_124),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_133),
.B(n_137),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_128),
.B(n_130),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_131),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_131),
.A2(n_132),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_142),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_153),
.B2(n_161),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_152),
.C(n_161),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_149),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_153),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_157),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_165),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_177),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_179),
.C(n_181),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_172),
.B2(n_176),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_173),
.C(n_174),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_172),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_175),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_178),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_185),
.B(n_186),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_200),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_187)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_188),
.B(n_199),
.C(n_200),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_194),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_197),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_208),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_207),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g304 ( 
.A1(n_215),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_233),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_216),
.B(n_233),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_227),
.C(n_232),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_217),
.B(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_232),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_230),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_251),
.B2(n_252),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_236),
.B(n_241),
.C(n_252),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_239),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_247),
.C(n_250),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_244),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_251),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_255),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_275),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_258),
.B(n_275),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_268),
.C(n_274),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_259),
.A2(n_260),
.B1(n_268),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_264),
.C(n_266),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_273),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_270),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_269),
.A2(n_288),
.B(n_292),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_271),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_271),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_272),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_301),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_295),
.B2(n_296),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_286),
.B2(n_287),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_287),
.C(n_296),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_283),
.B(n_285),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_283),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_284),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_285),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_285),
.A2(n_311),
.B1(n_320),
.B2(n_333),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_294),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_290),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_298),
.A2(n_304),
.B(n_307),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_322),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_322),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_320),
.C(n_321),
.Y(n_310)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_313),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_318),
.C(n_319),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_324),
.C(n_328),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_316),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_332),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_328),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_341),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_341),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_338),
.Y(n_340)
);


endmodule