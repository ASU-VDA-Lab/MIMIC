module fake_jpeg_25281_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

AND2x2_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_3),
.Y(n_7)
);

INVx3_ASAP7_75t_SL g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_0),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_0),
.C(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_15),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_8),
.A2(n_6),
.B1(n_13),
.B2(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_18),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_2),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_20),
.B1(n_6),
.B2(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_20),
.B(n_12),
.Y(n_28)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_14),
.C(n_9),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_16),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_21),
.C(n_26),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_R g32 ( 
.A(n_28),
.B(n_31),
.C(n_23),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_22),
.Y(n_35)
);

OAI22x1_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_11),
.B1(n_9),
.B2(n_12),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_33),
.B1(n_31),
.B2(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_21),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_35),
.C(n_33),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_26),
.C(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_26),
.C(n_21),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_23),
.B(n_1),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_23),
.C(n_24),
.Y(n_43)
);

OAI321xp33_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_44),
.A3(n_42),
.B1(n_11),
.B2(n_24),
.C(n_40),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_24),
.Y(n_46)
);


endmodule