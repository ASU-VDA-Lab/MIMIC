module fake_aes_12393_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x4_ASAP7_75t_L g13 ( .A(n_7), .B(n_10), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_5), .B(n_11), .Y(n_14) );
AOI22xp5_ASAP7_75t_L g15 ( .A1(n_0), .A2(n_2), .B1(n_9), .B2(n_6), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
NAND2xp33_ASAP7_75t_L g17 ( .A(n_1), .B(n_5), .Y(n_17) );
AND2x6_ASAP7_75t_L g18 ( .A(n_6), .B(n_12), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
AOI221xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_17), .B1(n_15), .B2(n_13), .C(n_14), .Y(n_21) );
A2O1A1Ixp33_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_18), .B(n_2), .C(n_3), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
AOI211xp5_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_21), .B(n_19), .C(n_24), .Y(n_26) );
AOI211xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_24), .B(n_18), .C(n_4), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_24), .B1(n_18), .B2(n_4), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
AOI322xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_1), .A3(n_3), .B1(n_7), .B2(n_8), .C1(n_18), .C2(n_26), .Y(n_30) );
endmodule