module fake_jpeg_21265_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_20),
.B1(n_19),
.B2(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_30),
.B1(n_23),
.B2(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_36),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_28),
.B1(n_29),
.B2(n_20),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_60),
.B1(n_30),
.B2(n_22),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_28),
.B1(n_29),
.B2(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_61),
.B(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_69),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_20),
.Y(n_65)
);

NAND2x1p5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_38),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_31),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_37),
.B1(n_28),
.B2(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_71),
.A2(n_73),
.B1(n_93),
.B2(n_106),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_77),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_37),
.B1(n_45),
.B2(n_42),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_SL g138 ( 
.A(n_74),
.B(n_105),
.C(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_75),
.B(n_87),
.Y(n_132)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_86),
.Y(n_119)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_45),
.B1(n_40),
.B2(n_39),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_83),
.A2(n_85),
.B1(n_90),
.B2(n_95),
.Y(n_147)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_45),
.B1(n_39),
.B2(n_22),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_18),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_33),
.B1(n_46),
.B2(n_18),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_56),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_109),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_16),
.B1(n_35),
.B2(n_25),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_68),
.B1(n_65),
.B2(n_63),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_96),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_57),
.A2(n_25),
.B1(n_35),
.B2(n_16),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_103),
.B1(n_24),
.B2(n_33),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_56),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_101),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_38),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_38),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_59),
.B(n_16),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_39),
.B1(n_44),
.B2(n_43),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_38),
.B1(n_23),
.B2(n_27),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_38),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_62),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g108 ( 
.A(n_59),
.B(n_34),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_59),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_18),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_110),
.B(n_18),
.Y(n_112)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_112),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_39),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_127),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_121),
.B1(n_141),
.B2(n_145),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_105),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_75),
.A2(n_38),
.B1(n_44),
.B2(n_43),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_26),
.B(n_23),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_130),
.B(n_100),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_88),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_135),
.B1(n_140),
.B2(n_143),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_82),
.B(n_111),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_109),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_0),
.B(n_1),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_27),
.B(n_26),
.C(n_24),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_146),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_78),
.A2(n_46),
.B1(n_33),
.B2(n_34),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_83),
.A2(n_34),
.B1(n_17),
.B2(n_0),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_99),
.A2(n_17),
.B1(n_8),
.B2(n_2),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_81),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_108),
.B(n_100),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_151),
.A2(n_152),
.B(n_161),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_121),
.Y(n_193)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_76),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_98),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_160),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_138),
.B(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_77),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_104),
.B(n_1),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_167),
.B(n_145),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_122),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_169),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_102),
.B(n_84),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_96),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_107),
.C(n_79),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_115),
.C(n_112),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_125),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_172),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_119),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_134),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_176),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_91),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_113),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_174),
.A2(n_147),
.B1(n_114),
.B2(n_123),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_197),
.B1(n_207),
.B2(n_175),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_126),
.B1(n_147),
.B2(n_141),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_184),
.A2(n_166),
.B1(n_154),
.B2(n_151),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_SL g185 ( 
.A1(n_171),
.A2(n_142),
.B(n_133),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_185),
.A2(n_190),
.B(n_211),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_162),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_123),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_193),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_200),
.C(n_206),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_146),
.B1(n_116),
.B2(n_106),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_115),
.C(n_131),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_161),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_171),
.A2(n_106),
.B1(n_137),
.B2(n_144),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_170),
.A2(n_144),
.B(n_92),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_210),
.A2(n_177),
.B(n_173),
.C(n_169),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_152),
.A2(n_4),
.B(n_5),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_212),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_205),
.Y(n_214)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_165),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_225),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_210),
.B(n_204),
.Y(n_253)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_201),
.B(n_155),
.Y(n_222)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_227),
.B1(n_228),
.B2(n_232),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_172),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_226),
.A2(n_186),
.B1(n_199),
.B2(n_89),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_203),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_180),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_229),
.B(n_231),
.C(n_235),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_167),
.C(n_153),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_194),
.C(n_202),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_158),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_191),
.B(n_156),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_191),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_184),
.A2(n_176),
.B1(n_175),
.B2(n_164),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_200),
.B(n_163),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_153),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_195),
.A2(n_167),
.B1(n_179),
.B2(n_178),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_202),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_242),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_195),
.B1(n_192),
.B2(n_182),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_239),
.A2(n_236),
.B1(n_252),
.B2(n_214),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_196),
.B(n_193),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_253),
.B(n_224),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_206),
.C(n_190),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_254),
.C(n_216),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_211),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_255),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_207),
.C(n_189),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_192),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_256),
.A2(n_214),
.B1(n_219),
.B2(n_215),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_217),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_261),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_237),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_240),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_267),
.B1(n_253),
.B2(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_266),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

NAND3xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_270),
.C(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_220),
.C(n_221),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_273),
.C(n_274),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_199),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_226),
.C(n_215),
.Y(n_274)
);

OAI321xp33_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_219),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_279),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_280),
.B(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_242),
.C(n_255),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_287),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_288),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_243),
.C(n_250),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_256),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_271),
.C(n_265),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_293),
.C(n_297),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_291),
.A2(n_276),
.B1(n_277),
.B2(n_284),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_265),
.C(n_269),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_260),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_261),
.C(n_219),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_279),
.C(n_262),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_305),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_306),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_SL g303 ( 
.A1(n_295),
.A2(n_288),
.B(n_280),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_304),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_286),
.B(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_311),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_293),
.C(n_294),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_294),
.C(n_302),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_9),
.C(n_11),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_313),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_316),
.B1(n_312),
.B2(n_310),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_11),
.B(n_13),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_14),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_321),
.B(n_14),
.Y(n_322)
);


endmodule