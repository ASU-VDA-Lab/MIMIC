module fake_jpeg_19164_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_44),
.Y(n_51)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_9),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx2_ASAP7_75t_R g96 ( 
.A(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_50),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_63),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_23),
.B1(n_28),
.B2(n_24),
.Y(n_87)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_56),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_29),
.B1(n_27),
.B2(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_22),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_43),
.B(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_24),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_64),
.B(n_69),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_32),
.B1(n_42),
.B2(n_41),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_65),
.A2(n_77),
.B1(n_88),
.B2(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_75),
.Y(n_135)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_73),
.Y(n_113)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_59),
.B1(n_62),
.B2(n_47),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_79),
.B(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_82),
.Y(n_125)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_84),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_46),
.B(n_61),
.C(n_50),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_17),
.B(n_34),
.C(n_0),
.Y(n_133)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_103),
.B1(n_25),
.B2(n_41),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_26),
.B1(n_28),
.B2(n_23),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_92),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_43),
.B(n_38),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_26),
.B1(n_21),
.B2(n_27),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_16),
.B1(n_35),
.B2(n_30),
.Y(n_120)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_100),
.Y(n_131)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_99),
.Y(n_105)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_16),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_29),
.Y(n_102)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_102),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g103 ( 
.A1(n_46),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_56),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_25),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_110),
.A2(n_120),
.B1(n_1),
.B2(n_15),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_85),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_38),
.B1(n_35),
.B2(n_30),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_72),
.B1(n_100),
.B2(n_95),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_78),
.A2(n_16),
.B(n_34),
.C(n_20),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_124),
.B(n_130),
.C(n_89),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_85),
.A2(n_0),
.B(n_1),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_133),
.B(n_116),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_85),
.B(n_79),
.C(n_96),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g130 ( 
.A1(n_67),
.A2(n_34),
.A3(n_20),
.B1(n_30),
.B2(n_17),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_68),
.B(n_17),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_92),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_141),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_74),
.B1(n_72),
.B2(n_97),
.Y(n_138)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_145),
.B(n_149),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_148),
.Y(n_168)
);

INVx6_ASAP7_75t_SL g143 ( 
.A(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_144),
.Y(n_176)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_66),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_133),
.B1(n_110),
.B2(n_148),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_77),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_65),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_98),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_11),
.CI(n_2),
.CON(n_150),
.SN(n_150)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_81),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_122),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_10),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_105),
.B(n_1),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_162),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_114),
.B(n_10),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_11),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_107),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_159)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_8),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_115),
.B(n_8),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_163),
.A2(n_164),
.B1(n_131),
.B2(n_107),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_112),
.C(n_124),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_172),
.C(n_175),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_106),
.C(n_127),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_127),
.C(n_120),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_178),
.B(n_182),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_144),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_115),
.C(n_117),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_126),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_133),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_150),
.B(n_134),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_118),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_156),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_190),
.A2(n_125),
.B1(n_126),
.B2(n_108),
.Y(n_222)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_146),
.B1(n_151),
.B2(n_155),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_109),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_193),
.B(n_164),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_109),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_177),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_199),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_180),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_198),
.B(n_206),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_145),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_208),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_207),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_166),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_180),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_170),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_212),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_150),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_188),
.B(n_154),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_215),
.B(n_224),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_163),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_223),
.C(n_169),
.Y(n_229)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_174),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_167),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_111),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_189),
.B(n_167),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_226),
.A2(n_243),
.B1(n_212),
.B2(n_201),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_239),
.Y(n_254)
);

FAx1_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_190),
.CI(n_189),
.CON(n_232),
.SN(n_232)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_232),
.A2(n_186),
.B(n_208),
.C(n_195),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_200),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_241),
.Y(n_250)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_166),
.C(n_191),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_220),
.C(n_217),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_211),
.A2(n_171),
.B1(n_173),
.B2(n_196),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_218),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_246),
.B(n_248),
.Y(n_266)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_205),
.CI(n_223),
.CON(n_247),
.SN(n_247)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_252),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_257),
.C(n_259),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_217),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_228),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_222),
.B1(n_216),
.B2(n_225),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_179),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_258),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_203),
.C(n_209),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_194),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_203),
.C(n_210),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_210),
.C(n_211),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_261),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_240),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_230),
.A2(n_185),
.B1(n_214),
.B2(n_181),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_264),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_230),
.B(n_228),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_225),
.A2(n_173),
.B1(n_171),
.B2(n_208),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_242),
.B1(n_244),
.B2(n_256),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_265),
.A2(n_260),
.B1(n_263),
.B2(n_232),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_267),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_269),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_244),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_275),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_263),
.A2(n_234),
.B(n_231),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_235),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_263),
.A2(n_231),
.B(n_232),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_251),
.B(n_174),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_249),
.C(n_259),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_284),
.C(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_254),
.C(n_247),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_111),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_265),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_280),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_295),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_273),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_297),
.B(n_298),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_279),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_267),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_294),
.A2(n_274),
.B1(n_290),
.B2(n_271),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_292),
.A2(n_284),
.B(n_286),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_302),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_286),
.B(n_287),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_303),
.A2(n_125),
.B(n_3),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_307),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_301),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_305),
.B(n_300),
.C(n_304),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_309),
.Y(n_311)
);

OAI321xp33_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_12),
.A3(n_4),
.B1(n_6),
.B2(n_8),
.C(n_15),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_6),
.Y(n_313)
);


endmodule