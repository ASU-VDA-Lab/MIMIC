module fake_jpeg_24735_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_45),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_19),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_0),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_32),
.B(n_1),
.Y(n_64)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_28),
.A2(n_22),
.B1(n_33),
.B2(n_36),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_18),
.B1(n_33),
.B2(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_55),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_18),
.B1(n_36),
.B2(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_37),
.B1(n_28),
.B2(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_38),
.B1(n_40),
.B2(n_17),
.Y(n_84)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_46),
.Y(n_80)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_70),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_50),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_75),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_46),
.B1(n_30),
.B2(n_35),
.Y(n_115)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_79),
.Y(n_129)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_90),
.CON(n_106),
.SN(n_106)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_98),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_45),
.B1(n_48),
.B2(n_37),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_82),
.A2(n_30),
.B1(n_21),
.B2(n_35),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_97),
.B1(n_39),
.B2(n_56),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_17),
.B1(n_24),
.B2(n_25),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_86),
.B(n_87),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_17),
.B1(n_25),
.B2(n_40),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_94),
.Y(n_124)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_54),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_59),
.A2(n_17),
.B1(n_38),
.B2(n_19),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_55),
.B(n_29),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_100),
.B(n_20),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_39),
.B1(n_47),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_104),
.B1(n_118),
.B2(n_71),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_102),
.A2(n_115),
.B1(n_130),
.B2(n_93),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_47),
.B1(n_57),
.B2(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_46),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_116),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_46),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_32),
.Y(n_157)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_43),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_45),
.B1(n_43),
.B2(n_21),
.Y(n_118)
);

INVxp67_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_78),
.B(n_32),
.Y(n_143)
);

CKINVDCx12_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_69),
.B(n_45),
.C(n_43),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_96),
.C(n_73),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_92),
.B(n_75),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_143),
.B(n_149),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_139),
.B1(n_127),
.B2(n_124),
.Y(n_174)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_77),
.B1(n_95),
.B2(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_61),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_152),
.Y(n_178)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_20),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_0),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_150),
.A2(n_155),
.B1(n_156),
.B2(n_99),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_127),
.B1(n_124),
.B2(n_104),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_107),
.B(n_67),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_154),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_32),
.B(n_1),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_99),
.A2(n_110),
.B1(n_114),
.B2(n_79),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_118),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_102),
.B1(n_101),
.B2(n_130),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_172),
.B1(n_135),
.B2(n_134),
.Y(n_200)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_177),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_160),
.Y(n_209)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_171),
.B1(n_173),
.B2(n_187),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_154),
.A2(n_109),
.B1(n_118),
.B2(n_100),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_SL g197 ( 
.A(n_164),
.B(n_10),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_123),
.B(n_118),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_168),
.B(n_174),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_132),
.B1(n_138),
.B2(n_155),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_126),
.B1(n_127),
.B2(n_124),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_181),
.B1(n_184),
.B2(n_135),
.Y(n_204)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_179),
.A2(n_23),
.B(n_3),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_136),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_180),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_107),
.B1(n_103),
.B2(n_117),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_21),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_103),
.B1(n_26),
.B2(n_27),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_188),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_26),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_203),
.Y(n_237)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_149),
.B(n_141),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_195),
.A2(n_210),
.B(n_2),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_23),
.Y(n_226)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_204),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_200),
.A2(n_208),
.B1(n_188),
.B2(n_185),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_134),
.C(n_141),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_206),
.C(n_220),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_142),
.Y(n_205)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_142),
.C(n_150),
.Y(n_206)
);

AOI22x1_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_88),
.B1(n_112),
.B2(n_128),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_23),
.B(n_3),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_137),
.B1(n_140),
.B2(n_34),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_0),
.Y(n_210)
);

OAI21x1_ASAP7_75t_SL g212 ( 
.A1(n_174),
.A2(n_30),
.B(n_23),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_167),
.B1(n_177),
.B2(n_23),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_216),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_164),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_207),
.B1(n_204),
.B2(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_113),
.Y(n_215)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_159),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_158),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_165),
.B(n_170),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_221),
.A2(n_224),
.B(n_195),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_241),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_211),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_175),
.B(n_165),
.C(n_181),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_238),
.C(n_243),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_226),
.A2(n_231),
.B1(n_191),
.B2(n_189),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_158),
.B1(n_180),
.B2(n_183),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_233),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_203),
.B1(n_213),
.B2(n_214),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_192),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_230),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_158),
.Y(n_234)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_205),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_236),
.A2(n_194),
.B1(n_218),
.B2(n_199),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_158),
.C(n_167),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_242),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_186),
.C(n_4),
.Y(n_243)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_266),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_219),
.B1(n_189),
.B2(n_194),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_237),
.B(n_190),
.Y(n_253)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_259),
.B1(n_260),
.B2(n_263),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_243),
.B(n_198),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_256),
.B(n_258),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_244),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_261),
.A2(n_252),
.B1(n_267),
.B2(n_251),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_221),
.Y(n_280)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_227),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_210),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_246),
.C(n_240),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_271),
.C(n_276),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_233),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_273),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_265),
.C(n_225),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_228),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_242),
.C(n_222),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_235),
.B1(n_251),
.B2(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_277),
.A2(n_241),
.B1(n_210),
.B2(n_12),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_223),
.C(n_191),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_284),
.C(n_285),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_241),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_250),
.A2(n_224),
.B1(n_198),
.B2(n_231),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_282),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_208),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_16),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_226),
.C(n_195),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_260),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_273),
.B(n_247),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_15),
.C(n_14),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_290),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_252),
.B1(n_261),
.B2(n_249),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_289),
.A2(n_293),
.B1(n_299),
.B2(n_284),
.Y(n_301)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_292),
.B(n_296),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_276),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_16),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_271),
.C(n_269),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_305),
.C(n_309),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_307),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_285),
.C(n_278),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_286),
.B(n_300),
.CI(n_290),
.CON(n_307),
.SN(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_287),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_308),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_2),
.C(n_4),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_311),
.C(n_5),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_5),
.C(n_6),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_294),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_300),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_313),
.B(n_316),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_291),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_307),
.B(n_315),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_320),
.B1(n_311),
.B2(n_310),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_11),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_13),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_323),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_319),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_303),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_327),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_317),
.A2(n_305),
.B(n_15),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_326),
.A2(n_5),
.B(n_6),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_314),
.A2(n_15),
.B1(n_6),
.B2(n_7),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_331),
.B(n_332),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_334),
.B(n_325),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_330),
.C(n_328),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_6),
.B(n_7),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_7),
.B(n_8),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_8),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_8),
.B(n_320),
.Y(n_341)
);


endmodule