module fake_jpeg_1283_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_5),
.B(n_2),
.Y(n_6)
);

INVx11_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_14),
.Y(n_17)
);

INVx3_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

AND2x6_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_0),
.Y(n_16)
);

NAND2xp33_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_6),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_6),
.C(n_14),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_10),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_14),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_10),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_13),
.C(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_22),
.B1(n_13),
.B2(n_15),
.Y(n_27)
);

AOI322xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_12),
.A3(n_8),
.B1(n_11),
.B2(n_7),
.C1(n_2),
.C2(n_4),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_30),
.B(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_1),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_11),
.B1(n_7),
.B2(n_12),
.Y(n_33)
);


endmodule