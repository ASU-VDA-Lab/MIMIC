module fake_netlist_6_574_n_37 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_37);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;

output n_37;

wire n_16;
wire n_34;
wire n_9;
wire n_8;
wire n_18;
wire n_10;
wire n_24;
wire n_21;
wire n_15;
wire n_33;
wire n_27;
wire n_14;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_13;
wire n_35;
wire n_11;
wire n_28;
wire n_23;
wire n_17;
wire n_12;
wire n_20;
wire n_30;
wire n_19;
wire n_29;
wire n_31;
wire n_25;

INVx2_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

CKINVDCx5p33_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx5p33_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx5p33_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_R g15 ( 
.A(n_11),
.B(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_12),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_2),
.B(n_3),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_10),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_19),
.Y(n_28)
);

NOR2x1_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_18),
.Y(n_29)
);

XNOR2x2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_10),
.Y(n_30)
);

OAI322xp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_28),
.A3(n_26),
.B1(n_21),
.B2(n_17),
.C1(n_16),
.C2(n_4),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_17),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_16),
.C(n_15),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_R g34 ( 
.A(n_32),
.B(n_31),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_34),
.B1(n_2),
.B2(n_4),
.Y(n_37)
);


endmodule