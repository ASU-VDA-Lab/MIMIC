module real_aes_6377_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g494 ( .A(n_0), .Y(n_494) );
AOI22xp5_ASAP7_75t_SL g267 ( .A1(n_1), .A2(n_182), .B1(n_268), .B2(n_272), .Y(n_267) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_2), .A2(n_12), .B1(n_299), .B2(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g359 ( .A(n_3), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_4), .A2(n_92), .B1(n_287), .B2(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_5), .A2(n_47), .B1(n_300), .B2(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_6), .A2(n_13), .B1(n_253), .B2(n_560), .Y(n_702) );
INVx1_ASAP7_75t_L g477 ( .A(n_7), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_8), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_9), .A2(n_108), .B1(n_412), .B2(n_565), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_10), .A2(n_121), .B1(n_414), .B2(n_532), .Y(n_531) );
AOI222xp33_ASAP7_75t_L g638 ( .A1(n_11), .A2(n_105), .B1(n_170), .B2(n_287), .C1(n_351), .C2(n_449), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_14), .A2(n_90), .B1(n_326), .B2(n_328), .C(n_329), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g282 ( .A(n_15), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_16), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_17), .A2(n_59), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_18), .A2(n_138), .B1(n_560), .B2(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g487 ( .A(n_19), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_20), .Y(n_393) );
AO22x2_ASAP7_75t_L g242 ( .A1(n_21), .A2(n_70), .B1(n_243), .B2(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g656 ( .A(n_21), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_22), .A2(n_132), .B1(n_579), .B2(n_581), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_23), .A2(n_157), .B1(n_412), .B2(n_419), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_24), .A2(n_221), .B1(n_272), .B2(n_371), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g295 ( .A1(n_25), .A2(n_167), .B1(n_296), .B2(n_299), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_26), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_27), .B(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_28), .A2(n_130), .B1(n_264), .B2(n_275), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_29), .A2(n_202), .B1(n_253), .B2(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g483 ( .A(n_30), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_31), .B(n_517), .Y(n_636) );
AOI222xp33_ASAP7_75t_L g703 ( .A1(n_32), .A2(n_114), .B1(n_163), .B2(n_351), .C1(n_552), .C2(n_704), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_33), .A2(n_425), .B1(n_459), .B2(n_460), .Y(n_424) );
INVx1_ASAP7_75t_L g459 ( .A(n_33), .Y(n_459) );
INVx1_ASAP7_75t_L g522 ( .A(n_34), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g671 ( .A1(n_35), .A2(n_144), .B1(n_300), .B2(n_619), .Y(n_671) );
AO22x2_ASAP7_75t_L g246 ( .A1(n_36), .A2(n_74), .B1(n_243), .B2(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g657 ( .A(n_36), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_37), .A2(n_131), .B1(n_268), .B2(n_371), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_38), .A2(n_211), .B1(n_304), .B2(n_340), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_39), .A2(n_133), .B1(n_275), .B2(n_277), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_40), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_41), .A2(n_73), .B1(n_335), .B2(n_432), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_42), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_43), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_44), .A2(n_192), .B1(n_277), .B2(n_419), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_45), .A2(n_117), .B1(n_300), .B2(n_388), .Y(n_699) );
AOI222xp33_ASAP7_75t_L g623 ( .A1(n_46), .A2(n_154), .B1(n_206), .B2(n_296), .C1(n_552), .C2(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_48), .Y(n_428) );
AOI22xp5_ASAP7_75t_SL g259 ( .A1(n_49), .A2(n_127), .B1(n_260), .B2(n_264), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_50), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_51), .A2(n_80), .B1(n_339), .B2(n_340), .C(n_341), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_52), .A2(n_314), .B1(n_315), .B2(n_356), .Y(n_313) );
INVx1_ASAP7_75t_L g356 ( .A(n_52), .Y(n_356) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_53), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_54), .A2(n_217), .B1(n_364), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_55), .A2(n_123), .B1(n_299), .B2(n_388), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_56), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_57), .A2(n_149), .B1(n_277), .B2(n_414), .Y(n_621) );
AOI22xp33_ASAP7_75t_SL g673 ( .A1(n_58), .A2(n_159), .B1(n_414), .B2(n_562), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_60), .Y(n_377) );
AOI22xp5_ASAP7_75t_SL g235 ( .A1(n_61), .A2(n_115), .B1(n_236), .B2(n_253), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_62), .A2(n_174), .B1(n_304), .B2(n_307), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_63), .Y(n_548) );
AO22x2_ASAP7_75t_L g540 ( .A1(n_64), .A2(n_541), .B1(n_566), .B2(n_567), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_64), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_65), .A2(n_180), .B1(n_433), .B2(n_560), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_66), .Y(n_443) );
AOI22xp5_ASAP7_75t_SL g362 ( .A1(n_67), .A2(n_120), .B1(n_253), .B2(n_275), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_68), .A2(n_122), .B1(n_369), .B2(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g533 ( .A(n_69), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g350 ( .A1(n_71), .A2(n_91), .B1(n_112), .B2(n_351), .C1(n_352), .C2(n_354), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_72), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_75), .A2(n_164), .B1(n_278), .B2(n_336), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_76), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_77), .Y(n_450) );
AND2x2_ASAP7_75t_L g229 ( .A(n_78), .B(n_230), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_79), .A2(n_160), .B1(n_414), .B2(n_415), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_81), .A2(n_110), .B1(n_328), .B2(n_419), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_82), .B(n_505), .Y(n_504) );
AOI22xp5_ASAP7_75t_SL g367 ( .A1(n_83), .A2(n_184), .B1(n_368), .B2(n_369), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_84), .A2(n_152), .B1(n_387), .B2(n_388), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_85), .A2(n_101), .B1(n_369), .B2(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g226 ( .A(n_86), .Y(n_226) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_87), .A2(n_137), .B1(n_419), .B2(n_420), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_88), .A2(n_119), .B1(n_288), .B2(n_296), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_89), .B(n_340), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_93), .A2(n_134), .B1(n_618), .B2(n_619), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_94), .A2(n_187), .B1(n_322), .B2(n_565), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_95), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_96), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_97), .A2(n_140), .B1(n_265), .B2(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g496 ( .A(n_98), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_99), .A2(n_201), .B1(n_601), .B2(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g509 ( .A(n_100), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_102), .Y(n_446) );
INVx1_ASAP7_75t_L g333 ( .A(n_103), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_104), .A2(n_473), .B1(n_510), .B2(n_511), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g510 ( .A(n_104), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_106), .A2(n_139), .B1(n_364), .B2(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_107), .A2(n_189), .B1(n_597), .B2(n_599), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_109), .A2(n_181), .B1(n_336), .B2(n_420), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g317 ( .A1(n_111), .A2(n_158), .B1(n_236), .B2(n_318), .C(n_320), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_113), .A2(n_148), .B1(n_287), .B2(n_292), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_116), .Y(n_639) );
INVx2_ASAP7_75t_L g230 ( .A(n_118), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_124), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_125), .A2(n_166), .B1(n_335), .B2(n_594), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_126), .A2(n_190), .B1(n_489), .B2(n_491), .Y(n_488) );
AND2x6_ASAP7_75t_L g225 ( .A(n_128), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_128), .Y(n_650) );
AO22x2_ASAP7_75t_L g250 ( .A1(n_129), .A2(n_178), .B1(n_243), .B2(n_247), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_135), .A2(n_198), .B1(n_364), .B2(n_415), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_136), .A2(n_161), .B1(n_236), .B2(n_527), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_141), .Y(n_385) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_142), .A2(n_205), .B1(n_275), .B2(n_415), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_143), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_145), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_146), .Y(n_422) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_147), .A2(n_223), .B(n_231), .C(n_658), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_150), .A2(n_204), .B1(n_564), .B2(n_565), .Y(n_563) );
AO22x1_ASAP7_75t_L g320 ( .A1(n_151), .A2(n_176), .B1(n_321), .B2(n_323), .Y(n_320) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_153), .A2(n_195), .B1(n_369), .B2(n_412), .Y(n_677) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_155), .A2(n_193), .B1(n_243), .B2(n_244), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_156), .A2(n_196), .B1(n_502), .B2(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_162), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_165), .A2(n_218), .B1(n_355), .B2(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_168), .B(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_SL g678 ( .A1(n_169), .A2(n_197), .B1(n_236), .B2(n_264), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_171), .A2(n_194), .B1(n_336), .B2(n_433), .Y(n_622) );
INVx1_ASAP7_75t_L g503 ( .A(n_172), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_173), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_175), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_177), .A2(n_183), .B1(n_322), .B2(n_529), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_178), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_179), .B(n_340), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_185), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_186), .A2(n_203), .B1(n_340), .B2(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g507 ( .A(n_188), .Y(n_507) );
INVx1_ASAP7_75t_L g330 ( .A(n_191), .Y(n_330) );
INVx1_ASAP7_75t_L g653 ( .A(n_193), .Y(n_653) );
INVx1_ASAP7_75t_L g480 ( .A(n_199), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_200), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_207), .B(n_339), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_208), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_209), .Y(n_344) );
INVx1_ASAP7_75t_L g243 ( .A(n_210), .Y(n_243) );
INVx1_ASAP7_75t_L g245 ( .A(n_210), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_212), .Y(n_686) );
XOR2xp5_ASAP7_75t_L g659 ( .A(n_213), .B(n_660), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_214), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_215), .Y(n_454) );
INVx1_ASAP7_75t_L g500 ( .A(n_216), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_219), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_220), .A2(n_571), .B1(n_605), .B2(n_606), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_220), .Y(n_605) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_226), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_227), .A2(n_648), .B(n_685), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_466), .B1(n_643), .B2(n_644), .C(n_645), .Y(n_231) );
INVx1_ASAP7_75t_L g643 ( .A(n_232), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_309), .B1(n_464), .B2(n_465), .Y(n_232) );
INVx2_ASAP7_75t_L g464 ( .A(n_233), .Y(n_464) );
XOR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_308), .Y(n_233) );
NAND4xp75_ASAP7_75t_SL g234 ( .A(n_235), .B(n_259), .C(n_266), .D(n_280), .Y(n_234) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx4_ASAP7_75t_L g368 ( .A(n_237), .Y(n_368) );
OAI221xp5_ASAP7_75t_SL g427 ( .A1(n_237), .A2(n_428), .B1(n_429), .B2(n_430), .C(n_431), .Y(n_427) );
INVx2_ASAP7_75t_SL g479 ( .A(n_237), .Y(n_479) );
INVx11_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx11_ASAP7_75t_L g416 ( .A(n_238), .Y(n_416) );
AND2x6_ASAP7_75t_L g238 ( .A(n_239), .B(n_248), .Y(n_238) );
AND2x4_ASAP7_75t_L g306 ( .A(n_239), .B(n_279), .Y(n_306) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g383 ( .A(n_240), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_246), .Y(n_240) );
AND2x2_ASAP7_75t_L g258 ( .A(n_241), .B(n_246), .Y(n_258) );
AND2x2_ASAP7_75t_L g262 ( .A(n_241), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g285 ( .A(n_242), .B(n_246), .Y(n_285) );
AND2x2_ASAP7_75t_L g291 ( .A(n_242), .B(n_250), .Y(n_291) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g247 ( .A(n_245), .Y(n_247) );
INVx2_ASAP7_75t_L g263 ( .A(n_246), .Y(n_263) );
INVx1_ASAP7_75t_L g302 ( .A(n_246), .Y(n_302) );
AND2x2_ASAP7_75t_L g261 ( .A(n_248), .B(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g265 ( .A(n_248), .B(n_258), .Y(n_265) );
AND2x6_ASAP7_75t_L g284 ( .A(n_248), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
AND2x2_ASAP7_75t_L g279 ( .A(n_249), .B(n_252), .Y(n_279) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g256 ( .A(n_250), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_250), .B(n_252), .Y(n_271) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g257 ( .A(n_252), .Y(n_257) );
INVx1_ASAP7_75t_L g290 ( .A(n_252), .Y(n_290) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx5_ASAP7_75t_L g420 ( .A(n_254), .Y(n_420) );
INVx2_ASAP7_75t_L g433 ( .A(n_254), .Y(n_433) );
BUFx3_ASAP7_75t_L g490 ( .A(n_254), .Y(n_490) );
INVx1_ASAP7_75t_L g675 ( .A(n_254), .Y(n_675) );
INVx8_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_258), .Y(n_255) );
AND2x2_ASAP7_75t_L g276 ( .A(n_256), .B(n_262), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_256), .B(n_258), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_256), .B(n_262), .Y(n_486) );
INVx1_ASAP7_75t_L g293 ( .A(n_257), .Y(n_293) );
AND2x6_ASAP7_75t_L g307 ( .A(n_258), .B(n_279), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g376 ( .A(n_258), .B(n_279), .Y(n_376) );
BUFx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
INVx2_ASAP7_75t_L g365 ( .A(n_261), .Y(n_365) );
AND2x4_ASAP7_75t_L g269 ( .A(n_262), .B(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g278 ( .A(n_262), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g273 ( .A(n_263), .Y(n_273) );
AND2x2_ASAP7_75t_L g298 ( .A(n_263), .B(n_290), .Y(n_298) );
BUFx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx6_ASAP7_75t_L g327 ( .A(n_265), .Y(n_327) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_274), .Y(n_266) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx3_ASAP7_75t_L g324 ( .A(n_269), .Y(n_324) );
BUFx3_ASAP7_75t_L g369 ( .A(n_269), .Y(n_369) );
BUFx2_ASAP7_75t_L g532 ( .A(n_269), .Y(n_532) );
BUFx3_ASAP7_75t_L g565 ( .A(n_269), .Y(n_565) );
AND2x2_ASAP7_75t_L g272 ( .A(n_270), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OR2x6_ASAP7_75t_L g337 ( .A(n_271), .B(n_302), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_273), .B(n_291), .Y(n_343) );
BUFx2_ASAP7_75t_L g328 ( .A(n_275), .Y(n_328) );
BUFx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx3_ASAP7_75t_L g412 ( .A(n_276), .Y(n_412) );
BUFx3_ASAP7_75t_L g603 ( .A(n_276), .Y(n_603) );
BUFx3_ASAP7_75t_L g695 ( .A(n_276), .Y(n_695) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_277), .Y(n_438) );
BUFx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx3_ASAP7_75t_L g322 ( .A(n_278), .Y(n_322) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_278), .Y(n_371) );
BUFx3_ASAP7_75t_L g562 ( .A(n_278), .Y(n_562) );
INVx2_ASAP7_75t_L g592 ( .A(n_278), .Y(n_592) );
INVx1_ASAP7_75t_L g384 ( .A(n_279), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_294), .Y(n_280) );
OAI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_286), .Y(n_281) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_284), .Y(n_351) );
INVx4_ASAP7_75t_L g390 ( .A(n_284), .Y(n_390) );
INVx2_ASAP7_75t_L g402 ( .A(n_284), .Y(n_402) );
BUFx3_ASAP7_75t_L g550 ( .A(n_284), .Y(n_550) );
AND2x4_ASAP7_75t_L g292 ( .A(n_285), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g348 ( .A(n_285), .Y(n_348) );
INVx2_ASAP7_75t_L g553 ( .A(n_287), .Y(n_553) );
BUFx12f_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_288), .Y(n_355) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_288), .Y(n_387) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g297 ( .A(n_291), .B(n_298), .Y(n_297) );
AND2x4_ASAP7_75t_L g300 ( .A(n_291), .B(n_301), .Y(n_300) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_292), .Y(n_388) );
BUFx2_ASAP7_75t_SL g404 ( .A(n_292), .Y(n_404) );
BUFx2_ASAP7_75t_SL g524 ( .A(n_292), .Y(n_524) );
BUFx3_ASAP7_75t_L g619 ( .A(n_292), .Y(n_619) );
INVx1_ASAP7_75t_L g349 ( .A(n_293), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_303), .Y(n_294) );
INVx4_ASAP7_75t_L g353 ( .A(n_296), .Y(n_353) );
INVx2_ASAP7_75t_L g392 ( .A(n_296), .Y(n_392) );
BUFx2_ASAP7_75t_L g704 ( .A(n_296), .Y(n_704) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx4f_ASAP7_75t_SL g407 ( .A(n_297), .Y(n_407) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_297), .Y(n_449) );
BUFx2_ASAP7_75t_L g502 ( .A(n_297), .Y(n_502) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_297), .Y(n_520) );
BUFx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g580 ( .A(n_300), .Y(n_580) );
BUFx2_ASAP7_75t_L g618 ( .A(n_300), .Y(n_618) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_304), .Y(n_339) );
INVx5_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g517 ( .A(n_305), .Y(n_517) );
INVx2_ASAP7_75t_L g616 ( .A(n_305), .Y(n_616) );
INVx2_ASAP7_75t_L g670 ( .A(n_305), .Y(n_670) );
INVx4_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx4f_ASAP7_75t_L g340 ( .A(n_307), .Y(n_340) );
INVx1_ASAP7_75t_L g465 ( .A(n_309), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_396), .B2(n_463), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_357), .B1(n_394), .B2(n_395), .Y(n_311) );
INVx1_ASAP7_75t_L g394 ( .A(n_312), .Y(n_394) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND4x1_ASAP7_75t_L g316 ( .A(n_317), .B(n_325), .C(n_338), .D(n_350), .Y(n_316) );
INVx1_ASAP7_75t_SL g476 ( .A(n_318), .Y(n_476) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx3_ASAP7_75t_L g435 ( .A(n_319), .Y(n_435) );
BUFx3_ASAP7_75t_L g590 ( .A(n_319), .Y(n_590) );
BUFx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g429 ( .A(n_324), .Y(n_429) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g419 ( .A(n_327), .Y(n_419) );
OAI221xp5_ASAP7_75t_SL g482 ( .A1(n_327), .A2(n_483), .B1(n_484), .B2(n_487), .C(n_488), .Y(n_482) );
INVx2_ASAP7_75t_L g527 ( .A(n_327), .Y(n_527) );
INVx2_ASAP7_75t_L g599 ( .A(n_327), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B1(n_333), .B2(n_334), .Y(n_329) );
BUFx2_ASAP7_75t_R g331 ( .A(n_332), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_335), .Y(n_334) );
BUFx4f_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g560 ( .A(n_336), .Y(n_560) );
INVx6_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g491 ( .A(n_337), .Y(n_491) );
INVx1_ASAP7_75t_SL g529 ( .A(n_337), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_344), .B2(n_345), .Y(n_341) );
INVx4_ASAP7_75t_L g379 ( .A(n_343), .Y(n_379) );
BUFx3_ASAP7_75t_L g457 ( .A(n_343), .Y(n_457) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_345), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_345), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_506) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_347), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_347), .A2(n_508), .B1(n_555), .B2(n_556), .Y(n_554) );
OR2x6_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx2_ASAP7_75t_L g451 ( .A(n_351), .Y(n_451) );
INVx2_ASAP7_75t_SL g499 ( .A(n_351), .Y(n_499) );
INVx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g453 ( .A(n_354), .Y(n_453) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g395 ( .A(n_357), .Y(n_395) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
XNOR2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NAND3x1_ASAP7_75t_SL g360 ( .A(n_361), .B(n_366), .C(n_372), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g414 ( .A(n_365), .Y(n_414) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_370), .Y(n_366) );
BUFx2_ASAP7_75t_L g604 ( .A(n_369), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_381), .C(n_389), .Y(n_372) );
OAI22xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_377), .B1(n_378), .B2(n_380), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_374), .A2(n_443), .B1(n_444), .B2(n_446), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_374), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_543) );
OA211x2_ASAP7_75t_L g696 ( .A1(n_374), .A2(n_697), .B(n_698), .C(n_699), .Y(n_696) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx3_ASAP7_75t_L g497 ( .A(n_376), .Y(n_497) );
INVx3_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g508 ( .A(n_379), .Y(n_508) );
OAI21xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_385), .B(n_386), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g445 ( .A(n_383), .Y(n_445) );
BUFx4f_ASAP7_75t_L g505 ( .A(n_387), .Y(n_505) );
INVx1_ASAP7_75t_SL g582 ( .A(n_388), .Y(n_582) );
OAI22xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_391), .B1(n_392), .B2(n_393), .Y(n_389) );
INVx4_ASAP7_75t_L g624 ( .A(n_390), .Y(n_624) );
INVx1_ASAP7_75t_L g463 ( .A(n_396), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_423), .B1(n_461), .B2(n_462), .Y(n_396) );
INVx3_ASAP7_75t_SL g461 ( .A(n_397), .Y(n_461) );
XOR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_422), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_399), .B(n_409), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_400), .B(n_405), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_403), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_402), .A2(n_522), .B(n_523), .Y(n_521) );
OAI222xp33_ASAP7_75t_L g583 ( .A1(n_402), .A2(n_448), .B1(n_453), .B2(n_584), .C1(n_585), .C2(n_586), .Y(n_583) );
OAI21xp5_ASAP7_75t_SL g664 ( .A1(n_402), .A2(n_665), .B(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_417), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
INVx5_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g564 ( .A(n_416), .Y(n_564) );
INVx2_ASAP7_75t_L g693 ( .A(n_416), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_421), .Y(n_417) );
BUFx2_ASAP7_75t_L g594 ( .A(n_420), .Y(n_594) );
INVx3_ASAP7_75t_L g462 ( .A(n_423), .Y(n_462) );
BUFx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g460 ( .A(n_425), .Y(n_460) );
AND2x2_ASAP7_75t_SL g425 ( .A(n_426), .B(n_441), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_434), .Y(n_426) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
OAI221xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_436), .B1(n_437), .B2(n_439), .C(n_440), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_447), .C(n_455), .Y(n_441) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g495 ( .A(n_445), .Y(n_495) );
INVx2_ASAP7_75t_L g545 ( .A(n_445), .Y(n_545) );
OAI222xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_450), .B1(n_451), .B2(n_452), .C1(n_453), .C2(n_454), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g644 ( .A(n_466), .Y(n_644) );
AOI22xp5_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_607), .B1(n_608), .B2(n_642), .Y(n_466) );
INVx1_ASAP7_75t_L g642 ( .A(n_467), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_536), .B2(n_537), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_512), .B1(n_534), .B2(n_535), .Y(n_469) );
INVx1_ASAP7_75t_SL g534 ( .A(n_470), .Y(n_534) );
BUFx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g511 ( .A(n_473), .Y(n_511) );
AND2x2_ASAP7_75t_SL g473 ( .A(n_474), .B(n_492), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_482), .Y(n_474) );
OAI221xp5_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_477), .B1(n_478), .B2(n_480), .C(n_481), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_498), .C(n_506), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_493) );
INVx2_ASAP7_75t_L g576 ( .A(n_497), .Y(n_576) );
OA211x2_ASAP7_75t_L g634 ( .A1(n_497), .A2(n_635), .B(n_636), .C(n_637), .Y(n_634) );
OAI221xp5_ASAP7_75t_SL g498 ( .A1(n_499), .A2(n_500), .B1(n_501), .B2(n_503), .C(n_504), .Y(n_498) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g535 ( .A(n_512), .Y(n_535) );
XOR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_533), .Y(n_512) );
NAND4xp75_ASAP7_75t_SL g513 ( .A(n_514), .B(n_525), .C(n_530), .D(n_531), .Y(n_513) );
NOR2xp67_ASAP7_75t_SL g514 ( .A(n_515), .B(n_521), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .C(n_519), .Y(n_515) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
XOR2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_568), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_SL g566 ( .A(n_541), .Y(n_566) );
AND2x2_ASAP7_75t_SL g541 ( .A(n_542), .B(n_557), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .C(n_554), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_545), .A2(n_574), .B1(n_575), .B2(n_577), .C(n_578), .Y(n_573) );
OAI21xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B(n_551), .Y(n_547) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND4x1_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .C(n_561), .D(n_563), .Y(n_557) );
INVx1_ASAP7_75t_L g598 ( .A(n_564), .Y(n_598) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g606 ( .A(n_571), .Y(n_606) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_587), .Y(n_571) );
NOR2xp33_ASAP7_75t_SL g572 ( .A(n_573), .B(n_583), .Y(n_572) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_595), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_593), .Y(n_588) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_596), .B(n_600), .Y(n_595) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AO22x1_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_626), .B1(n_640), .B2(n_641), .Y(n_608) );
INVx2_ASAP7_75t_SL g640 ( .A(n_609), .Y(n_640) );
XOR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_625), .Y(n_609) );
NAND4xp75_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .C(n_620), .D(n_623), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_SL g614 ( .A(n_615), .B(n_617), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx2_ASAP7_75t_SL g641 ( .A(n_626), .Y(n_641) );
XOR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_639), .Y(n_626) );
NAND4xp75_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .C(n_634), .D(n_638), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NOR2x1_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .Y(n_646) );
OR2x2_ASAP7_75t_SL g705 ( .A(n_647), .B(n_652), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_648), .Y(n_680) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_649), .B(n_682), .Y(n_685) );
CKINVDCx16_ASAP7_75t_R g682 ( .A(n_650), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
OAI322xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_679), .A3(n_681), .B1(n_683), .B2(n_686), .C1(n_687), .C2(n_705), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND3x1_ASAP7_75t_L g662 ( .A(n_663), .B(n_672), .C(n_676), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .C(n_671), .Y(n_667) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
BUFx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
XOR2x2_ASAP7_75t_L g689 ( .A(n_686), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND4xp75_ASAP7_75t_L g690 ( .A(n_691), .B(n_696), .C(n_700), .D(n_703), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
endmodule