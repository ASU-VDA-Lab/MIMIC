module fake_jpeg_31597_n_33 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_16),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_17),
.B(n_20),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_6),
.B(n_9),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_18),
.A2(n_21),
.B(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_14),
.B(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_5),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_26),
.B1(n_14),
.B2(n_11),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_31),
.B(n_29),
.C(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);


endmodule