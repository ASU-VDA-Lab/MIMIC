module fake_jpeg_57_n_32 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_32;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_15;

INVx4_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_SL g11 ( 
.A(n_7),
.Y(n_11)
);

INVx4_ASAP7_75t_SL g12 ( 
.A(n_9),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_0),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.C(n_19),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.C(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_2),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_24),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_16),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_R g27 ( 
.A(n_26),
.B(n_13),
.Y(n_27)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_29),
.B(n_25),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_18),
.C(n_13),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_28),
.A2(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_31)
);

AOI321xp33_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C(n_30),
.Y(n_32)
);


endmodule