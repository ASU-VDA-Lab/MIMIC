module real_aes_8014_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g562 ( .A1(n_0), .A2(n_200), .B(n_563), .C(n_566), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_1), .B(n_551), .Y(n_567) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_3), .A2(n_129), .B1(n_130), .B2(n_133), .Y(n_128) );
INVx1_ASAP7_75t_L g133 ( .A(n_3), .Y(n_133) );
INVx1_ASAP7_75t_L g218 ( .A(n_4), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_5), .B(n_189), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_6), .A2(n_466), .B(n_545), .Y(n_544) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_7), .A2(n_165), .B(n_513), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_8), .A2(n_39), .B1(n_145), .B2(n_154), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_9), .B(n_165), .Y(n_229) );
AND2x6_ASAP7_75t_L g163 ( .A(n_10), .B(n_164), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_11), .A2(n_163), .B(n_469), .C(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_12), .B(n_40), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_12), .B(n_40), .Y(n_126) );
INVx1_ASAP7_75t_L g161 ( .A(n_13), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_14), .B(n_152), .Y(n_172) );
INVx1_ASAP7_75t_L g210 ( .A(n_15), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_16), .B(n_189), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_17), .B(n_166), .Y(n_234) );
AO32x2_ASAP7_75t_L g197 ( .A1(n_18), .A2(n_162), .A3(n_165), .B1(n_198), .B2(n_202), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_19), .A2(n_106), .B1(n_116), .B2(n_772), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_20), .B(n_154), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_21), .B(n_166), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_22), .A2(n_56), .B1(n_145), .B2(n_154), .Y(n_201) );
AOI22xp33_ASAP7_75t_SL g151 ( .A1(n_23), .A2(n_83), .B1(n_152), .B2(n_154), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_24), .B(n_154), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_25), .A2(n_162), .B(n_469), .C(n_471), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_26), .A2(n_448), .B1(n_753), .B2(n_754), .C1(n_763), .C2(n_767), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_27), .A2(n_162), .B(n_469), .C(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_28), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_29), .B(n_157), .Y(n_254) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_30), .A2(n_758), .B1(n_761), .B2(n_762), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_30), .Y(n_762) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_31), .A2(n_466), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_32), .B(n_157), .Y(n_195) );
INVx2_ASAP7_75t_L g147 ( .A(n_33), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_34), .A2(n_490), .B(n_499), .C(n_501), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_35), .B(n_154), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_36), .B(n_157), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_37), .A2(n_77), .B1(n_759), .B2(n_760), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_37), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_38), .B(n_174), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_41), .B(n_465), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_42), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_42), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_43), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_44), .B(n_189), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_45), .B(n_466), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_46), .A2(n_490), .B(n_499), .C(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_47), .A2(n_81), .B1(n_440), .B2(n_441), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_47), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_47), .A2(n_440), .B1(n_451), .B2(n_452), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_48), .B(n_154), .Y(n_224) );
INVx1_ASAP7_75t_L g564 ( .A(n_49), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_50), .A2(n_91), .B1(n_145), .B2(n_148), .Y(n_144) );
INVx1_ASAP7_75t_L g537 ( .A(n_51), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_52), .B(n_154), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_53), .B(n_154), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_54), .B(n_466), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_55), .B(n_216), .Y(n_228) );
AOI22xp33_ASAP7_75t_SL g238 ( .A1(n_57), .A2(n_61), .B1(n_152), .B2(n_154), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_58), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_59), .B(n_154), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_60), .B(n_154), .Y(n_253) );
INVx1_ASAP7_75t_L g164 ( .A(n_62), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_63), .B(n_466), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_64), .A2(n_100), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_64), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_64), .B(n_551), .Y(n_550) );
A2O1A1Ixp33_ASAP7_75t_L g547 ( .A1(n_65), .A2(n_213), .B(n_216), .C(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_66), .B(n_154), .Y(n_219) );
INVx1_ASAP7_75t_L g160 ( .A(n_67), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_68), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_69), .B(n_189), .Y(n_503) );
AO32x2_ASAP7_75t_L g142 ( .A1(n_70), .A2(n_143), .A3(n_156), .B1(n_162), .B2(n_165), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_71), .B(n_155), .Y(n_527) );
INVx1_ASAP7_75t_L g252 ( .A(n_72), .Y(n_252) );
INVx1_ASAP7_75t_L g187 ( .A(n_73), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g561 ( .A(n_74), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_75), .B(n_473), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_76), .A2(n_469), .B(n_486), .C(n_490), .Y(n_485) );
INVx1_ASAP7_75t_L g760 ( .A(n_77), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_78), .B(n_152), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_79), .Y(n_546) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_81), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_82), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_84), .B(n_145), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_85), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_86), .B(n_152), .Y(n_192) );
INVx2_ASAP7_75t_L g158 ( .A(n_87), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_88), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_89), .B(n_149), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_90), .B(n_152), .Y(n_225) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_92), .B(n_112), .C(n_113), .Y(n_111) );
OR2x2_ASAP7_75t_L g123 ( .A(n_92), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g455 ( .A(n_92), .B(n_125), .Y(n_455) );
INVx2_ASAP7_75t_L g752 ( .A(n_92), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_93), .A2(n_104), .B1(n_152), .B2(n_153), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_94), .B(n_466), .Y(n_497) );
INVx1_ASAP7_75t_L g502 ( .A(n_95), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_96), .B(n_444), .Y(n_443) );
INVxp67_ASAP7_75t_L g549 ( .A(n_97), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_98), .B(n_152), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_99), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g131 ( .A(n_100), .Y(n_131) );
INVx1_ASAP7_75t_L g487 ( .A(n_101), .Y(n_487) );
INVx1_ASAP7_75t_L g523 ( .A(n_102), .Y(n_523) );
AND2x2_ASAP7_75t_L g539 ( .A(n_103), .B(n_157), .Y(n_539) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx12_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g773 ( .A(n_109), .Y(n_773) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x2_ASAP7_75t_L g125 ( .A(n_112), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
OA21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_446), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g771 ( .A(n_119), .Y(n_771) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_127), .B(n_443), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_123), .Y(n_445) );
NOR2x2_ASAP7_75t_L g769 ( .A(n_124), .B(n_752), .Y(n_769) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g751 ( .A(n_125), .B(n_752), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_134), .B1(n_135), .B2(n_442), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_128), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
XOR2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_439), .Y(n_135) );
INVx2_ASAP7_75t_L g451 ( .A(n_136), .Y(n_451) );
AND3x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_359), .C(n_407), .Y(n_136) );
NOR4xp25_ASAP7_75t_L g137 ( .A(n_138), .B(n_287), .C(n_332), .D(n_346), .Y(n_137) );
OAI311xp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_203), .A3(n_230), .B1(n_240), .C1(n_255), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_167), .Y(n_139) );
OAI21xp33_ASAP7_75t_L g240 ( .A1(n_140), .A2(n_241), .B(n_243), .Y(n_240) );
AND2x2_ASAP7_75t_L g348 ( .A(n_140), .B(n_275), .Y(n_348) );
AND2x2_ASAP7_75t_L g405 ( .A(n_140), .B(n_291), .Y(n_405) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g298 ( .A(n_141), .B(n_196), .Y(n_298) );
AND2x2_ASAP7_75t_L g355 ( .A(n_141), .B(n_303), .Y(n_355) );
INVx1_ASAP7_75t_L g396 ( .A(n_141), .Y(n_396) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_142), .Y(n_264) );
AND2x2_ASAP7_75t_L g305 ( .A(n_142), .B(n_196), .Y(n_305) );
AND2x2_ASAP7_75t_L g309 ( .A(n_142), .B(n_197), .Y(n_309) );
INVx1_ASAP7_75t_L g321 ( .A(n_142), .Y(n_321) );
OAI22xp5_ASAP7_75t_SL g143 ( .A1(n_144), .A2(n_149), .B1(n_151), .B2(n_155), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx3_ASAP7_75t_L g148 ( .A(n_146), .Y(n_148) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
AND2x6_ASAP7_75t_L g469 ( .A(n_146), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g217 ( .A(n_147), .Y(n_217) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_148), .Y(n_504) );
INVx2_ASAP7_75t_L g566 ( .A(n_148), .Y(n_566) );
INVx2_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_149), .A2(n_199), .B1(n_200), .B2(n_201), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_149), .A2(n_200), .B1(n_237), .B2(n_238), .Y(n_236) );
INVx4_ASAP7_75t_L g565 ( .A(n_149), .Y(n_565) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g155 ( .A(n_150), .Y(n_155) );
INVx1_ASAP7_75t_L g174 ( .A(n_150), .Y(n_174) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
AND2x2_ASAP7_75t_L g467 ( .A(n_150), .B(n_217), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_150), .Y(n_470) );
INVx2_ASAP7_75t_L g211 ( .A(n_152), .Y(n_211) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_154), .Y(n_489) );
INVx5_ASAP7_75t_L g189 ( .A(n_155), .Y(n_189) );
INVx1_ASAP7_75t_L g476 ( .A(n_156), .Y(n_476) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_157), .A2(n_169), .B(n_179), .Y(n_168) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_157), .A2(n_184), .B(n_195), .Y(n_183) );
INVx1_ASAP7_75t_L g479 ( .A(n_157), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_157), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_157), .A2(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AND2x2_ASAP7_75t_L g166 ( .A(n_158), .B(n_159), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NAND3xp33_ASAP7_75t_L g235 ( .A(n_162), .B(n_236), .C(n_239), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_162), .A2(n_248), .B(n_251), .Y(n_247) );
BUFx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_163), .A2(n_170), .B(n_175), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_163), .A2(n_185), .B(n_190), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_163), .A2(n_209), .B(n_214), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_163), .A2(n_223), .B(n_226), .Y(n_222) );
AND2x4_ASAP7_75t_L g466 ( .A(n_163), .B(n_467), .Y(n_466) );
INVx4_ASAP7_75t_SL g491 ( .A(n_163), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g524 ( .A(n_163), .B(n_467), .Y(n_524) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_165), .A2(n_222), .B(n_229), .Y(n_221) );
INVx4_ASAP7_75t_L g239 ( .A(n_165), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_165), .A2(n_514), .B(n_515), .Y(n_513) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_165), .Y(n_543) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g202 ( .A(n_166), .Y(n_202) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_180), .Y(n_167) );
AND2x2_ASAP7_75t_L g242 ( .A(n_168), .B(n_196), .Y(n_242) );
INVx2_ASAP7_75t_L g276 ( .A(n_168), .Y(n_276) );
AND2x2_ASAP7_75t_L g291 ( .A(n_168), .B(n_197), .Y(n_291) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_168), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_168), .B(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g311 ( .A(n_168), .B(n_274), .Y(n_311) );
INVx1_ASAP7_75t_L g323 ( .A(n_168), .Y(n_323) );
INVx1_ASAP7_75t_L g364 ( .A(n_168), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_168), .B(n_264), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_173), .Y(n_170) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_178), .Y(n_175) );
O2A1O1Ixp5_ASAP7_75t_L g251 ( .A1(n_178), .A2(n_215), .B(n_252), .C(n_253), .Y(n_251) );
NOR2xp67_ASAP7_75t_L g180 ( .A(n_181), .B(n_196), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g241 ( .A(n_182), .B(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_182), .Y(n_269) );
AND2x2_ASAP7_75t_SL g322 ( .A(n_182), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g326 ( .A(n_182), .B(n_196), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_182), .B(n_321), .Y(n_384) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g274 ( .A(n_183), .Y(n_274) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_183), .Y(n_290) );
OR2x2_ASAP7_75t_L g363 ( .A(n_183), .B(n_364), .Y(n_363) );
O2A1O1Ixp5_ASAP7_75t_SL g185 ( .A1(n_186), .A2(n_187), .B(n_188), .C(n_189), .Y(n_185) );
INVx2_ASAP7_75t_L g200 ( .A(n_189), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_189), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_189), .A2(n_249), .B(n_250), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_189), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
INVx1_ASAP7_75t_L g213 ( .A(n_193), .Y(n_213) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g473 ( .A(n_194), .Y(n_473) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g270 ( .A(n_197), .Y(n_270) );
AND2x2_ASAP7_75t_L g275 ( .A(n_197), .B(n_276), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_200), .A2(n_215), .B(n_218), .C(n_219), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_200), .A2(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g207 ( .A(n_202), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_202), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_203), .B(n_258), .Y(n_421) );
INVx1_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g391 ( .A(n_204), .B(n_232), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_221), .Y(n_204) );
AND2x2_ASAP7_75t_L g267 ( .A(n_205), .B(n_258), .Y(n_267) );
INVx2_ASAP7_75t_L g279 ( .A(n_205), .Y(n_279) );
AND2x2_ASAP7_75t_L g313 ( .A(n_205), .B(n_261), .Y(n_313) );
AND2x2_ASAP7_75t_L g380 ( .A(n_205), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_206), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g260 ( .A(n_206), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g300 ( .A(n_206), .B(n_221), .Y(n_300) );
AND2x2_ASAP7_75t_L g317 ( .A(n_206), .B(n_318), .Y(n_317) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_220), .Y(n_206) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_207), .A2(n_247), .B(n_254), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .C(n_213), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_211), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_211), .A2(n_527), .B(n_528), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g486 ( .A1(n_213), .A2(n_487), .B(n_488), .C(n_489), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_215), .A2(n_472), .B(n_474), .Y(n_471) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g243 ( .A(n_221), .B(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g261 ( .A(n_221), .Y(n_261) );
AND2x2_ASAP7_75t_L g266 ( .A(n_221), .B(n_246), .Y(n_266) );
AND2x2_ASAP7_75t_L g339 ( .A(n_221), .B(n_318), .Y(n_339) );
AND2x2_ASAP7_75t_L g404 ( .A(n_221), .B(n_394), .Y(n_404) );
OAI311xp33_ASAP7_75t_L g287 ( .A1(n_230), .A2(n_288), .A3(n_292), .B1(n_294), .C1(n_314), .Y(n_287) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g299 ( .A(n_231), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g358 ( .A(n_231), .B(n_266), .Y(n_358) );
AND2x2_ASAP7_75t_L g432 ( .A(n_231), .B(n_313), .Y(n_432) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_232), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g367 ( .A(n_232), .Y(n_367) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g258 ( .A(n_233), .Y(n_258) );
NOR2x1_ASAP7_75t_L g330 ( .A(n_233), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g387 ( .A(n_233), .B(n_261), .Y(n_387) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
INVx1_ASAP7_75t_L g284 ( .A(n_234), .Y(n_284) );
AO21x1_ASAP7_75t_L g283 ( .A1(n_236), .A2(n_239), .B(n_284), .Y(n_283) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_239), .A2(n_484), .B(n_493), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_239), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_239), .B(n_506), .Y(n_505) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_239), .A2(n_522), .B(n_529), .Y(n_521) );
INVx3_ASAP7_75t_L g551 ( .A(n_239), .Y(n_551) );
AND2x2_ASAP7_75t_L g262 ( .A(n_242), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g315 ( .A(n_242), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g395 ( .A(n_242), .B(n_396), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_243), .A2(n_275), .B1(n_295), .B2(n_299), .C(n_301), .Y(n_294) );
INVx1_ASAP7_75t_L g419 ( .A(n_244), .Y(n_419) );
OR2x2_ASAP7_75t_L g385 ( .A(n_245), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g280 ( .A(n_246), .B(n_261), .Y(n_280) );
OR2x2_ASAP7_75t_L g282 ( .A(n_246), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g307 ( .A(n_246), .Y(n_307) );
INVx2_ASAP7_75t_L g318 ( .A(n_246), .Y(n_318) );
AND2x2_ASAP7_75t_L g345 ( .A(n_246), .B(n_283), .Y(n_345) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_246), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_262), .B1(n_265), .B2(n_268), .C(n_271), .Y(n_255) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g356 ( .A(n_258), .B(n_266), .Y(n_356) );
AND2x2_ASAP7_75t_L g406 ( .A(n_258), .B(n_260), .Y(n_406) );
INVx2_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g293 ( .A(n_260), .B(n_264), .Y(n_293) );
AND2x2_ASAP7_75t_L g372 ( .A(n_260), .B(n_345), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_261), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g331 ( .A(n_261), .Y(n_331) );
OAI21xp33_ASAP7_75t_L g341 ( .A1(n_262), .A2(n_342), .B(n_344), .Y(n_341) );
OR2x2_ASAP7_75t_L g285 ( .A(n_263), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g351 ( .A(n_263), .B(n_311), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_263), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g328 ( .A(n_264), .B(n_297), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_264), .B(n_411), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_265), .B(n_291), .Y(n_401) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x2_ASAP7_75t_L g324 ( .A(n_266), .B(n_279), .Y(n_324) );
INVx1_ASAP7_75t_L g340 ( .A(n_267), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_277), .B1(n_281), .B2(n_285), .Y(n_271) );
INVx2_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
INVx1_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
INVx1_ASAP7_75t_L g286 ( .A(n_275), .Y(n_286) );
AND2x2_ASAP7_75t_L g357 ( .A(n_275), .B(n_303), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_275), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
OR2x2_ASAP7_75t_L g281 ( .A(n_278), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_278), .B(n_394), .Y(n_393) );
NOR2xp67_ASAP7_75t_L g425 ( .A(n_278), .B(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g428 ( .A(n_280), .B(n_380), .Y(n_428) );
INVx1_ASAP7_75t_SL g394 ( .A(n_282), .Y(n_394) );
AND2x2_ASAP7_75t_L g334 ( .A(n_283), .B(n_318), .Y(n_334) );
INVx1_ASAP7_75t_L g381 ( .A(n_283), .Y(n_381) );
OAI222xp33_ASAP7_75t_L g422 ( .A1(n_288), .A2(n_378), .B1(n_423), .B2(n_424), .C1(n_427), .C2(n_429), .Y(n_422) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g343 ( .A(n_290), .Y(n_343) );
AND2x2_ASAP7_75t_L g354 ( .A(n_291), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_291), .B(n_396), .Y(n_423) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_293), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g398 ( .A(n_295), .Y(n_398) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g336 ( .A(n_298), .Y(n_336) );
AND2x2_ASAP7_75t_L g415 ( .A(n_298), .B(n_376), .Y(n_415) );
AND2x2_ASAP7_75t_L g438 ( .A(n_298), .B(n_322), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_300), .B(n_334), .Y(n_333) );
OAI32xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_304), .A3(n_306), .B1(n_308), .B2(n_312), .Y(n_301) );
BUFx2_ASAP7_75t_L g376 ( .A(n_303), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_304), .B(n_322), .Y(n_403) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g342 ( .A(n_305), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g410 ( .A(n_305), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g399 ( .A(n_306), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g370 ( .A(n_309), .B(n_343), .Y(n_370) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
OAI221xp5_ASAP7_75t_SL g332 ( .A1(n_311), .A2(n_333), .B1(n_335), .B2(n_337), .C(n_341), .Y(n_332) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g344 ( .A(n_313), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g350 ( .A(n_313), .B(n_334), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B1(n_319), .B2(n_324), .C(n_325), .Y(n_314) );
INVx1_ASAP7_75t_L g433 ( .A(n_315), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_316), .B(n_410), .Y(n_409) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_317), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_322), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g388 ( .A(n_322), .Y(n_388) );
BUFx3_ASAP7_75t_L g411 ( .A(n_323), .Y(n_411) );
INVx1_ASAP7_75t_SL g352 ( .A(n_324), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_324), .B(n_366), .Y(n_365) );
AOI21xp33_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_327), .B(n_329), .Y(n_325) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_326), .A2(n_427), .B1(n_431), .B2(n_433), .C(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g373 ( .A(n_331), .B(n_334), .Y(n_373) );
INVx1_ASAP7_75t_L g437 ( .A(n_331), .Y(n_437) );
INVx2_ASAP7_75t_L g426 ( .A(n_334), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_334), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g379 ( .A(n_339), .B(n_380), .Y(n_379) );
OAI221xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_349), .B1(n_351), .B2(n_352), .C(n_353), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B1(n_357), .B2(n_358), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_355), .A2(n_417), .B1(n_418), .B2(n_420), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_358), .A2(n_435), .B(n_438), .Y(n_434) );
NOR4xp25_ASAP7_75t_SL g359 ( .A(n_360), .B(n_368), .C(n_377), .D(n_397), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_365), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_371), .B1(n_374), .B2(n_375), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g413 ( .A(n_373), .Y(n_413) );
OAI221xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_382), .B1(n_385), .B2(n_388), .C(n_389), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g400 ( .A(n_380), .Y(n_400) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI21xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_392), .B(n_395), .Y(n_389) );
INVx1_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_401), .C(n_402), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_405), .B2(n_406), .Y(n_402) );
CKINVDCx14_ASAP7_75t_R g412 ( .A(n_406), .Y(n_412) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_422), .C(n_430), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .B1(n_413), .B2(n_414), .C(n_416), .Y(n_408) );
INVxp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_443), .B(n_447), .C(n_770), .Y(n_446) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI22xp5_ASAP7_75t_SL g448 ( .A1(n_449), .A2(n_453), .B1(n_456), .B2(n_749), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g763 ( .A1(n_450), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_763) );
INVx2_ASAP7_75t_L g452 ( .A(n_451), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g764 ( .A(n_454), .Y(n_764) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g765 ( .A(n_457), .Y(n_765) );
AND3x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_653), .C(n_710), .Y(n_457) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_598), .C(n_634), .Y(n_458) );
OAI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_507), .B(n_553), .C(n_585), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_480), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g556 ( .A(n_462), .B(n_557), .Y(n_556) );
INVx5_ASAP7_75t_L g584 ( .A(n_462), .Y(n_584) );
AND2x2_ASAP7_75t_L g657 ( .A(n_462), .B(n_573), .Y(n_657) );
AND2x2_ASAP7_75t_L g695 ( .A(n_462), .B(n_601), .Y(n_695) );
AND2x2_ASAP7_75t_L g715 ( .A(n_462), .B(n_558), .Y(n_715) );
OR2x6_ASAP7_75t_L g462 ( .A(n_463), .B(n_477), .Y(n_462) );
AOI21xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_468), .B(n_476), .Y(n_463) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx5_ASAP7_75t_L g500 ( .A(n_469), .Y(n_500) );
INVx2_ASAP7_75t_L g475 ( .A(n_473), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_475), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_475), .A2(n_504), .B(n_537), .C(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_480), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_495), .Y(n_480) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_481), .Y(n_596) );
AND2x2_ASAP7_75t_L g610 ( .A(n_481), .B(n_557), .Y(n_610) );
INVx1_ASAP7_75t_L g633 ( .A(n_481), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_481), .B(n_584), .Y(n_672) );
OR2x2_ASAP7_75t_L g709 ( .A(n_481), .B(n_555), .Y(n_709) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_482), .Y(n_645) );
AND2x2_ASAP7_75t_L g652 ( .A(n_482), .B(n_558), .Y(n_652) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g573 ( .A(n_483), .B(n_558), .Y(n_573) );
BUFx2_ASAP7_75t_L g601 ( .A(n_483), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_492), .Y(n_484) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_L g545 ( .A1(n_491), .A2(n_500), .B(n_546), .C(n_547), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_SL g560 ( .A1(n_491), .A2(n_500), .B(n_561), .C(n_562), .Y(n_560) );
INVx5_ASAP7_75t_L g555 ( .A(n_495), .Y(n_555) );
BUFx2_ASAP7_75t_L g577 ( .A(n_495), .Y(n_577) );
AND2x2_ASAP7_75t_L g734 ( .A(n_495), .B(n_588), .Y(n_734) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_505), .Y(n_495) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_540), .Y(n_508) );
OAI221xp5_ASAP7_75t_L g634 ( .A1(n_509), .A2(n_635), .B1(n_642), .B2(n_643), .C(n_646), .Y(n_634) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
AND2x2_ASAP7_75t_L g541 ( .A(n_510), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_510), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g569 ( .A(n_511), .B(n_520), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_511), .B(n_521), .Y(n_579) );
OR2x2_ASAP7_75t_L g590 ( .A(n_511), .B(n_542), .Y(n_590) );
AND2x2_ASAP7_75t_L g593 ( .A(n_511), .B(n_581), .Y(n_593) );
AND2x2_ASAP7_75t_L g609 ( .A(n_511), .B(n_531), .Y(n_609) );
OR2x2_ASAP7_75t_L g625 ( .A(n_511), .B(n_521), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_511), .B(n_542), .Y(n_687) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_512), .B(n_531), .Y(n_679) );
AND2x2_ASAP7_75t_L g682 ( .A(n_512), .B(n_521), .Y(n_682) );
OR2x2_ASAP7_75t_L g603 ( .A(n_519), .B(n_590), .Y(n_603) );
INVx2_ASAP7_75t_L g629 ( .A(n_519), .Y(n_629) );
OR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_531), .Y(n_519) );
AND2x2_ASAP7_75t_L g552 ( .A(n_520), .B(n_532), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_520), .B(n_542), .Y(n_608) );
OR2x2_ASAP7_75t_L g619 ( .A(n_520), .B(n_532), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_520), .B(n_581), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g711 ( .A1(n_520), .A2(n_712), .B1(n_714), .B2(n_716), .C(n_719), .Y(n_711) );
INVx5_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_521), .B(n_542), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_525), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_531), .B(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_531), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g597 ( .A(n_531), .B(n_569), .Y(n_597) );
OR2x2_ASAP7_75t_L g641 ( .A(n_531), .B(n_542), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_531), .B(n_593), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_531), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g706 ( .A(n_531), .B(n_707), .Y(n_706) );
INVx5_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_SL g570 ( .A(n_532), .B(n_541), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_SL g574 ( .A1(n_532), .A2(n_575), .B(n_578), .C(n_582), .Y(n_574) );
OR2x2_ASAP7_75t_L g612 ( .A(n_532), .B(n_608), .Y(n_612) );
OR2x2_ASAP7_75t_L g648 ( .A(n_532), .B(n_590), .Y(n_648) );
OAI311xp33_ASAP7_75t_L g654 ( .A1(n_532), .A2(n_593), .A3(n_655), .B1(n_658), .C1(n_665), .Y(n_654) );
AND2x2_ASAP7_75t_L g705 ( .A(n_532), .B(n_542), .Y(n_705) );
AND2x2_ASAP7_75t_L g713 ( .A(n_532), .B(n_568), .Y(n_713) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_532), .Y(n_731) );
AND2x2_ASAP7_75t_L g748 ( .A(n_532), .B(n_569), .Y(n_748) );
OR2x6_ASAP7_75t_L g532 ( .A(n_533), .B(n_539), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_552), .Y(n_540) );
AND2x2_ASAP7_75t_L g576 ( .A(n_541), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g732 ( .A(n_541), .Y(n_732) );
AND2x2_ASAP7_75t_L g568 ( .A(n_542), .B(n_569), .Y(n_568) );
INVx3_ASAP7_75t_L g581 ( .A(n_542), .Y(n_581) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_542), .Y(n_624) );
INVxp67_ASAP7_75t_L g663 ( .A(n_542), .Y(n_663) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B(n_550), .Y(n_542) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_551), .A2(n_559), .B(n_567), .Y(n_558) );
AND2x2_ASAP7_75t_L g741 ( .A(n_552), .B(n_589), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_568), .B1(n_570), .B2(n_571), .C(n_574), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_555), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g594 ( .A(n_555), .B(n_584), .Y(n_594) );
AND2x2_ASAP7_75t_L g602 ( .A(n_555), .B(n_557), .Y(n_602) );
OR2x2_ASAP7_75t_L g614 ( .A(n_555), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g632 ( .A(n_555), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g656 ( .A(n_555), .B(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_555), .Y(n_676) );
AND2x2_ASAP7_75t_L g728 ( .A(n_555), .B(n_652), .Y(n_728) );
OAI31xp33_ASAP7_75t_L g736 ( .A1(n_555), .A2(n_605), .A3(n_704), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_556), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g700 ( .A(n_556), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_556), .B(n_709), .Y(n_708) );
AND2x4_ASAP7_75t_L g588 ( .A(n_557), .B(n_584), .Y(n_588) );
INVx1_ASAP7_75t_L g675 ( .A(n_557), .Y(n_675) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g725 ( .A(n_558), .B(n_584), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_SL g735 ( .A(n_568), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_569), .B(n_640), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_570), .A2(n_682), .B1(n_720), .B2(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g583 ( .A(n_573), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g642 ( .A(n_573), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_573), .B(n_594), .Y(n_747) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g717 ( .A(n_576), .B(n_718), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_577), .A2(n_636), .B(n_638), .Y(n_635) );
OR2x2_ASAP7_75t_L g643 ( .A(n_577), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g664 ( .A(n_577), .B(n_652), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_577), .B(n_675), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_577), .B(n_715), .Y(n_714) );
OAI221xp5_ASAP7_75t_SL g691 ( .A1(n_578), .A2(n_692), .B1(n_697), .B2(n_700), .C(n_701), .Y(n_691) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OR2x2_ASAP7_75t_L g668 ( .A(n_579), .B(n_641), .Y(n_668) );
INVx1_ASAP7_75t_L g707 ( .A(n_579), .Y(n_707) );
INVx2_ASAP7_75t_L g683 ( .A(n_580), .Y(n_683) );
INVx1_ASAP7_75t_L g617 ( .A(n_581), .Y(n_617) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g622 ( .A(n_584), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_584), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g651 ( .A(n_584), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g739 ( .A(n_584), .B(n_709), .Y(n_739) );
AOI222xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_589), .B1(n_591), .B2(n_594), .C1(n_595), .C2(n_597), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g595 ( .A(n_588), .B(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_588), .A2(n_638), .B1(n_666), .B2(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_588), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OAI21xp33_ASAP7_75t_SL g626 ( .A1(n_597), .A2(n_627), .B(n_630), .Y(n_626) );
OAI211xp5_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_603), .B(n_604), .C(n_626), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_602), .A2(n_605), .B1(n_610), .B2(n_611), .C(n_613), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_602), .B(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g696 ( .A(n_602), .Y(n_696) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
AND2x2_ASAP7_75t_L g698 ( .A(n_607), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g615 ( .A(n_610), .Y(n_615) );
AND2x2_ASAP7_75t_L g621 ( .A(n_610), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B1(n_620), .B2(n_623), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_617), .B(n_629), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_618), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g718 ( .A(n_622), .Y(n_718) );
AND2x2_ASAP7_75t_L g737 ( .A(n_622), .B(n_652), .Y(n_737) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_629), .B(n_686), .Y(n_745) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_632), .B(n_700), .Y(n_743) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g666 ( .A(n_644), .Y(n_666) );
BUFx2_ASAP7_75t_L g690 ( .A(n_645), .Y(n_690) );
OAI21xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_649), .B(n_651), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_669), .C(n_691), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_661), .B(n_664), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_SL g669 ( .A1(n_670), .A2(n_673), .B(n_677), .C(n_680), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_670), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NOR2xp67_ASAP7_75t_SL g674 ( .A(n_675), .B(n_676), .Y(n_674) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g699 ( .A(n_679), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B(n_688), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
AND2x2_ASAP7_75t_L g704 ( .A(n_682), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B1(n_706), .B2(n_708), .Y(n_701) );
INVx2_ASAP7_75t_SL g722 ( .A(n_709), .Y(n_722) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_726), .C(n_738), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_722), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_729), .B1(n_733), .B2(n_735), .C(n_736), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g738 ( .A1(n_727), .A2(n_739), .B(n_740), .C(n_742), .Y(n_738) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_746), .B2(n_748), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g766 ( .A(n_750), .Y(n_766) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g761 ( .A(n_758), .Y(n_761) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx3_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
endmodule