module fake_jpeg_30837_n_531 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_531);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_531;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_417;
wire n_362;
wire n_142;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_58),
.Y(n_130)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_81),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_69),
.Y(n_158)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_71),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_18),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_102),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_73),
.Y(n_169)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_76),
.A2(n_41),
.B1(n_36),
.B2(n_50),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_78),
.Y(n_166)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_80),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_18),
.B(n_1),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_89),
.Y(n_173)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_96),
.Y(n_122)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_4),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_97),
.Y(n_160)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_98),
.Y(n_157)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g135 ( 
.A(n_100),
.Y(n_135)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_104),
.Y(n_123)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_35),
.B(n_4),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_31),
.C(n_36),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_28),
.Y(n_134)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_24),
.B(n_4),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_28),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_110),
.B(n_131),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_103),
.A2(n_23),
.B1(n_38),
.B2(n_42),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_112),
.A2(n_113),
.B1(n_132),
.B2(n_62),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_23),
.B1(n_38),
.B2(n_42),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_134),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_43),
.B(n_53),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_39),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_58),
.B(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_121),
.B(n_127),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_30),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_55),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_23),
.B1(n_38),
.B2(n_42),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_98),
.B(n_33),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_137),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_67),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_140),
.B(n_28),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_57),
.A2(n_44),
.B1(n_42),
.B2(n_38),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_144),
.A2(n_106),
.B1(n_102),
.B2(n_95),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_99),
.B(n_30),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_146),
.B(n_150),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_65),
.B(n_50),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_152),
.A2(n_39),
.B1(n_24),
.B2(n_27),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_76),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_93),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_80),
.C(n_56),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_175),
.B(n_216),
.C(n_125),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_115),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_185),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_43),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_211),
.Y(n_250)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_188),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_113),
.A2(n_69),
.B1(n_94),
.B2(n_100),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_189),
.A2(n_204),
.B1(n_226),
.B2(n_130),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_190),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_191),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_192),
.B(n_206),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_136),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_193),
.B(n_194),
.Y(n_253)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_196),
.B(n_202),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_135),
.A2(n_160),
.B1(n_53),
.B2(n_89),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_214),
.B1(n_222),
.B2(n_224),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx6_ASAP7_75t_SL g266 ( 
.A(n_198),
.Y(n_266)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_117),
.Y(n_199)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_227),
.B1(n_170),
.B2(n_147),
.Y(n_234)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_208),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_153),
.A2(n_77),
.B1(n_88),
.B2(n_87),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_205),
.A2(n_217),
.B1(n_45),
.B2(n_48),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_124),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_220),
.C(n_130),
.Y(n_236)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_173),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_209),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_122),
.A2(n_41),
.B(n_48),
.C(n_47),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_33),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_37),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_213),
.Y(n_267)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_126),
.Y(n_214)
);

BUFx16f_ASAP7_75t_L g215 ( 
.A(n_117),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_215),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_144),
.B(n_60),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_166),
.A2(n_86),
.B1(n_84),
.B2(n_78),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_219),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_117),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_221),
.A2(n_223),
.B1(n_147),
.B2(n_149),
.Y(n_268)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_225),
.A2(n_215),
.B1(n_199),
.B2(n_206),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_138),
.A2(n_75),
.B1(n_73),
.B2(n_83),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_228),
.B(n_232),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_201),
.B(n_27),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_203),
.A2(n_132),
.B(n_112),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_233),
.A2(n_259),
.B(n_262),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_234),
.A2(n_246),
.B1(n_261),
.B2(n_177),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_138),
.B1(n_155),
.B2(n_158),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_235),
.A2(n_209),
.B1(n_161),
.B2(n_180),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_244),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_174),
.B(n_175),
.C(n_187),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_192),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_183),
.B(n_37),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_258),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_174),
.B(n_155),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_263),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_179),
.B(n_45),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_200),
.A2(n_158),
.B1(n_141),
.B2(n_170),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_223),
.A2(n_125),
.B1(n_111),
.B2(n_164),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_174),
.B(n_161),
.Y(n_263)
);

INVx5_ASAP7_75t_SL g295 ( 
.A(n_268),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_216),
.B1(n_205),
.B2(n_227),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_269),
.A2(n_278),
.B1(n_283),
.B2(n_284),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_264),
.C(n_237),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_141),
.B1(n_149),
.B2(n_189),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_272),
.A2(n_273),
.B1(n_287),
.B2(n_296),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_186),
.B1(n_198),
.B2(n_190),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_274),
.A2(n_296),
.B1(n_238),
.B2(n_240),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_233),
.A2(n_211),
.B(n_209),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_285),
.B(n_297),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_192),
.B1(n_191),
.B2(n_195),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_250),
.B(n_210),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_281),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_253),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_248),
.Y(n_281)
);

OAI32xp33_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_257),
.A3(n_228),
.B1(n_249),
.B2(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_246),
.A2(n_213),
.B1(n_202),
.B2(n_188),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_265),
.A2(n_176),
.B(n_215),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_235),
.A2(n_181),
.B1(n_182),
.B2(n_129),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_185),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_290),
.B(n_300),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_255),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_291),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_292),
.B(n_298),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_214),
.B1(n_224),
.B2(n_145),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_230),
.A2(n_225),
.B(n_168),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_237),
.Y(n_298)
);

OAI21xp33_ASAP7_75t_SL g299 ( 
.A1(n_236),
.A2(n_148),
.B(n_221),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_299),
.A2(n_264),
.B(n_267),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_240),
.B(n_220),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_229),
.B(n_47),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_229),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_304),
.A2(n_314),
.B1(n_322),
.B2(n_326),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_306),
.B(n_318),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_276),
.B(n_264),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_SL g347 ( 
.A(n_312),
.B(n_275),
.Y(n_347)
);

INVx4_ASAP7_75t_SL g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_270),
.Y(n_333)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_288),
.Y(n_317)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_295),
.A2(n_266),
.B1(n_251),
.B2(n_252),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_319),
.Y(n_353)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_274),
.A2(n_272),
.B1(n_276),
.B2(n_281),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_277),
.Y(n_335)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_287),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_325),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_274),
.A2(n_264),
.B1(n_241),
.B2(n_267),
.Y(n_326)
);

NOR2x1_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_258),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_330),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_269),
.A2(n_266),
.B1(n_241),
.B2(n_251),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_329),
.A2(n_298),
.B1(n_291),
.B2(n_292),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_271),
.A2(n_238),
.B1(n_245),
.B2(n_254),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_275),
.A2(n_238),
.B(n_231),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_271),
.Y(n_340)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_326),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_321),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_334),
.B(n_343),
.Y(n_372)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_335),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_271),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_344),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_271),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_355),
.C(n_313),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_345),
.B(n_350),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_327),
.A2(n_303),
.B1(n_310),
.B2(n_332),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_342),
.A2(n_352),
.B1(n_360),
.B2(n_315),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_305),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_278),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_331),
.Y(n_345)
);

A2O1A1Ixp33_ASAP7_75t_SL g375 ( 
.A1(n_347),
.A2(n_312),
.B(n_315),
.C(n_308),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_280),
.Y(n_348)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_348),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_283),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_279),
.Y(n_355)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_303),
.A2(n_282),
.A3(n_290),
.B1(n_293),
.B2(n_284),
.Y(n_357)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_357),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_325),
.A2(n_295),
.B1(n_294),
.B2(n_297),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_302),
.B(n_313),
.Y(n_361)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_361),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_323),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_302),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_370),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_322),
.C(n_306),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_366),
.B(n_376),
.C(n_377),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_367),
.A2(n_373),
.B1(n_379),
.B2(n_381),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_357),
.Y(n_371)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_350),
.A2(n_330),
.B1(n_304),
.B2(n_320),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_390),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_333),
.B(n_339),
.C(n_336),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_285),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_378),
.B(n_252),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_350),
.A2(n_325),
.B1(n_295),
.B2(n_294),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_380),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_342),
.A2(n_305),
.B1(n_317),
.B2(n_309),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_356),
.B(n_309),
.C(n_307),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_383),
.C(n_389),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_301),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_384),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_340),
.A2(n_297),
.B(n_328),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_386),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_351),
.A2(n_328),
.B(n_289),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_354),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_54),
.Y(n_420)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_289),
.Y(n_389)
);

OA21x2_ASAP7_75t_L g390 ( 
.A1(n_341),
.A2(n_252),
.B(n_231),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_360),
.A2(n_242),
.B1(n_239),
.B2(n_254),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_393),
.B1(n_346),
.B2(n_358),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_359),
.A2(n_242),
.B1(n_239),
.B2(n_245),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_365),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_394),
.B(n_421),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_349),
.Y(n_397)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_397),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_391),
.A2(n_345),
.B(n_353),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_399),
.B(n_422),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_349),
.Y(n_400)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_400),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_364),
.Y(n_402)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_351),
.B1(n_353),
.B2(n_337),
.Y(n_403)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_368),
.A2(n_341),
.B1(n_345),
.B2(n_337),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_409),
.A2(n_416),
.B1(n_392),
.B2(n_379),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_390),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_410),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_346),
.Y(n_411)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_411),
.Y(n_436)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_389),
.A2(n_242),
.B1(n_254),
.B2(n_239),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_376),
.B(n_256),
.C(n_247),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_418),
.C(n_370),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_374),
.B(n_256),
.C(n_247),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_245),
.Y(n_419)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_419),
.Y(n_443)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_363),
.B(n_382),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_383),
.B(n_5),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_374),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_433),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_366),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_430),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_396),
.B(n_404),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_434),
.A2(n_442),
.B1(n_444),
.B2(n_403),
.Y(n_454)
);

XNOR2x1_ASAP7_75t_L g435 ( 
.A(n_407),
.B(n_375),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_SL g456 ( 
.A(n_435),
.B(n_399),
.C(n_401),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_404),
.B(n_377),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_445),
.C(n_418),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_405),
.A2(n_373),
.B1(n_375),
.B2(n_151),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_405),
.A2(n_375),
.B1(n_151),
.B2(n_142),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_142),
.Y(n_445)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_431),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_446),
.B(n_449),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_402),
.Y(n_447)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_447),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_428),
.A2(n_415),
.B1(n_412),
.B2(n_395),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_424),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_453),
.Y(n_479)
);

XNOR2x1_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_456),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_428),
.A2(n_410),
.B1(n_412),
.B2(n_411),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_452),
.A2(n_442),
.B1(n_434),
.B2(n_443),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_429),
.A2(n_395),
.B1(n_400),
.B2(n_419),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_454),
.A2(n_437),
.B1(n_441),
.B2(n_445),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_438),
.B(n_417),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_458),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_416),
.C(n_398),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_457),
.B(n_460),
.C(n_462),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_408),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_398),
.C(n_413),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_440),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_461),
.B(n_425),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_397),
.C(n_409),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g470 ( 
.A(n_463),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_429),
.A2(n_401),
.B1(n_408),
.B2(n_44),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_464),
.Y(n_466)
);

MAJx2_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_435),
.C(n_401),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_476),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_452),
.A2(n_436),
.B(n_423),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_467),
.A2(n_29),
.B(n_10),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_469),
.A2(n_454),
.B1(n_462),
.B2(n_463),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_472),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_450),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_451),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_475),
.A2(n_448),
.B1(n_6),
.B2(n_7),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_426),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_427),
.C(n_44),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_477),
.B(n_480),
.C(n_54),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_44),
.C(n_54),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_482),
.B(n_489),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_481),
.B(n_460),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_486),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_490),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_471),
.A2(n_448),
.B(n_6),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_496),
.B(n_494),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_467),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_491),
.B(n_492),
.Y(n_505)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_478),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_29),
.C(n_6),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_493),
.B(n_495),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_470),
.A2(n_29),
.B1(n_6),
.B2(n_9),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_494),
.A2(n_466),
.B1(n_475),
.B2(n_11),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_468),
.B(n_5),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_496),
.A2(n_466),
.B1(n_465),
.B2(n_11),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_497),
.B(n_508),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_490),
.A2(n_474),
.B(n_479),
.Y(n_498)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_498),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_499),
.B(n_504),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_502),
.A2(n_503),
.B1(n_488),
.B2(n_483),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g503 ( 
.A1(n_482),
.A2(n_474),
.B1(n_480),
.B2(n_476),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_487),
.A2(n_477),
.B1(n_10),
.B2(n_11),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_9),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_484),
.Y(n_509)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_509),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_501),
.Y(n_510)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_510),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_511),
.B(n_515),
.C(n_513),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_506),
.B(n_483),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_514),
.A2(n_507),
.B(n_497),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_489),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_518),
.B(n_519),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_503),
.C(n_508),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_11),
.C(n_12),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_520),
.A2(n_516),
.B(n_513),
.Y(n_522)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_522),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_523),
.A2(n_517),
.B(n_14),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_525),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_527),
.B(n_524),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_526),
.C(n_13),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_529),
.B(n_13),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_16),
.B(n_361),
.Y(n_531)
);


endmodule