module fake_jpeg_12811_n_181 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_4),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_36),
.B(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_9),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_50),
.Y(n_54)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_19),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_1),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_1),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_42),
.B1(n_49),
.B2(n_41),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_61),
.B1(n_65),
.B2(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_33),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_52),
.C(n_21),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_68),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_46),
.B1(n_35),
.B2(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_16),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_16),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_31),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_21),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx24_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_30),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_97),
.Y(n_121)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_100),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_52),
.C(n_22),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_102),
.C(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_13),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_52),
.B1(n_23),
.B2(n_22),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_99),
.B1(n_96),
.B2(n_66),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_22),
.B1(n_2),
.B2(n_11),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_3),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_2),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_66),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_57),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_115),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_87),
.A2(n_66),
.B1(n_63),
.B2(n_62),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_12),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_101),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_94),
.B(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_138),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_128),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_89),
.B1(n_84),
.B2(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_131),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_104),
.A2(n_106),
.B1(n_111),
.B2(n_116),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_92),
.B1(n_93),
.B2(n_99),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_94),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_137),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_145),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_110),
.C(n_112),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_147),
.B(n_150),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_103),
.C(n_108),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_130),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_113),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_155),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_127),
.B(n_123),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_154),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_135),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_157),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_126),
.B(n_127),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_123),
.B1(n_142),
.B2(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_144),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_158),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_141),
.C(n_137),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_159),
.C(n_163),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_157),
.A2(n_128),
.B1(n_118),
.B2(n_79),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_160),
.B(n_153),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_168),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_169),
.A2(n_171),
.B1(n_164),
.B2(n_67),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_166),
.A2(n_155),
.B1(n_79),
.B2(n_86),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_173),
.C(n_174),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_161),
.C(n_63),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_109),
.C(n_73),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_177),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_174),
.B(n_176),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_67),
.B(n_69),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_73),
.Y(n_181)
);


endmodule