module fake_jpeg_14950_n_359 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_359);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_18),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_49),
.Y(n_69)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_59),
.Y(n_85)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_31),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

OR2x4_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_23),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_35),
.Y(n_97)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_93),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_65),
.Y(n_117)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

BUFx16f_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_111),
.Y(n_120)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_101),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_53),
.B1(n_79),
.B2(n_83),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_112),
.B1(n_74),
.B2(n_32),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_53),
.B1(n_22),
.B2(n_25),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_97),
.B1(n_35),
.B2(n_84),
.Y(n_130)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_59),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_34),
.B1(n_36),
.B2(n_25),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_39),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_44),
.B1(n_34),
.B2(n_22),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_117),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_54),
.C(n_72),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_42),
.C(n_50),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_78),
.B1(n_70),
.B2(n_38),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_131),
.B1(n_135),
.B2(n_137),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_128),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_132),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_61),
.B1(n_44),
.B2(n_40),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_92),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_37),
.B(n_57),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_129),
.B(n_131),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_61),
.B1(n_40),
.B2(n_51),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_38),
.B1(n_43),
.B2(n_51),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_65),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_57),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_51),
.B1(n_50),
.B2(n_43),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_142),
.A2(n_86),
.B1(n_96),
.B2(n_91),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_100),
.B1(n_109),
.B2(n_90),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_157),
.B1(n_160),
.B2(n_142),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_96),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_158),
.C(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_91),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_155),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_150),
.A2(n_165),
.B(n_143),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_126),
.B1(n_141),
.B2(n_125),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_23),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_132),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_129),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_135),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_28),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_128),
.B1(n_123),
.B2(n_115),
.Y(n_160)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_27),
.B(n_29),
.Y(n_165)
);

CKINVDCx12_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_168),
.A2(n_122),
.B1(n_113),
.B2(n_99),
.Y(n_190)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_105),
.B1(n_103),
.B2(n_101),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_188),
.B1(n_133),
.B2(n_105),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_182),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_144),
.Y(n_179)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_114),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_28),
.C(n_23),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_164),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_114),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_186),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_147),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_160),
.B(n_121),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_126),
.B1(n_125),
.B2(n_136),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_28),
.CI(n_30),
.CON(n_189),
.SN(n_189)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_189),
.B(n_30),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_159),
.B1(n_163),
.B2(n_168),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_197),
.B(n_165),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_161),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_122),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_28),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_150),
.A2(n_143),
.B(n_86),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_146),
.B1(n_145),
.B2(n_151),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_199),
.A2(n_213),
.B1(n_223),
.B2(n_189),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_201),
.B1(n_214),
.B2(n_173),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_158),
.A3(n_151),
.B1(n_152),
.B2(n_157),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_204),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_197),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_28),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_216),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_0),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_210),
.B(n_222),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_170),
.B(n_2),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_174),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_212),
.B(n_215),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_181),
.A2(n_133),
.B1(n_161),
.B2(n_98),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_174),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_42),
.C(n_50),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_175),
.B1(n_182),
.B2(n_193),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_29),
.C(n_33),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_216),
.Y(n_247)
);

INVx13_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_221),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_10),
.B(n_16),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_176),
.A2(n_29),
.B1(n_33),
.B2(n_3),
.Y(n_223)
);

CKINVDCx12_ASAP7_75t_R g224 ( 
.A(n_172),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_188),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_247),
.C(n_179),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_215),
.Y(n_230)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_185),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_237),
.B1(n_244),
.B2(n_209),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_203),
.B(n_177),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_233),
.B(n_193),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_234),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_236),
.Y(n_261)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_238),
.A2(n_242),
.B1(n_245),
.B2(n_218),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_243),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g240 ( 
.A1(n_200),
.A2(n_210),
.B(n_213),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_199),
.B1(n_208),
.B2(n_221),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_195),
.B1(n_171),
.B2(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_190),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_187),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_249),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_245),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_209),
.B1(n_208),
.B2(n_205),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_254),
.A2(n_33),
.B1(n_3),
.B2(n_1),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_206),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_258),
.C(n_263),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_223),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_267),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_187),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_227),
.A2(n_179),
.B1(n_10),
.B2(n_11),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_264),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_268),
.C(n_270),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_240),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_30),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_30),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_33),
.C(n_30),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_263),
.C(n_266),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_243),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_248),
.Y(n_284)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_252),
.B(n_225),
.CI(n_230),
.CON(n_277),
.SN(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_283),
.C(n_286),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_234),
.C(n_228),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_284),
.B(n_292),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_232),
.B1(n_244),
.B2(n_241),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_285),
.A2(n_288),
.B1(n_289),
.B2(n_291),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_250),
.C(n_248),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_249),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_287),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_259),
.A2(n_244),
.B1(n_8),
.B2(n_10),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_261),
.B1(n_255),
.B2(n_253),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_258),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_256),
.A2(n_7),
.B(n_14),
.Y(n_292)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_254),
.B(n_270),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_295),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_271),
.Y(n_296)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_7),
.B(n_4),
.C(n_5),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_298),
.A2(n_12),
.B(n_290),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_275),
.A2(n_1),
.B(n_4),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_301),
.A2(n_302),
.B(n_300),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_33),
.Y(n_303)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

OA21x2_ASAP7_75t_SL g304 ( 
.A1(n_283),
.A2(n_4),
.B(n_5),
.Y(n_304)
);

OAI21x1_ASAP7_75t_SL g319 ( 
.A1(n_304),
.A2(n_293),
.B(n_288),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_281),
.B(n_6),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_309),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_278),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_308),
.A2(n_291),
.B1(n_277),
.B2(n_12),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_277),
.B(n_12),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_274),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_312),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_282),
.C(n_274),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_311),
.B(n_322),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_280),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_280),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_316),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_319),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_300),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_299),
.Y(n_325)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_325),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_297),
.B1(n_294),
.B2(n_299),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_297),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_328),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_301),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_316),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_298),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_335),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_337),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_308),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_310),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_342),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_294),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_L g343 ( 
.A(n_333),
.B(n_311),
.C(n_314),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_326),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_339),
.A2(n_324),
.B(n_329),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_346),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_324),
.C(n_329),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_347),
.B(n_348),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_334),
.C(n_343),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_350),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_345),
.B(n_349),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_352),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_351),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_344),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_357),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_326),
.Y(n_359)
);


endmodule