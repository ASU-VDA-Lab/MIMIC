module real_jpeg_2848_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_1),
.A2(n_40),
.B1(n_48),
.B2(n_49),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_1),
.A2(n_40),
.B1(n_65),
.B2(n_66),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_57),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_2),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_3),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_96),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_96),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_96),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_164),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_5),
.B(n_47),
.C(n_49),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_5),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_5),
.B(n_46),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_5),
.B(n_62),
.C(n_65),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_199),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_5),
.B(n_86),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_5),
.B(n_67),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_199),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_54),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_10),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_70),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_13),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_135),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_135),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_135),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_14),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_14),
.A2(n_28),
.B1(n_48),
.B2(n_49),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_28),
.B1(n_65),
.B2(n_66),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_15),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_163),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_15),
.A2(n_48),
.B1(n_49),
.B2(n_163),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_163),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_110),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_108),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_20),
.B(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_78),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_72),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_41),
.B2(n_71),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_22),
.A2(n_23),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_23),
.B(n_42),
.C(n_59),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_31),
.B2(n_39),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_24),
.A2(n_31),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_25),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_26),
.A2(n_29),
.B(n_199),
.C(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_26),
.B(n_199),
.Y(n_200)
);

AOI32xp33_ASAP7_75t_L g211 ( 
.A1(n_26),
.A2(n_33),
.A3(n_35),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_29),
.A2(n_31),
.B1(n_39),
.B2(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_29),
.A2(n_133),
.B(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_30),
.A2(n_134),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_38),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_31),
.B(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_31),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_31),
.A2(n_93),
.B(n_285),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_33),
.B1(n_47),
.B2(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_32),
.B(n_189),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g213 ( 
.A(n_32),
.B(n_36),
.Y(n_213)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_53),
.B1(n_55),
.B2(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_44),
.A2(n_55),
.B1(n_56),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_44),
.A2(n_55),
.B1(n_74),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_44),
.A2(n_55),
.B1(n_172),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_44),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_44),
.A2(n_203),
.B(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_45),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_46),
.B(n_160),
.Y(n_265)
);

AO22x1_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_46)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_49),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_49),
.B(n_238),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_55),
.A2(n_131),
.B(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_55),
.A2(n_159),
.B(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_59),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_67),
.B(n_68),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_60),
.A2(n_67),
.B1(n_91),
.B2(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_60),
.A2(n_67),
.B1(n_129),
.B2(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_60),
.A2(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_60),
.B(n_185),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_69),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_76),
.B1(n_77),
.B2(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_64),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_64),
.A2(n_206),
.B(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_64),
.A2(n_76),
.B1(n_182),
.B2(n_232),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_65),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_67),
.B(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_76),
.A2(n_184),
.B(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B(n_92),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_79),
.A2(n_80),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_89),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_82),
.B1(n_92),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_81),
.A2(n_82),
.B1(n_89),
.B2(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_86),
.B(n_87),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_83),
.A2(n_86),
.B1(n_126),
.B2(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_83),
.A2(n_199),
.B(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_84),
.A2(n_85),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_84),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_84),
.A2(n_85),
.B1(n_179),
.B2(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_84),
.A2(n_224),
.B(n_225),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_84),
.A2(n_85),
.B1(n_224),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_85),
.A2(n_178),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_85),
.B(n_193),
.Y(n_226)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_86),
.A2(n_192),
.B(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_89),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_138),
.B(n_313),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_112),
.B(n_114),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_121),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_130),
.C(n_132),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_123),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_124),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_132),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_137),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_165),
.B(n_312),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_144),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_141),
.B(n_144),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_150),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_145),
.B(n_148),
.Y(n_310)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_150),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_157),
.C(n_161),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_151),
.A2(n_152),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_153),
.B(n_155),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_154),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_156),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_161),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_162),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_307),
.B(n_311),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_276),
.B(n_304),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_218),
.B(n_275),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_194),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_169),
.B(n_194),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.C(n_186),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_170),
.B(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_174),
.C(n_177),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_180),
.B(n_186),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_208),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_195),
.B(n_209),
.C(n_217),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_207),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_196),
.B(n_202),
.C(n_204),
.Y(n_289)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_200),
.Y(n_212)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_217),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_210),
.B(n_215),
.Y(n_280)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_270),
.B(n_274),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_259),
.B(n_269),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_241),
.B(n_258),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_235),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_235),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_227),
.B1(n_233),
.B2(n_234),
.Y(n_222)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_227),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_230),
.C(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_252),
.B(n_257),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_247),
.B(n_251),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_250),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_255),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_261),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_267),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_266),
.C(n_267),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_291),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_290),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_290),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_279),
.B(n_288),
.C(n_289),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_282),
.C(n_286),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_286),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_303),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_303),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_297),
.C(n_299),
.Y(n_308)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_300),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_309),
.Y(n_311)
);


endmodule