module real_jpeg_23548_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_249;
wire n_288;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx8_ASAP7_75t_SL g68 ( 
.A(n_3),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_4),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_4),
.B(n_75),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_4),
.B(n_31),
.C(n_50),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_161),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_4),
.B(n_122),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_4),
.A2(n_91),
.B1(n_229),
.B2(n_232),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_5),
.A2(n_46),
.B1(n_69),
.B2(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_46),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_6),
.A2(n_35),
.B1(n_69),
.B2(n_70),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_6),
.A2(n_35),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_7),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_7),
.A2(n_69),
.B1(n_70),
.B2(n_116),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_116),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_116),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_8),
.A2(n_60),
.B1(n_69),
.B2(n_70),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_60),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_60),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_9),
.A2(n_32),
.B1(n_61),
.B2(n_63),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_9),
.A2(n_32),
.B1(n_69),
.B2(n_70),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_9),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_55),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_10),
.A2(n_55),
.B1(n_69),
.B2(n_70),
.Y(n_123)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_11),
.B(n_68),
.C(n_69),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_13),
.A2(n_62),
.B1(n_137),
.B2(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_13),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_13),
.A2(n_69),
.B1(n_70),
.B2(n_165),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_165),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_165),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_15),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_148),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_146),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_117),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_19),
.B(n_117),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_88),
.C(n_99),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_20),
.A2(n_21),
.B1(n_88),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_56),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_22),
.B(n_76),
.C(n_87),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_25),
.A2(n_91),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_27),
.A2(n_33),
.B(n_179),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_29),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_29),
.A2(n_91),
.B(n_104),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_37),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_31),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_30),
.B(n_235),
.Y(n_234)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_34),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_36),
.A2(n_103),
.B1(n_105),
.B2(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_36),
.A2(n_105),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_38),
.Y(n_233)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_42),
.A2(n_52),
.B(n_109),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_44),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_43),
.A2(n_80),
.B(n_244),
.C(n_246),
.Y(n_243)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_44),
.B(n_204),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_L g246 ( 
.A(n_44),
.B(n_69),
.C(n_79),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_47),
.B(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_47),
.A2(n_96),
.B(n_126),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_47),
.A2(n_53),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_47),
.A2(n_53),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_48),
.A2(n_52),
.B1(n_208),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_48),
.A2(n_125),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_52),
.B(n_161),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_53),
.B(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_54),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_76),
.B1(n_77),
.B2(n_87),
.Y(n_56)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_64),
.B(n_73),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_59),
.A2(n_65),
.B1(n_75),
.B2(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_63),
.B1(n_67),
.B2(n_68),
.Y(n_72)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_64),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_64),
.A2(n_66),
.B1(n_164),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_65),
.A2(n_75),
.B1(n_160),
.B2(n_163),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_67),
.A2(n_70),
.B(n_162),
.C(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_70),
.B1(n_79),
.B2(n_80),
.Y(n_84)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g245 ( 
.A(n_70),
.B(n_161),
.CON(n_245),
.SN(n_245)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_74),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_75),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_82),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_78),
.A2(n_173),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_83),
.A2(n_122),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_83),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_83),
.A2(n_122),
.B1(n_194),
.B2(n_245),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_88),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_98),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_89),
.A2(n_90),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_93),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_91),
.A2(n_106),
.B1(n_222),
.B2(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_92),
.B(n_161),
.Y(n_235)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_99),
.B(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_111),
.C(n_114),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_100),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_108),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_108),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_111),
.B(n_114),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_112),
.B(n_122),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_115),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_117)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_128),
.B1(n_141),
.B2(n_142),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_124),
.B(n_127),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_124),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_140),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_161),
.Y(n_162)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_143),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_286),
.B(n_291),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_196),
.B(n_277),
.C(n_285),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_183),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_151),
.B(n_183),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_166),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_153),
.B(n_154),
.C(n_166),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.C(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_185),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_175),
.B2(n_182),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_169),
.B(n_171),
.C(n_182),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B(n_174),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_177),
.B1(n_180),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_184),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_186),
.B(n_188),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.C(n_192),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_192),
.B(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_276),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_271),
.B(n_275),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_256),
.B(n_270),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_239),
.B(n_255),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_218),
.B(n_238),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_205),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_213),
.C(n_216),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_217),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_225),
.B(n_237),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_224),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_230),
.B(n_236),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_228),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_254),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_254),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_249),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_250),
.C(n_251),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_247),
.B2(n_248),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_258),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_266),
.C(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_282),
.C(n_284),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);


endmodule