module real_aes_7414_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g229 ( .A1(n_0), .A2(n_230), .B(n_231), .C(n_235), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_1), .B(n_171), .Y(n_236) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_2), .B(n_105), .C(n_106), .Y(n_104) );
INVx1_ASAP7_75t_L g454 ( .A(n_2), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_3), .B(n_143), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_4), .A2(n_129), .B(n_134), .C(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_5), .A2(n_124), .B(n_536), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_6), .A2(n_124), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_7), .B(n_171), .Y(n_542) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_8), .A2(n_159), .B(n_175), .Y(n_174) );
AND2x6_ASAP7_75t_L g129 ( .A(n_9), .B(n_130), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_10), .A2(n_129), .B(n_134), .C(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g480 ( .A(n_11), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_12), .B(n_40), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_12), .B(n_40), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_13), .B(n_234), .Y(n_500) );
INVx1_ASAP7_75t_L g153 ( .A(n_14), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_15), .B(n_143), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_16), .A2(n_144), .B(n_488), .C(n_490), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_17), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_18), .B(n_171), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_19), .B(n_208), .Y(n_579) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_20), .A2(n_134), .B(n_185), .C(n_204), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_21), .A2(n_183), .B(n_233), .C(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_22), .B(n_234), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_23), .B(n_234), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g527 ( .A(n_24), .Y(n_527) );
INVx1_ASAP7_75t_L g519 ( .A(n_25), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_26), .A2(n_134), .B(n_178), .C(n_185), .Y(n_177) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_27), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_28), .Y(n_496) );
INVx1_ASAP7_75t_L g576 ( .A(n_29), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_30), .A2(n_124), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g127 ( .A(n_31), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_32), .A2(n_132), .B(n_147), .C(n_193), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_33), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_34), .A2(n_233), .B(n_539), .C(n_541), .Y(n_538) );
INVxp67_ASAP7_75t_L g577 ( .A(n_35), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_36), .B(n_180), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_37), .A2(n_134), .B(n_185), .C(n_518), .Y(n_517) );
CKINVDCx14_ASAP7_75t_R g537 ( .A(n_38), .Y(n_537) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_39), .A2(n_98), .B1(n_462), .B2(n_739), .C1(n_740), .C2(n_743), .Y(n_461) );
INVx1_ASAP7_75t_L g739 ( .A(n_39), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_41), .A2(n_235), .B(n_478), .C(n_479), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_42), .B(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_43), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_44), .A2(n_116), .B1(n_117), .B2(n_447), .Y(n_115) );
INVx1_ASAP7_75t_L g447 ( .A(n_44), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_45), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_46), .B(n_124), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_47), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_48), .Y(n_573) );
A2O1A1Ixp33_ASAP7_75t_L g131 ( .A1(n_49), .A2(n_132), .B(n_137), .C(n_147), .Y(n_131) );
INVx1_ASAP7_75t_L g232 ( .A(n_50), .Y(n_232) );
INVx1_ASAP7_75t_L g138 ( .A(n_51), .Y(n_138) );
INVx1_ASAP7_75t_L g508 ( .A(n_52), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_53), .B(n_124), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_54), .Y(n_211) );
CKINVDCx14_ASAP7_75t_R g476 ( .A(n_55), .Y(n_476) );
INVx1_ASAP7_75t_L g130 ( .A(n_56), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_57), .B(n_124), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_58), .B(n_171), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_59), .A2(n_165), .B(n_167), .C(n_169), .Y(n_164) );
INVx1_ASAP7_75t_L g152 ( .A(n_60), .Y(n_152) );
INVx1_ASAP7_75t_SL g540 ( .A(n_61), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_62), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_63), .B(n_143), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_64), .B(n_171), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_65), .B(n_144), .Y(n_246) );
INVx1_ASAP7_75t_L g530 ( .A(n_66), .Y(n_530) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_67), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_68), .B(n_140), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_69), .A2(n_134), .B(n_147), .C(n_217), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g163 ( .A(n_70), .Y(n_163) );
INVx1_ASAP7_75t_L g108 ( .A(n_71), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_72), .A2(n_124), .B(n_475), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_73), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_74), .A2(n_124), .B(n_485), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_75), .A2(n_202), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g486 ( .A(n_76), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_77), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_78), .B(n_139), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_79), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_80), .A2(n_124), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g489 ( .A(n_81), .Y(n_489) );
INVx2_ASAP7_75t_L g150 ( .A(n_82), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_83), .A2(n_100), .B1(n_109), .B2(n_747), .Y(n_99) );
INVx1_ASAP7_75t_L g499 ( .A(n_84), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_85), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_86), .B(n_234), .Y(n_247) );
INVx2_ASAP7_75t_L g105 ( .A(n_87), .Y(n_105) );
OR2x2_ASAP7_75t_L g451 ( .A(n_87), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g738 ( .A(n_87), .B(n_453), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_88), .A2(n_134), .B(n_147), .C(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_89), .B(n_124), .Y(n_191) );
INVx1_ASAP7_75t_L g194 ( .A(n_90), .Y(n_194) );
INVxp67_ASAP7_75t_L g168 ( .A(n_91), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_92), .B(n_159), .Y(n_481) );
INVx2_ASAP7_75t_L g511 ( .A(n_93), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_94), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g218 ( .A(n_95), .Y(n_218) );
INVx1_ASAP7_75t_L g242 ( .A(n_96), .Y(n_242) );
AND2x2_ASAP7_75t_L g154 ( .A(n_97), .B(n_149), .Y(n_154) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_SL g747 ( .A(n_102), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_104), .Y(n_102) );
OR2x2_ASAP7_75t_L g467 ( .A(n_105), .B(n_453), .Y(n_467) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_105), .B(n_452), .Y(n_742) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OA21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_114), .B(n_460), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g746 ( .A(n_113), .Y(n_746) );
OAI21xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_448), .B(n_456), .Y(n_114) );
AOI22x1_ASAP7_75t_SL g744 ( .A1(n_116), .A2(n_464), .B1(n_735), .B2(n_745), .Y(n_744) );
INVx4_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_117), .A2(n_464), .B1(n_468), .B2(n_735), .Y(n_463) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OR5x1_ASAP7_75t_L g118 ( .A(n_119), .B(n_320), .C(n_398), .D(n_422), .E(n_439), .Y(n_118) );
OAI211xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_186), .B(n_237), .C(n_297), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_155), .Y(n_120) );
AND2x2_ASAP7_75t_L g251 ( .A(n_121), .B(n_157), .Y(n_251) );
INVx5_ASAP7_75t_SL g279 ( .A(n_121), .Y(n_279) );
AND2x2_ASAP7_75t_L g315 ( .A(n_121), .B(n_300), .Y(n_315) );
OR2x2_ASAP7_75t_L g354 ( .A(n_121), .B(n_156), .Y(n_354) );
OR2x2_ASAP7_75t_L g385 ( .A(n_121), .B(n_276), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_121), .B(n_289), .Y(n_421) );
AND2x2_ASAP7_75t_L g433 ( .A(n_121), .B(n_276), .Y(n_433) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_154), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_131), .B(n_149), .Y(n_122) );
BUFx2_ASAP7_75t_L g202 ( .A(n_124), .Y(n_202) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_125), .B(n_129), .Y(n_243) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
INVx1_ASAP7_75t_L g169 ( .A(n_126), .Y(n_169) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g135 ( .A(n_127), .Y(n_135) );
INVx1_ASAP7_75t_L g184 ( .A(n_127), .Y(n_184) );
INVx1_ASAP7_75t_L g136 ( .A(n_128), .Y(n_136) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_128), .Y(n_141) );
INVx3_ASAP7_75t_L g144 ( .A(n_128), .Y(n_144) );
INVx1_ASAP7_75t_L g180 ( .A(n_128), .Y(n_180) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_128), .Y(n_234) );
INVx4_ASAP7_75t_SL g148 ( .A(n_129), .Y(n_148) );
BUFx3_ASAP7_75t_L g185 ( .A(n_129), .Y(n_185) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_133), .A2(n_148), .B(n_163), .C(n_164), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_SL g227 ( .A1(n_133), .A2(n_148), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_133), .A2(n_148), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g485 ( .A1(n_133), .A2(n_148), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_133), .A2(n_148), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_133), .A2(n_148), .B(n_537), .C(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_SL g572 ( .A1(n_133), .A2(n_148), .B(n_573), .C(n_574), .Y(n_572) );
INVx5_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx3_ASAP7_75t_L g146 ( .A(n_135), .Y(n_146) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_135), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_142), .C(n_145), .Y(n_137) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_139), .A2(n_145), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp5_ASAP7_75t_L g498 ( .A1(n_139), .A2(n_499), .B(n_500), .C(n_501), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_139), .A2(n_501), .B(n_530), .C(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g166 ( .A(n_141), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_143), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g230 ( .A(n_143), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_143), .A2(n_207), .B(n_519), .C(n_520), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_143), .A2(n_166), .B1(n_576), .B2(n_577), .Y(n_575) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_144), .B(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g235 ( .A(n_146), .Y(n_235) );
INVx1_ASAP7_75t_L g490 ( .A(n_146), .Y(n_490) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_149), .A2(n_191), .B(n_192), .Y(n_190) );
INVx2_ASAP7_75t_L g209 ( .A(n_149), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_149), .A2(n_474), .B(n_481), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_149), .A2(n_243), .B(n_516), .C(n_517), .Y(n_515) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_L g160 ( .A(n_150), .B(n_151), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
AND2x2_ASAP7_75t_L g432 ( .A(n_155), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
OR2x2_ASAP7_75t_L g295 ( .A(n_156), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_173), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_157), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_157), .Y(n_288) );
INVx3_ASAP7_75t_L g303 ( .A(n_157), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_157), .B(n_173), .Y(n_327) );
OR2x2_ASAP7_75t_L g336 ( .A(n_157), .B(n_279), .Y(n_336) );
AND2x2_ASAP7_75t_L g340 ( .A(n_157), .B(n_300), .Y(n_340) );
AND2x2_ASAP7_75t_L g346 ( .A(n_157), .B(n_347), .Y(n_346) );
INVxp67_ASAP7_75t_L g383 ( .A(n_157), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_157), .B(n_240), .Y(n_397) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_161), .B(n_170), .Y(n_157) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_158), .A2(n_484), .B(n_491), .Y(n_483) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_158), .A2(n_506), .B(n_512), .Y(n_505) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_158), .A2(n_535), .B(n_542), .Y(n_534) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g172 ( .A(n_159), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_159), .A2(n_176), .B(n_177), .Y(n_175) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g250 ( .A(n_160), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_165), .A2(n_218), .B(n_219), .C(n_220), .Y(n_217) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_166), .B(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_166), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g207 ( .A(n_169), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_169), .B(n_575), .Y(n_574) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_171), .A2(n_226), .B(n_236), .Y(n_225) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_172), .B(n_197), .Y(n_196) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_172), .A2(n_215), .B(n_223), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_172), .B(n_224), .Y(n_223) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_172), .A2(n_241), .B(n_248), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_172), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_172), .B(n_522), .Y(n_521) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_172), .A2(n_526), .B(n_532), .Y(n_525) );
OR2x2_ASAP7_75t_L g289 ( .A(n_173), .B(n_240), .Y(n_289) );
AND2x2_ASAP7_75t_L g300 ( .A(n_173), .B(n_276), .Y(n_300) );
AND2x2_ASAP7_75t_L g312 ( .A(n_173), .B(n_303), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_173), .B(n_240), .Y(n_335) );
INVx1_ASAP7_75t_SL g347 ( .A(n_173), .Y(n_347) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g239 ( .A(n_174), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_174), .B(n_279), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_181), .B(n_182), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_182), .A2(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_198), .Y(n_187) );
AND2x2_ASAP7_75t_L g260 ( .A(n_188), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_188), .B(n_213), .Y(n_264) );
AND2x2_ASAP7_75t_L g267 ( .A(n_188), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_188), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g292 ( .A(n_188), .B(n_283), .Y(n_292) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_188), .Y(n_311) );
AND2x2_ASAP7_75t_L g332 ( .A(n_188), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g342 ( .A(n_188), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g388 ( .A(n_188), .B(n_271), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_188), .B(n_294), .Y(n_415) );
INVx5_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g285 ( .A(n_189), .Y(n_285) );
AND2x2_ASAP7_75t_L g351 ( .A(n_189), .B(n_283), .Y(n_351) );
AND2x2_ASAP7_75t_L g435 ( .A(n_189), .B(n_303), .Y(n_435) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_196), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_198), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_198), .Y(n_424) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_213), .Y(n_198) );
AND2x2_ASAP7_75t_L g254 ( .A(n_199), .B(n_255), .Y(n_254) );
AND2x4_ASAP7_75t_L g263 ( .A(n_199), .B(n_261), .Y(n_263) );
INVx5_ASAP7_75t_L g271 ( .A(n_199), .Y(n_271) );
AND2x2_ASAP7_75t_L g294 ( .A(n_199), .B(n_225), .Y(n_294) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_199), .Y(n_331) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_210), .Y(n_199) );
AOI21xp5_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_203), .B(n_208), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_209), .B(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_212), .A2(n_495), .B(n_502), .Y(n_494) );
INVx1_ASAP7_75t_L g372 ( .A(n_213), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_213), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g405 ( .A(n_213), .B(n_271), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_213), .A2(n_328), .B(n_435), .C(n_436), .Y(n_434) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_225), .Y(n_213) );
BUFx2_ASAP7_75t_L g255 ( .A(n_214), .Y(n_255) );
INVx2_ASAP7_75t_L g259 ( .A(n_214), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_222), .Y(n_215) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx3_ASAP7_75t_L g541 ( .A(n_221), .Y(n_541) );
INVx2_ASAP7_75t_L g261 ( .A(n_225), .Y(n_261) );
AND2x2_ASAP7_75t_L g268 ( .A(n_225), .B(n_259), .Y(n_268) );
AND2x2_ASAP7_75t_L g359 ( .A(n_225), .B(n_271), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_233), .B(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g478 ( .A(n_234), .Y(n_478) );
INVx2_ASAP7_75t_L g501 ( .A(n_235), .Y(n_501) );
AOI211x1_ASAP7_75t_SL g237 ( .A1(n_238), .A2(n_252), .B(n_265), .C(n_290), .Y(n_237) );
INVx1_ASAP7_75t_L g356 ( .A(n_238), .Y(n_356) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_251), .Y(n_238) );
INVx5_ASAP7_75t_SL g276 ( .A(n_240), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_240), .B(n_346), .Y(n_345) );
AOI311xp33_ASAP7_75t_L g364 ( .A1(n_240), .A2(n_365), .A3(n_367), .B(n_368), .C(n_374), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_240), .A2(n_312), .B(n_400), .C(n_403), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_244), .Y(n_241) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_243), .A2(n_496), .B(n_497), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_243), .A2(n_527), .B(n_528), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g569 ( .A(n_250), .Y(n_569) );
INVxp67_ASAP7_75t_L g319 ( .A(n_251), .Y(n_319) );
NAND4xp25_ASAP7_75t_SL g252 ( .A(n_253), .B(n_256), .C(n_262), .D(n_264), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_253), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g310 ( .A(n_254), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_257), .B(n_263), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_257), .B(n_270), .Y(n_390) );
BUFx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_258), .B(n_271), .Y(n_408) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g283 ( .A(n_259), .Y(n_283) );
INVxp67_ASAP7_75t_L g318 ( .A(n_260), .Y(n_318) );
AND2x4_ASAP7_75t_L g270 ( .A(n_261), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g344 ( .A(n_261), .B(n_283), .Y(n_344) );
INVx1_ASAP7_75t_L g371 ( .A(n_261), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_261), .B(n_358), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_262), .B(n_332), .Y(n_352) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_263), .B(n_285), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_263), .B(n_332), .Y(n_431) );
INVx1_ASAP7_75t_L g442 ( .A(n_264), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_269), .B(n_272), .C(n_280), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g284 ( .A(n_268), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g322 ( .A(n_268), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g304 ( .A(n_269), .Y(n_304) );
AND2x2_ASAP7_75t_L g281 ( .A(n_270), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_270), .B(n_332), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_270), .B(n_351), .Y(n_375) );
OR2x2_ASAP7_75t_L g291 ( .A(n_271), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g323 ( .A(n_271), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_271), .B(n_283), .Y(n_338) );
AND2x2_ASAP7_75t_L g395 ( .A(n_271), .B(n_351), .Y(n_395) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_271), .Y(n_402) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_273), .A2(n_285), .B1(n_407), .B2(n_409), .C(n_412), .Y(n_406) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g296 ( .A(n_276), .B(n_279), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_276), .B(n_346), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_276), .B(n_303), .Y(n_411) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g396 ( .A(n_278), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g410 ( .A(n_278), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_279), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g307 ( .A(n_279), .B(n_300), .Y(n_307) );
AND2x2_ASAP7_75t_L g377 ( .A(n_279), .B(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_279), .B(n_326), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_279), .B(n_427), .Y(n_426) );
OAI21xp5_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_284), .B(n_286), .Y(n_280) );
INVx2_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g333 ( .A(n_283), .Y(n_333) );
OR2x2_ASAP7_75t_L g337 ( .A(n_285), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g440 ( .A(n_285), .B(n_408), .Y(n_440) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AOI21xp33_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_293), .B(n_295), .Y(n_290) );
INVx1_ASAP7_75t_L g444 ( .A(n_291), .Y(n_444) );
INVx2_ASAP7_75t_SL g358 ( .A(n_292), .Y(n_358) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g439 ( .A1(n_295), .A2(n_376), .B(n_440), .C(n_441), .Y(n_439) );
OAI322xp33_ASAP7_75t_SL g308 ( .A1(n_296), .A2(n_309), .A3(n_312), .B1(n_313), .B2(n_314), .C1(n_316), .C2(n_319), .Y(n_308) );
INVx2_ASAP7_75t_L g328 ( .A(n_296), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B1(n_305), .B2(n_307), .C(n_308), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI22xp33_ASAP7_75t_SL g374 ( .A1(n_299), .A2(n_375), .B1(n_376), .B2(n_379), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_300), .B(n_303), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_300), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g373 ( .A(n_302), .B(n_335), .Y(n_373) );
INVx1_ASAP7_75t_L g363 ( .A(n_303), .Y(n_363) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_307), .A2(n_417), .B(n_419), .Y(n_416) );
AOI21xp33_ASAP7_75t_L g341 ( .A1(n_309), .A2(n_342), .B(n_345), .Y(n_341) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2xp67_ASAP7_75t_SL g370 ( .A(n_311), .B(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_311), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g427 ( .A(n_312), .Y(n_427) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND4xp25_ASAP7_75t_L g320 ( .A(n_321), .B(n_348), .C(n_364), .D(n_380), .Y(n_320) );
AOI211xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B(n_329), .C(n_341), .Y(n_321) );
INVx1_ASAP7_75t_L g413 ( .A(n_322), .Y(n_413) );
AND2x2_ASAP7_75t_L g361 ( .A(n_323), .B(n_344), .Y(n_361) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_328), .B(n_363), .Y(n_362) );
OAI22xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_334), .B1(n_337), .B2(n_339), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_331), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g379 ( .A(n_332), .Y(n_379) );
O2A1O1Ixp33_ASAP7_75t_L g393 ( .A1(n_332), .A2(n_371), .B(n_394), .C(n_396), .Y(n_393) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g378 ( .A(n_335), .Y(n_378) );
INVx1_ASAP7_75t_L g438 ( .A(n_336), .Y(n_438) );
NAND2xp33_ASAP7_75t_SL g428 ( .A(n_337), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g367 ( .A(n_346), .Y(n_367) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B(n_353), .C(n_355), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_360), .B2(n_362), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_358), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_363), .B(n_384), .Y(n_446) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI21xp33_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_372), .B(n_373), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_386), .B1(n_389), .B2(n_391), .C(n_393), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_396), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_412) );
NAND3xp33_ASAP7_75t_SL g398 ( .A(n_399), .B(n_406), .C(n_416), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B(n_425), .C(n_434), .Y(n_422) );
INVx1_ASAP7_75t_L g443 ( .A(n_423), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B1(n_430), .B2(n_432), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B1(n_444), .B2(n_445), .Y(n_441) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g459 ( .A(n_451), .Y(n_459) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_456), .B(n_461), .C(n_746), .Y(n_460) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g745 ( .A(n_468), .Y(n_745) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_665), .Y(n_468) );
NAND5xp2_ASAP7_75t_L g469 ( .A(n_470), .B(n_580), .C(n_612), .D(n_629), .E(n_652), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_513), .B1(n_543), .B2(n_547), .C(n_551), .Y(n_470) );
INVx1_ASAP7_75t_L g692 ( .A(n_471), .Y(n_692) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_492), .Y(n_471) );
AND3x2_ASAP7_75t_L g667 ( .A(n_472), .B(n_494), .C(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_482), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_473), .B(n_549), .Y(n_548) );
BUFx3_ASAP7_75t_L g558 ( .A(n_473), .Y(n_558) );
AND2x2_ASAP7_75t_L g562 ( .A(n_473), .B(n_504), .Y(n_562) );
INVx2_ASAP7_75t_L g589 ( .A(n_473), .Y(n_589) );
OR2x2_ASAP7_75t_L g600 ( .A(n_473), .B(n_505), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_473), .B(n_493), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_473), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g679 ( .A(n_473), .B(n_505), .Y(n_679) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_482), .Y(n_561) );
AND2x2_ASAP7_75t_L g620 ( .A(n_482), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_482), .B(n_493), .Y(n_639) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g550 ( .A(n_483), .B(n_493), .Y(n_550) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_483), .Y(n_557) );
AND2x2_ASAP7_75t_L g606 ( .A(n_483), .B(n_505), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_483), .B(n_492), .C(n_589), .Y(n_631) );
AND2x2_ASAP7_75t_L g696 ( .A(n_483), .B(n_494), .Y(n_696) );
AND2x2_ASAP7_75t_L g730 ( .A(n_483), .B(n_493), .Y(n_730) );
INVxp67_ASAP7_75t_L g559 ( .A(n_492), .Y(n_559) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_504), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_493), .B(n_589), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_493), .B(n_620), .Y(n_628) );
AND2x2_ASAP7_75t_L g678 ( .A(n_493), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g706 ( .A(n_493), .Y(n_706) );
INVx4_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g613 ( .A(n_494), .B(n_606), .Y(n_613) );
BUFx3_ASAP7_75t_L g645 ( .A(n_494), .Y(n_645) );
INVx2_ASAP7_75t_L g621 ( .A(n_504), .Y(n_621) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_505), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_513), .A2(n_681), .B1(n_683), .B2(n_684), .Y(n_680) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .Y(n_513) );
AND2x2_ASAP7_75t_L g543 ( .A(n_514), .B(n_544), .Y(n_543) );
INVx3_ASAP7_75t_SL g554 ( .A(n_514), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_514), .B(n_584), .Y(n_616) );
OR2x2_ASAP7_75t_L g635 ( .A(n_514), .B(n_524), .Y(n_635) );
AND2x2_ASAP7_75t_L g640 ( .A(n_514), .B(n_592), .Y(n_640) );
AND2x2_ASAP7_75t_L g643 ( .A(n_514), .B(n_585), .Y(n_643) );
AND2x2_ASAP7_75t_L g655 ( .A(n_514), .B(n_534), .Y(n_655) );
AND2x2_ASAP7_75t_L g671 ( .A(n_514), .B(n_525), .Y(n_671) );
AND2x4_ASAP7_75t_L g674 ( .A(n_514), .B(n_545), .Y(n_674) );
OR2x2_ASAP7_75t_L g691 ( .A(n_514), .B(n_627), .Y(n_691) );
OR2x2_ASAP7_75t_L g722 ( .A(n_514), .B(n_567), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_514), .B(n_650), .Y(n_724) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_521), .Y(n_514) );
AND2x2_ASAP7_75t_L g598 ( .A(n_523), .B(n_565), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_523), .B(n_585), .Y(n_717) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_534), .Y(n_523) );
AND2x2_ASAP7_75t_L g553 ( .A(n_524), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g584 ( .A(n_524), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g592 ( .A(n_524), .B(n_567), .Y(n_592) );
AND2x2_ASAP7_75t_L g610 ( .A(n_524), .B(n_545), .Y(n_610) );
OR2x2_ASAP7_75t_L g627 ( .A(n_524), .B(n_585), .Y(n_627) );
INVx2_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
BUFx2_ASAP7_75t_L g546 ( .A(n_525), .Y(n_546) );
AND2x2_ASAP7_75t_L g650 ( .A(n_525), .B(n_534), .Y(n_650) );
INVx2_ASAP7_75t_L g545 ( .A(n_534), .Y(n_545) );
INVx1_ASAP7_75t_L g662 ( .A(n_534), .Y(n_662) );
AND2x2_ASAP7_75t_L g712 ( .A(n_534), .B(n_554), .Y(n_712) );
AND2x2_ASAP7_75t_L g564 ( .A(n_544), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g596 ( .A(n_544), .B(n_554), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_544), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
AND2x2_ASAP7_75t_L g583 ( .A(n_545), .B(n_554), .Y(n_583) );
OR2x2_ASAP7_75t_L g699 ( .A(n_546), .B(n_673), .Y(n_699) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_549), .B(n_679), .Y(n_685) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
OAI32xp33_ASAP7_75t_L g641 ( .A1(n_550), .A2(n_642), .A3(n_644), .B1(n_646), .B2(n_647), .Y(n_641) );
OR2x2_ASAP7_75t_L g658 ( .A(n_550), .B(n_600), .Y(n_658) );
OAI21xp33_ASAP7_75t_SL g683 ( .A1(n_550), .A2(n_560), .B(n_588), .Y(n_683) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_555), .B1(n_560), .B2(n_563), .Y(n_551) );
INVxp33_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_553), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_554), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g609 ( .A(n_554), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g709 ( .A(n_554), .B(n_650), .Y(n_709) );
OR2x2_ASAP7_75t_L g733 ( .A(n_554), .B(n_627), .Y(n_733) );
AOI21xp33_ASAP7_75t_L g716 ( .A1(n_555), .A2(n_615), .B(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g593 ( .A(n_557), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_557), .B(n_562), .Y(n_611) );
AND2x2_ASAP7_75t_L g633 ( .A(n_558), .B(n_606), .Y(n_633) );
INVx1_ASAP7_75t_L g646 ( .A(n_558), .Y(n_646) );
OR2x2_ASAP7_75t_L g651 ( .A(n_558), .B(n_585), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_561), .B(n_600), .Y(n_599) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_562), .A2(n_582), .B1(n_587), .B2(n_591), .Y(n_581) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_565), .A2(n_624), .B1(n_631), .B2(n_632), .Y(n_630) );
AND2x2_ASAP7_75t_L g708 ( .A(n_565), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_567), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g727 ( .A(n_567), .B(n_610), .Y(n_727) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B(n_578), .Y(n_567) );
INVx1_ASAP7_75t_L g586 ( .A(n_568), .Y(n_586) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OA21x2_ASAP7_75t_L g585 ( .A1(n_571), .A2(n_579), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_593), .B1(n_594), .B2(n_599), .C(n_601), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_583), .B(n_585), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_583), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g602 ( .A(n_584), .Y(n_602) );
O2A1O1Ixp33_ASAP7_75t_L g689 ( .A1(n_584), .A2(n_690), .B(n_691), .C(n_692), .Y(n_689) );
AND2x2_ASAP7_75t_L g694 ( .A(n_584), .B(n_674), .Y(n_694) );
O2A1O1Ixp33_ASAP7_75t_SL g732 ( .A1(n_584), .A2(n_673), .B(n_733), .C(n_734), .Y(n_732) );
BUFx3_ASAP7_75t_L g624 ( .A(n_585), .Y(n_624) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_588), .B(n_645), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g707 ( .A1(n_588), .A2(n_708), .B(n_710), .C(n_716), .Y(n_707) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVxp67_ASAP7_75t_L g668 ( .A(n_590), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_592), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
AOI211xp5_ASAP7_75t_L g612 ( .A1(n_596), .A2(n_613), .B(n_614), .C(n_622), .Y(n_612) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g697 ( .A(n_600), .Y(n_697) );
OR2x2_ASAP7_75t_L g714 ( .A(n_600), .B(n_644), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B1(n_608), .B2(n_611), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g614 ( .A1(n_603), .A2(n_615), .B1(n_616), .B2(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_607), .Y(n_604) );
OR2x2_ASAP7_75t_L g701 ( .A(n_605), .B(n_645), .Y(n_701) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g656 ( .A(n_606), .B(n_646), .Y(n_656) );
INVx1_ASAP7_75t_L g664 ( .A(n_607), .Y(n_664) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_610), .B(n_624), .Y(n_672) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_620), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g729 ( .A(n_621), .Y(n_729) );
AOI21xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .B(n_628), .Y(n_622) );
INVx1_ASAP7_75t_L g659 ( .A(n_623), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_624), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_624), .B(n_655), .Y(n_654) );
NAND2x1p5_ASAP7_75t_L g675 ( .A(n_624), .B(n_650), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_624), .B(n_671), .Y(n_682) );
OAI211xp5_ASAP7_75t_L g686 ( .A1(n_624), .A2(n_634), .B(n_674), .C(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
AOI221xp5_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_634), .B1(n_636), .B2(n_640), .C(n_641), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_638), .B(n_646), .Y(n_720) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g731 ( .A1(n_640), .A2(n_655), .B(n_657), .C(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_643), .B(n_650), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_644), .B(n_697), .Y(n_734) );
CKINVDCx16_ASAP7_75t_R g644 ( .A(n_645), .Y(n_644) );
INVxp33_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
AOI21xp33_ASAP7_75t_SL g660 ( .A1(n_649), .A2(n_661), .B(n_663), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_649), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_650), .B(n_704), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B1(n_657), .B2(n_659), .C(n_660), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_656), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g690 ( .A(n_662), .Y(n_690) );
NAND5xp2_ASAP7_75t_L g665 ( .A(n_666), .B(n_693), .C(n_707), .D(n_718), .E(n_731), .Y(n_665) );
AOI211xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B(n_676), .C(n_689), .Y(n_666) );
INVx2_ASAP7_75t_SL g713 ( .A(n_667), .Y(n_713) );
NAND4xp25_ASAP7_75t_SL g669 ( .A(n_670), .B(n_672), .C(n_673), .D(n_675), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI211xp5_ASAP7_75t_SL g676 ( .A1(n_675), .A2(n_677), .B(n_680), .C(n_686), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_678), .A2(n_719), .B1(n_721), .B2(n_723), .C(n_725), .Y(n_718) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI221xp5_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_695), .B1(n_698), .B2(n_700), .C(n_702), .Y(n_693) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_701), .A2(n_724), .B1(n_726), .B2(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_710) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
endmodule