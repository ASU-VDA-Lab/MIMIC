module fake_jpeg_4514_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_42),
.Y(n_72)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx12_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_52),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_23),
.B1(n_43),
.B2(n_36),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_32),
.B1(n_25),
.B2(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_16),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_61),
.C(n_19),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_23),
.B1(n_33),
.B2(n_21),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_50),
.A2(n_63),
.B1(n_64),
.B2(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_21),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_21),
.Y(n_54)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_33),
.B1(n_16),
.B2(n_22),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_32),
.B1(n_22),
.B2(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_36),
.A2(n_32),
.B1(n_22),
.B2(n_29),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_17),
.B1(n_20),
.B2(n_25),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_76),
.B1(n_83),
.B2(n_85),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_24),
.B1(n_28),
.B2(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_19),
.C(n_28),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_93),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_24),
.B1(n_28),
.B2(n_18),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_89),
.B1(n_92),
.B2(n_95),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_55),
.B1(n_58),
.B2(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_69),
.B1(n_59),
.B2(n_67),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_17),
.B1(n_19),
.B2(n_11),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_31),
.B1(n_19),
.B2(n_27),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_56),
.C(n_60),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_88),
.C(n_94),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_49),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_109),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_76),
.B(n_72),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_53),
.B1(n_68),
.B2(n_72),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_110),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_114),
.B1(n_116),
.B2(n_77),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_117),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_48),
.B1(n_62),
.B2(n_31),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_48),
.B1(n_62),
.B2(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_81),
.B(n_78),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_120),
.Y(n_146)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_57),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_98),
.B1(n_87),
.B2(n_115),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_138),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_81),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_143),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_80),
.B1(n_89),
.B2(n_79),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_132),
.A2(n_137),
.B1(n_147),
.B2(n_74),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_45),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_117),
.C(n_103),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_92),
.B(n_79),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_122),
.B(n_101),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_79),
.B1(n_87),
.B2(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_77),
.B1(n_82),
.B2(n_87),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_99),
.A2(n_87),
.B1(n_88),
.B2(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_108),
.A2(n_95),
.B(n_94),
.C(n_74),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_114),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_108),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_160),
.C(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_154),
.B(n_156),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_155),
.A2(n_180),
.B(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_157),
.B(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_99),
.B1(n_108),
.B2(n_104),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_169),
.A2(n_74),
.B1(n_139),
.B2(n_124),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_129),
.A2(n_108),
.B(n_109),
.C(n_100),
.D(n_107),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_134),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_179),
.B(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_177),
.B1(n_148),
.B2(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_202),
.C(n_180),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_190),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_204),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_141),
.B1(n_144),
.B2(n_143),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_185),
.A2(n_199),
.B1(n_201),
.B2(n_154),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_131),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_192),
.Y(n_233)
);

NOR2x1_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_173),
.Y(n_189)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_167),
.C(n_121),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_135),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_197),
.B(n_198),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_128),
.B(n_152),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_128),
.B(n_126),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_151),
.B1(n_132),
.B2(n_147),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_151),
.B1(n_125),
.B2(n_126),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_136),
.C(n_130),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_130),
.B(n_105),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_57),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_164),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_166),
.B1(n_139),
.B2(n_66),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_179),
.C(n_157),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_169),
.C(n_170),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_188),
.C(n_198),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_218),
.C(n_197),
.Y(n_240)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_162),
.C(n_161),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_224),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_205),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_174),
.Y(n_222)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_150),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_223),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_172),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_184),
.B(n_185),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_199),
.Y(n_242)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_230),
.B1(n_231),
.B2(n_57),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_232),
.B1(n_191),
.B2(n_201),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_167),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_229),
.B(n_27),
.Y(n_250)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_238),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_248),
.C(n_249),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_243),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_186),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_186),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_27),
.C(n_65),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_27),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_250),
.B(n_254),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_27),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_66),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_46),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_46),
.C(n_1),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_220),
.B1(n_229),
.B2(n_209),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_256),
.A2(n_260),
.B1(n_266),
.B2(n_3),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_246),
.B(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_240),
.A2(n_212),
.B1(n_213),
.B2(n_218),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_227),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_251),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_221),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_267),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_232),
.B1(n_46),
.B2(n_2),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_15),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_272),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_0),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_15),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_14),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_248),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_275),
.B(n_283),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_284),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_235),
.B(n_249),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_278),
.A2(n_280),
.B(n_282),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_235),
.B(n_1),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_0),
.C(n_1),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_14),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_2),
.C(n_3),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_2),
.B(n_3),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_285),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_290),
.B(n_13),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_285),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_13),
.B(n_12),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_273),
.B1(n_267),
.B2(n_264),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_292),
.B(n_294),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_265),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_303),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_261),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_280),
.C(n_290),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_302),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_264),
.B1(n_259),
.B2(n_261),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_282),
.B(n_259),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_284),
.C(n_11),
.Y(n_313)
);

INVx11_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_8),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_281),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_306),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_300),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_298),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_314),
.A2(n_295),
.B1(n_292),
.B2(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_315),
.B(n_318),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_312),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_317),
.A2(n_320),
.B(n_313),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_305),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_311),
.A2(n_299),
.B(n_9),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_8),
.Y(n_321)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_321),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_10),
.C(n_309),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_323),
.A2(n_327),
.B(n_326),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_311),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_324),
.A2(n_328),
.B(n_317),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_330),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_325),
.C(n_316),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_314),
.Y(n_333)
);


endmodule