module fake_jpeg_29398_n_347 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_347);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_347;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_0),
.B(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_19),
.B(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_8),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_31),
.B1(n_16),
.B2(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_64),
.B1(n_26),
.B2(n_25),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_54),
.B(n_56),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_55),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_49),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_31),
.B1(n_16),
.B2(n_24),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_67),
.B(n_74),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_29),
.B1(n_23),
.B2(n_21),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_78),
.B1(n_80),
.B2(n_25),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_21),
.B1(n_29),
.B2(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_72),
.B1(n_18),
.B2(n_24),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_37),
.A2(n_29),
.B1(n_23),
.B2(n_21),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_30),
.B1(n_34),
.B2(n_21),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_29),
.B1(n_23),
.B2(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_32),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_27),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_85),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_36),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_52),
.B1(n_50),
.B2(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_87),
.A2(n_120),
.B1(n_75),
.B2(n_79),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_88),
.A2(n_97),
.B1(n_32),
.B2(n_27),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_90),
.B(n_95),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_96),
.Y(n_137)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_61),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_25),
.B1(n_20),
.B2(n_26),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_26),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_98),
.Y(n_140)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_81),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_100),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_65),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_121),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_59),
.A2(n_19),
.B1(n_16),
.B2(n_33),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_54),
.A2(n_28),
.B1(n_17),
.B2(n_26),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_70),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_65),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_25),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_118),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_56),
.Y(n_118)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_20),
.B1(n_28),
.B2(n_17),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_67),
.B(n_9),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_27),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_125),
.B1(n_77),
.B2(n_71),
.Y(n_131)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_149),
.B1(n_97),
.B2(n_95),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_131),
.A2(n_123),
.B(n_110),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_77),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_136),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_86),
.A2(n_75),
.B1(n_79),
.B2(n_71),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_144),
.B1(n_147),
.B2(n_155),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_76),
.B1(n_60),
.B2(n_27),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_100),
.A2(n_60),
.B1(n_27),
.B2(n_32),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_87),
.B1(n_105),
.B2(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_158),
.A2(n_165),
.B1(n_174),
.B2(n_182),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_101),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_160),
.B(n_162),
.Y(n_206)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_121),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_145),
.B(n_89),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_166),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_93),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_164),
.B(n_175),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_98),
.B1(n_103),
.B2(n_117),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_89),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_186),
.Y(n_193)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_98),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_170),
.C(n_172),
.Y(n_221)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_96),
.C(n_113),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_137),
.B(n_96),
.CI(n_120),
.CON(n_171),
.SN(n_171)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_177),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_96),
.C(n_93),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_120),
.B1(n_115),
.B2(n_109),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_156),
.B(n_106),
.Y(n_175)
);

OR2x2_ASAP7_75t_SL g176 ( 
.A(n_128),
.B(n_136),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_181),
.B(n_135),
.Y(n_214)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

BUFx4f_ASAP7_75t_SL g178 ( 
.A(n_142),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_183),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_120),
.C(n_114),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_187),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_126),
.A2(n_122),
.B1(n_92),
.B2(n_99),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_112),
.C(n_11),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_125),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_55),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_32),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_144),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_143),
.A2(n_32),
.B(n_2),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_139),
.B(n_127),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_189),
.A2(n_182),
.B1(n_190),
.B2(n_180),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_0),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_149),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_129),
.A2(n_55),
.B1(n_9),
.B2(n_11),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_148),
.B1(n_146),
.B2(n_127),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_194),
.A2(n_198),
.B1(n_200),
.B2(n_204),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_187),
.B1(n_173),
.B2(n_158),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_199),
.A2(n_2),
.B(n_3),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_165),
.B1(n_171),
.B2(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_201),
.B(n_5),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_215),
.B1(n_6),
.B2(n_12),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_139),
.B1(n_142),
.B2(n_151),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_151),
.B1(n_135),
.B2(n_130),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_5),
.B1(n_200),
.B2(n_199),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_132),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_216),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_176),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_224),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_189),
.B(n_167),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_172),
.A2(n_152),
.B1(n_132),
.B2(n_133),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_0),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_0),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_4),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_219),
.Y(n_240)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_220),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_55),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_222),
.A2(n_167),
.B(n_178),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_191),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_225),
.B(n_237),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_206),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_226),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_236),
.B(n_201),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_6),
.C(n_13),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_218),
.Y(n_266)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_196),
.A2(n_6),
.B1(n_12),
.B2(n_14),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_241),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_214),
.Y(n_259)
);

AO22x1_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_239),
.B(n_247),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_203),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_14),
.C(n_4),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_221),
.C(n_194),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_246),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_210),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_244),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_5),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_197),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_193),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_193),
.B(n_212),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_224),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_207),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_252),
.B(n_254),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_255),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_223),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_238),
.Y(n_255)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_266),
.Y(n_286)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_269),
.Y(n_288)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_216),
.C(n_223),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_209),
.C(n_215),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_230),
.C(n_242),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_208),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_225),
.Y(n_289)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_243),
.B1(n_250),
.B2(n_196),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_281),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_234),
.B1(n_239),
.B2(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_248),
.B1(n_236),
.B2(n_227),
.Y(n_280)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_263),
.A2(n_248),
.B1(n_245),
.B2(n_235),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_286),
.Y(n_294)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_285),
.Y(n_299)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_256),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_272),
.Y(n_300)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_290),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_265),
.A2(n_246),
.B1(n_231),
.B2(n_222),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_291),
.A2(n_293),
.B1(n_270),
.B2(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_292),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_264),
.A2(n_251),
.B1(n_229),
.B2(n_231),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_300),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_274),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_307),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_268),
.C(n_273),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_308),
.C(n_277),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_263),
.B1(n_253),
.B2(n_262),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_305),
.A2(n_293),
.B1(n_291),
.B2(n_284),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_259),
.B1(n_262),
.B2(n_274),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_229),
.C(n_266),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_276),
.Y(n_309)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_309),
.Y(n_328)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_312),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_288),
.C(n_289),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_314),
.Y(n_323)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_319),
.C(n_320),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_252),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_294),
.B(n_258),
.C(n_292),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_290),
.C(n_285),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_304),
.A2(n_275),
.B1(n_267),
.B2(n_230),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_306),
.C(n_300),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_325),
.B(n_311),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_295),
.Y(n_327)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_327),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_310),
.A2(n_295),
.B(n_307),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_320),
.B(n_267),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_328),
.B(n_326),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_331),
.A2(n_333),
.B(n_334),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_336),
.Y(n_338)
);

OAI21x1_ASAP7_75t_SL g333 ( 
.A1(n_329),
.A2(n_302),
.B(n_303),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_322),
.A2(n_316),
.B(n_298),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_322),
.A2(n_192),
.B(n_220),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_337),
.A2(n_325),
.B(n_324),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_341),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_330),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_247),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_339),
.C(n_228),
.Y(n_344)
);

AOI322xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_192),
.A3(n_228),
.B1(n_205),
.B2(n_342),
.C1(n_233),
.C2(n_232),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_205),
.Y(n_346)
);

NAND2xp33_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_237),
.Y(n_347)
);


endmodule