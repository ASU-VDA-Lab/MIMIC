module fake_jpeg_8597_n_113 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_0),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_67),
.B(n_68),
.C(n_57),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_65),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_0),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_16),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_48),
.B1(n_45),
.B2(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_75),
.B1(n_80),
.B2(n_38),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_58),
.B1(n_52),
.B2(n_50),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_76),
.B1(n_81),
.B2(n_85),
.Y(n_88)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_49),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_77),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_86),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_89),
.Y(n_98)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_20),
.C(n_23),
.Y(n_92)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_25),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_99),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_100),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_96),
.B(n_98),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_88),
.C(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_92),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_95),
.C(n_97),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_91),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_107),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_31),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_94),
.B(n_34),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g113 ( 
.A(n_112),
.Y(n_113)
);


endmodule