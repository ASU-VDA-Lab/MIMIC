module fake_jpeg_8888_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_294;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_33),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_53),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_24),
.B1(n_30),
.B2(n_18),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_21),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_22),
.B1(n_17),
.B2(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_61),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_41),
.B1(n_37),
.B2(n_42),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_41),
.B1(n_42),
.B2(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_66),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_81),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_42),
.B(n_8),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_31),
.B(n_2),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_94),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_91),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_84),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_41),
.B1(n_28),
.B2(n_32),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_77),
.A2(n_86),
.B1(n_96),
.B2(n_98),
.Y(n_127)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_82),
.B(n_83),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_42),
.B(n_26),
.C(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_0),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_41),
.B1(n_27),
.B2(n_32),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_33),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_31),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_35),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_95),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_39),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_63),
.A2(n_26),
.B1(n_19),
.B2(n_34),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_64),
.B(n_38),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_43),
.B1(n_39),
.B2(n_38),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_34),
.B1(n_31),
.B2(n_39),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_34),
.Y(n_119)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_43),
.Y(n_100)
);

OR2x4_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_43),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_12),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_29),
.Y(n_129)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_120),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_85),
.B(n_94),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_72),
.B1(n_101),
.B2(n_80),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_11),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_126),
.A2(n_128),
.B1(n_131),
.B2(n_73),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_75),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_149),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_78),
.C(n_71),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_155),
.C(n_118),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_140),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_81),
.B1(n_74),
.B2(n_71),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_148),
.B1(n_157),
.B2(n_117),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_147),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_162),
.Y(n_185)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_108),
.A2(n_110),
.B1(n_128),
.B2(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_106),
.A2(n_83),
.B(n_85),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_156),
.B(n_132),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_78),
.B1(n_76),
.B2(n_87),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_113),
.B1(n_93),
.B2(n_124),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_125),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_153),
.A2(n_154),
.B1(n_158),
.B2(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_84),
.C(n_69),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_93),
.B1(n_75),
.B2(n_79),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_94),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_43),
.B1(n_65),
.B2(n_52),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_164),
.B(n_174),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_119),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_172),
.C(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_169),
.A2(n_192),
.B1(n_193),
.B2(n_3),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_176),
.B(n_177),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_175),
.B(n_179),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_112),
.B(n_123),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_122),
.B(n_120),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_181),
.B1(n_184),
.B2(n_179),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_111),
.B(n_105),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_186),
.B(n_163),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_136),
.A2(n_105),
.B1(n_93),
.B2(n_98),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_149),
.C(n_135),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_142),
.C(n_144),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_156),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_98),
.B1(n_102),
.B2(n_104),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_103),
.B(n_29),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_161),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_9),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_137),
.A2(n_98),
.B1(n_124),
.B2(n_34),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_139),
.A2(n_92),
.B1(n_39),
.B2(n_65),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_137),
.A2(n_43),
.B1(n_29),
.B2(n_1),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_199),
.B1(n_215),
.B2(n_173),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_177),
.B(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_205),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_160),
.B1(n_153),
.B2(n_138),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_210),
.B1(n_212),
.B2(n_216),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_214),
.C(n_218),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_176),
.A2(n_142),
.B1(n_140),
.B2(n_143),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_217),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_143),
.B1(n_29),
.B2(n_1),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_2),
.C(n_3),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_180),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_220),
.A2(n_224),
.B1(n_227),
.B2(n_215),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_205),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_204),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_172),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_228),
.C(n_233),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_198),
.B(n_185),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_197),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_237),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_170),
.B1(n_188),
.B2(n_174),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_185),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_216),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_181),
.B(n_169),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_231),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_192),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_203),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_167),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_241),
.Y(n_256)
);

BUFx12_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_251),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_208),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_233),
.C(n_214),
.Y(n_263)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_219),
.B(n_211),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_250),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_201),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_234),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_254),
.B1(n_226),
.B2(n_235),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_207),
.B1(n_196),
.B2(n_213),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_235),
.B1(n_196),
.B2(n_227),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_230),
.C(n_222),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_257),
.C(n_259),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_230),
.C(n_243),
.Y(n_257)
);

OAI211xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_206),
.B(n_231),
.C(n_224),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_242),
.B(n_266),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_208),
.C(n_228),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_267),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_264),
.C(n_195),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_214),
.C(n_210),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_241),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_271),
.Y(n_282)
);

NOR2x1_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_240),
.Y(n_269)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_270),
.B(n_6),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_257),
.Y(n_271)
);

OAI221xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_253),
.B1(n_240),
.B2(n_212),
.C(n_194),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_273),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_252),
.C(n_248),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_276),
.B(n_5),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_195),
.B(n_193),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_278),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_4),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_4),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_7),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_4),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_285),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_284),
.C(n_7),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_5),
.B(n_6),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_279),
.A2(n_280),
.B1(n_274),
.B2(n_285),
.Y(n_287)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_291),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_292),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_272),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_268),
.C(n_9),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_7),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_10),
.B(n_13),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g297 ( 
.A1(n_295),
.A2(n_289),
.A3(n_10),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_9),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_298),
.Y(n_299)
);

AOI321xp33_ASAP7_75t_SL g300 ( 
.A1(n_299),
.A2(n_294),
.A3(n_293),
.B1(n_296),
.B2(n_14),
.C(n_15),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_15),
.Y(n_301)
);


endmodule