module fake_jpeg_22408_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_42),
.Y(n_46)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_40),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_29),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_26),
.B1(n_25),
.B2(n_36),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_30),
.B1(n_29),
.B2(n_23),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_52),
.B1(n_36),
.B2(n_32),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_25),
.B(n_31),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_54),
.B(n_60),
.C(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_30),
.B1(n_27),
.B2(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_21),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_33),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_67),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_80),
.B1(n_85),
.B2(n_49),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_1),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_72),
.C(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_70),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_74),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_55),
.B1(n_47),
.B2(n_43),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_16),
.B1(n_33),
.B2(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_41),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_18),
.B(n_14),
.Y(n_100)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_49),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_55),
.B(n_43),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_106),
.B(n_86),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_92),
.A2(n_98),
.B1(n_101),
.B2(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_2),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_64),
.B1(n_77),
.B2(n_73),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_2),
.B(n_3),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_63),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_116),
.B(n_119),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_74),
.C(n_68),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_104),
.C(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_67),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_89),
.B(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_83),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.C(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_76),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_96),
.B1(n_91),
.B2(n_101),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_130),
.B1(n_116),
.B2(n_122),
.Y(n_143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_95),
.B(n_104),
.C(n_100),
.D(n_106),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_129),
.C(n_132),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_94),
.C(n_105),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_94),
.C(n_90),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_140),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_142),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_112),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_147),
.B1(n_132),
.B2(n_134),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_114),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_146),
.B(n_114),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_121),
.B(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_107),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_144),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_127),
.B(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_150),
.Y(n_160)
);

NAND4xp25_ASAP7_75t_SL g150 ( 
.A(n_142),
.B(n_102),
.C(n_133),
.D(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_110),
.C(n_108),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_140),
.B(n_128),
.C(n_117),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_158),
.Y(n_162)
);

OAI21x1_ASAP7_75t_SL g163 ( 
.A1(n_157),
.A2(n_159),
.B(n_153),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_149),
.B(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_128),
.B1(n_62),
.B2(n_76),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_164),
.B(n_166),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_154),
.B(n_151),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_4),
.C(n_5),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_165),
.B(n_5),
.Y(n_168)
);

AOI321xp33_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_161),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_159),
.C(n_7),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_169),
.A2(n_9),
.B(n_167),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_9),
.B(n_170),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_172),
.Y(n_173)
);


endmodule