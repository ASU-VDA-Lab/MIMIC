module real_jpeg_24757_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_288;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_1),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_1),
.A2(n_31),
.B1(n_56),
.B2(n_57),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_1),
.A2(n_31),
.B1(n_53),
.B2(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_2),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_28),
.B1(n_56),
.B2(n_57),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_2),
.A2(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_2),
.A2(n_60),
.B(n_164),
.C(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_2),
.B(n_55),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_2),
.A2(n_57),
.B(n_72),
.C(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_2),
.B(n_26),
.C(n_38),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_2),
.B(n_129),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_2),
.B(n_21),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_2),
.B(n_36),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_43),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_7),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_64),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_64),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_64),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_275),
.B1(n_288),
.B2(n_289),
.Y(n_13)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_14),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_133),
.B(n_274),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_110),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_16),
.B(n_110),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_81),
.C(n_89),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_17),
.B(n_81),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_48),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_18),
.B(n_49),
.C(n_68),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_34),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_19),
.B(n_34),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_20),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_24),
.A2(n_32),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_24),
.B(n_32),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_26),
.B(n_230),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_28),
.A2(n_57),
.B(n_59),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_28),
.A2(n_40),
.B(n_74),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_29),
.A2(n_93),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_29),
.B(n_223),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_32),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_32),
.B(n_217),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_33),
.Y(n_167)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_33),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B(n_44),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_35),
.B(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_35),
.A2(n_86),
.B(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_36),
.B(n_47),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_36),
.B(n_193),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_39),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_41),
.B1(n_72),
.B2(n_74),
.Y(n_71)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_41),
.B(n_206),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_44),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_44),
.B(n_203),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_45),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_45),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_67),
.B2(n_68),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_61),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_55),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_52),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_52),
.B(n_65),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_66)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_62),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_55),
.B(n_107),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_57),
.B1(n_72),
.B2(n_74),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_61),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_63),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_65),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_75),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_69),
.B(n_155),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_69),
.A2(n_77),
.B(n_128),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_70),
.B(n_78),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_78),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_71),
.B(n_103),
.Y(n_157)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_76),
.B(n_148),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_78),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_82),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_85),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_88),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_82),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_82),
.A2(n_88),
.B1(n_188),
.B2(n_246),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g285 ( 
.A1(n_82),
.A2(n_114),
.B(n_116),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_87),
.B(n_192),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_89),
.B(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_102),
.C(n_104),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_90),
.A2(n_91),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_92),
.B(n_99),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_95),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_95),
.B(n_216),
.Y(n_235)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_100),
.B(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_102),
.A2(n_104),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_102),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_104),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_132),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_121),
.B2(n_122),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_112),
.B(n_122),
.C(n_132),
.Y(n_286)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_127),
.B(n_131),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_127),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_124),
.B(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B(n_130),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_130),
.B(n_147),
.Y(n_146)
);

FAx1_ASAP7_75t_L g277 ( 
.A(n_131),
.B(n_278),
.CI(n_285),
.CON(n_277),
.SN(n_277)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_269),
.B(n_273),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_181),
.B(n_255),
.C(n_268),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_169),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_136),
.B(n_169),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_152),
.B2(n_168),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_150),
.B2(n_151),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_139),
.B(n_151),
.C(n_168),
.Y(n_256)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_146),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_142),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_143),
.B(n_159),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_144),
.A2(n_145),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_162),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_154),
.B(n_161),
.C(n_162),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_166),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.C(n_176),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_171),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_176),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.C(n_179),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_180),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_254),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_197),
.B(n_253),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_194),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_184),
.B(n_194),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_190),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_187),
.B(n_190),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_188),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_248),
.B(n_252),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_239),
.B(n_247),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_220),
.B(n_238),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_201),
.B(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_214),
.B2(n_219),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_210),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_213),
.C(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_227),
.B(n_237),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_222),
.B(n_225),
.Y(n_237)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_236),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_234),
.B(n_235),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_241),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_244),
.C(n_245),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_256),
.B(n_257),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_267),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_265),
.B2(n_266),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_266),
.C(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_287),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_286),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_286),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_277),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_280),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);


endmodule