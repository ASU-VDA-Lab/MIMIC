module fake_ariane_3295_n_1567 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_439, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_432, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_429, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_438, n_314, n_16, n_440, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_430, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_428, n_159, n_358, n_105, n_30, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_425, n_431, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_1567);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_439;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_432;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_429;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_430;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_425;
input n_431;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_1567;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_1495;
wire n_661;
wire n_533;
wire n_1560;
wire n_1548;
wire n_1396;
wire n_1230;
wire n_612;
wire n_512;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_551;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_1521;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_519;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_1552;
wire n_750;
wire n_834;
wire n_800;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_975;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1458;
wire n_679;
wire n_663;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_504;
wire n_483;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_946;
wire n_757;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_1228;
wire n_1244;
wire n_484;
wire n_849;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g444 ( 
.A(n_247),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_266),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_359),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_7),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_101),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_379),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_8),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_25),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_82),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_7),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_186),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_65),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_102),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_54),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_160),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_122),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_12),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_361),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_124),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_194),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_424),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_423),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_253),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_156),
.Y(n_467)
);

BUFx5_ASAP7_75t_L g468 ( 
.A(n_356),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_432),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_50),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_15),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_184),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_317),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_140),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_63),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_350),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_409),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_158),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_119),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_115),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_89),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_162),
.Y(n_482)
);

BUFx2_ASAP7_75t_SL g483 ( 
.A(n_118),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_360),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_129),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_126),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_342),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_183),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_134),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_27),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_281),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_311),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_296),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_205),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_305),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_380),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_100),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_337),
.Y(n_498)
);

BUFx10_ASAP7_75t_L g499 ( 
.A(n_31),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_413),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_64),
.Y(n_501)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_288),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_255),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_386),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_382),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_121),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_127),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_370),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_353),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_79),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_146),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_107),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_259),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_123),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_128),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_120),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_75),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_19),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_80),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_419),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_91),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_291),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_180),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_242),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_295),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_63),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_275),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_143),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_144),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_349),
.Y(n_530)
);

CKINVDCx14_ASAP7_75t_R g531 ( 
.A(n_431),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_358),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_216),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_10),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_147),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_103),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_264),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_57),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_289),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_222),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_322),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_403),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_200),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_42),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_221),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_130),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_274),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_88),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_307),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_411),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_195),
.B(n_265),
.Y(n_551)
);

BUFx5_ASAP7_75t_L g552 ( 
.A(n_142),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_300),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_430),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_174),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_283),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_37),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_206),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_20),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_323),
.Y(n_561)
);

INVxp67_ASAP7_75t_SL g562 ( 
.A(n_250),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_202),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_290),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_327),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_23),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_6),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_85),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_154),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_324),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_282),
.B(n_81),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_277),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_40),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g574 ( 
.A(n_209),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_190),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_319),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_85),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_59),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_381),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_0),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_65),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_19),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_131),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_104),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_29),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_197),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_95),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_215),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_315),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_410),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_88),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_387),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_18),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_188),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_106),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_212),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_157),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_66),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_278),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_13),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_376),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_125),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_240),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_383),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_402),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_2),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_239),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_28),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_417),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_6),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_316),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_344),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_0),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_79),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_165),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_241),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_30),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_166),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_318),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_47),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_152),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_91),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_231),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_81),
.Y(n_624)
);

CKINVDCx14_ASAP7_75t_R g625 ( 
.A(n_301),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_364),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_326),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_204),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_207),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_201),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_519),
.B(n_566),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_492),
.Y(n_632)
);

CKINVDCx6p67_ASAP7_75t_R g633 ( 
.A(n_572),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_560),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_560),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_469),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_595),
.B(n_1),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_560),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_452),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_560),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_582),
.Y(n_641)
);

BUFx8_ASAP7_75t_SL g642 ( 
.A(n_536),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_492),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_472),
.A2(n_3),
.B1(n_1),
.B2(n_2),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_492),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_492),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_608),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_582),
.Y(n_648)
);

OAI22x1_ASAP7_75t_R g649 ( 
.A1(n_448),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_523),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_523),
.Y(n_651)
);

NOR2x1_ASAP7_75t_L g652 ( 
.A(n_509),
.B(n_111),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_581),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_542),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_581),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_542),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_542),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_582),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_625),
.A2(n_574),
.B1(n_531),
.B2(n_502),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_622),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_542),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_599),
.B(n_112),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_506),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_506),
.Y(n_664)
);

BUFx12f_ASAP7_75t_L g665 ( 
.A(n_499),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_556),
.B(n_4),
.Y(n_666)
);

OA21x2_ASAP7_75t_L g667 ( 
.A1(n_444),
.A2(n_466),
.B(n_463),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_SL g668 ( 
.A1(n_584),
.A2(n_9),
.B1(n_5),
.B2(n_8),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_480),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_484),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_556),
.B(n_9),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_629),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_622),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_485),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_622),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_629),
.Y(n_676)
);

BUFx8_ASAP7_75t_L g677 ( 
.A(n_590),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_629),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_447),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_629),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_491),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_455),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_599),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_621),
.B(n_10),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_451),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_460),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_475),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_481),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_515),
.A2(n_114),
.B(n_113),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_497),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_501),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_450),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_584),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_521),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_453),
.B(n_11),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_591),
.Y(n_696)
);

BUFx12f_ASAP7_75t_L g697 ( 
.A(n_499),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_456),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_580),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_522),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_598),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_543),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_498),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_473),
.B(n_11),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_600),
.Y(n_705)
);

AOI22x1_ASAP7_75t_SL g706 ( 
.A1(n_516),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_610),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_474),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_476),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_587),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_457),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_517),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_632),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_632),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_632),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_643),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_671),
.B(n_459),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_643),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_SL g719 ( 
.A(n_671),
.B(n_615),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_683),
.B(n_625),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_640),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_651),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_643),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_659),
.B(n_520),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_640),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_683),
.B(n_477),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_670),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_645),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_636),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_645),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_651),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_686),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_662),
.Y(n_733)
);

INVxp33_ASAP7_75t_L g734 ( 
.A(n_685),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_631),
.B(n_478),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_687),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_658),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_658),
.Y(n_738)
);

AOI21x1_ASAP7_75t_L g739 ( 
.A1(n_667),
.A2(n_488),
.B(n_486),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_690),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_674),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_654),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_663),
.B(n_664),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_698),
.B(n_562),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_634),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_647),
.B(n_517),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_712),
.B(n_547),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_662),
.Y(n_748)
);

AND3x2_ASAP7_75t_L g749 ( 
.A(n_666),
.B(n_562),
.C(n_569),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_684),
.B(n_594),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_639),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_669),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_660),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_660),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_682),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_654),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_682),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_673),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_635),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_722),
.B(n_667),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_755),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_757),
.A2(n_693),
.B(n_704),
.C(n_691),
.Y(n_762)
);

BUFx6f_ASAP7_75t_SL g763 ( 
.A(n_727),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_741),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_741),
.B(n_727),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_751),
.B(n_734),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_742),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_744),
.B(n_726),
.C(n_709),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_722),
.B(n_708),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_731),
.B(n_708),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_719),
.A2(n_644),
.B1(n_637),
.B2(n_633),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_751),
.B(n_711),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_746),
.B(n_637),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_721),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_720),
.B(n_731),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_724),
.B(n_665),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_746),
.B(n_653),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_732),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_736),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_719),
.B(n_695),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_743),
.B(n_695),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_717),
.A2(n_750),
.B1(n_747),
.B2(n_735),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_749),
.A2(n_623),
.B1(n_573),
.B2(n_740),
.Y(n_783)
);

AO221x1_ASAP7_75t_L g784 ( 
.A1(n_745),
.A2(n_668),
.B1(n_649),
.B2(n_706),
.C(n_647),
.Y(n_784)
);

BUFx5_ASAP7_75t_L g785 ( 
.A(n_733),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_725),
.B(n_662),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_725),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_733),
.B(n_681),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_733),
.B(n_703),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_737),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_742),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_748),
.B(n_571),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_748),
.B(n_677),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_729),
.B(n_655),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_729),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_737),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_748),
.B(n_677),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_748),
.B(n_697),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_752),
.B(n_445),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_738),
.B(n_700),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_753),
.B(n_700),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_752),
.B(n_700),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_742),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_753),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_754),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_754),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_758),
.B(n_702),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_758),
.B(n_702),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_739),
.B(n_702),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_745),
.B(n_646),
.Y(n_810)
);

NOR3xp33_ASAP7_75t_L g811 ( 
.A(n_759),
.B(n_471),
.C(n_470),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_713),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_739),
.B(n_638),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_713),
.B(n_641),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_714),
.B(n_648),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_715),
.Y(n_816)
);

NOR3xp33_ASAP7_75t_L g817 ( 
.A(n_715),
.B(n_510),
.C(n_490),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_716),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_716),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_718),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_742),
.B(n_512),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_718),
.B(n_518),
.Y(n_822)
);

OR2x2_ASAP7_75t_L g823 ( 
.A(n_723),
.B(n_692),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_723),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_728),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_728),
.B(n_688),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_756),
.A2(n_534),
.B1(n_538),
.B2(n_526),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_730),
.B(n_691),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_766),
.B(n_692),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_768),
.B(n_544),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_823),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_768),
.B(n_454),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_767),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_780),
.B(n_642),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_775),
.A2(n_689),
.B(n_494),
.Y(n_835)
);

BUFx2_ASAP7_75t_L g836 ( 
.A(n_794),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_795),
.B(n_548),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_764),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_776),
.B(n_558),
.Y(n_839)
);

AOI21xp33_ASAP7_75t_L g840 ( 
.A1(n_762),
.A2(n_568),
.B(n_567),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_777),
.B(n_577),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_773),
.B(n_500),
.Y(n_842)
);

O2A1O1Ixp5_ASAP7_75t_L g843 ( 
.A1(n_786),
.A2(n_761),
.B(n_770),
.C(n_769),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_796),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_816),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_778),
.B(n_525),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_804),
.A2(n_805),
.B(n_774),
.C(n_787),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_781),
.B(n_540),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_771),
.A2(n_483),
.B1(n_528),
.B2(n_527),
.Y(n_849)
);

AND2x4_ASAP7_75t_SL g850 ( 
.A(n_765),
.B(n_772),
.Y(n_850)
);

A2O1A1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_790),
.A2(n_530),
.B(n_535),
.C(n_532),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_779),
.B(n_578),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_760),
.A2(n_553),
.B(n_550),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_813),
.A2(n_565),
.B(n_557),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_765),
.B(n_585),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_782),
.B(n_546),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_765),
.B(n_593),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_806),
.B(n_559),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_767),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_788),
.B(n_606),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_826),
.A2(n_592),
.B(n_597),
.C(n_586),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_800),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_783),
.B(n_613),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_799),
.B(n_617),
.C(n_614),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_801),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_810),
.A2(n_652),
.B(n_551),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_793),
.B(n_679),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_789),
.B(n_620),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_797),
.B(n_701),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_802),
.B(n_699),
.Y(n_870)
);

OAI21xp33_ASAP7_75t_L g871 ( 
.A1(n_827),
.A2(n_624),
.B(n_811),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_763),
.Y(n_872)
);

AO22x1_ASAP7_75t_L g873 ( 
.A1(n_784),
.A2(n_705),
.B1(n_696),
.B2(n_694),
.Y(n_873)
);

INVx5_ASAP7_75t_L g874 ( 
.A(n_767),
.Y(n_874)
);

OR2x6_ASAP7_75t_L g875 ( 
.A(n_798),
.B(n_707),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_820),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_763),
.A2(n_604),
.B1(n_605),
.B2(n_601),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_828),
.B(n_446),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_808),
.Y(n_879)
);

AO21x1_ASAP7_75t_L g880 ( 
.A1(n_792),
.A2(n_618),
.B(n_616),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_814),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_817),
.A2(n_675),
.B(n_673),
.C(n_630),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_824),
.B(n_449),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_825),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_SL g885 ( 
.A(n_821),
.B(n_458),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_807),
.Y(n_886)
);

AOI211xp5_ASAP7_75t_L g887 ( 
.A1(n_822),
.A2(n_710),
.B(n_628),
.C(n_699),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_791),
.B(n_819),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_812),
.B(n_461),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_818),
.B(n_462),
.Y(n_890)
);

OAI21xp33_ASAP7_75t_L g891 ( 
.A1(n_815),
.A2(n_465),
.B(n_464),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_785),
.B(n_467),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_803),
.B(n_479),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_803),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_785),
.B(n_482),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_785),
.B(n_487),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_768),
.B(n_489),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_768),
.B(n_493),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_768),
.B(n_495),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_768),
.A2(n_503),
.B1(n_504),
.B2(n_496),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_765),
.B(n_549),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_768),
.B(n_505),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_767),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_775),
.A2(n_756),
.B(n_508),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_764),
.Y(n_905)
);

INVx11_ASAP7_75t_L g906 ( 
.A(n_763),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_766),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_766),
.B(n_507),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_775),
.A2(n_513),
.B(n_511),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_823),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_768),
.B(n_514),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_766),
.B(n_524),
.Y(n_912)
);

A2O1A1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_768),
.A2(n_555),
.B(n_554),
.C(n_533),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_SL g914 ( 
.A(n_766),
.B(n_529),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_780),
.A2(n_537),
.B1(n_541),
.B2(n_539),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_768),
.B(n_545),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_763),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_809),
.A2(n_657),
.B(n_650),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_761),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_766),
.B(n_561),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_823),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_768),
.B(n_563),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_763),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_786),
.A2(n_570),
.B(n_564),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_775),
.A2(n_576),
.B(n_575),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_816),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_768),
.B(n_579),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_765),
.B(n_16),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_764),
.B(n_650),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_777),
.A2(n_588),
.B(n_583),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_892),
.A2(n_596),
.B(n_589),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_843),
.A2(n_603),
.B(n_602),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_918),
.A2(n_552),
.B(n_468),
.Y(n_933)
);

OR2x4_ASAP7_75t_L g934 ( 
.A(n_855),
.B(n_17),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_839),
.B(n_607),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_917),
.B(n_650),
.Y(n_936)
);

CKINVDCx20_ASAP7_75t_R g937 ( 
.A(n_836),
.Y(n_937)
);

OAI21xp5_ASAP7_75t_L g938 ( 
.A1(n_847),
.A2(n_611),
.B(n_609),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_908),
.B(n_612),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_850),
.B(n_829),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_838),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_912),
.B(n_619),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_895),
.A2(n_627),
.B(n_626),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_924),
.A2(n_672),
.B(n_657),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_907),
.B(n_17),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_896),
.A2(n_672),
.B(n_657),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_904),
.A2(n_916),
.B(n_899),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_920),
.B(n_18),
.Y(n_948)
);

BUFx12f_ASAP7_75t_L g949 ( 
.A(n_917),
.Y(n_949)
);

OAI22x1_ASAP7_75t_L g950 ( 
.A1(n_849),
.A2(n_672),
.B1(n_22),
.B2(n_20),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_857),
.B(n_21),
.Y(n_951)
);

AND3x4_ASAP7_75t_L g952 ( 
.A(n_928),
.B(n_21),
.C(n_22),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_844),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_923),
.B(n_654),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_888),
.A2(n_661),
.B(n_656),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_832),
.B(n_24),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_853),
.A2(n_117),
.B(n_116),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_862),
.B(n_26),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_865),
.B(n_879),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_856),
.B(n_846),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_928),
.Y(n_961)
);

AO31x2_ASAP7_75t_L g962 ( 
.A1(n_880),
.A2(n_678),
.A3(n_680),
.B(n_676),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_854),
.A2(n_678),
.B(n_676),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_833),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_869),
.B(n_26),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_897),
.A2(n_902),
.B(n_911),
.C(n_898),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_906),
.Y(n_967)
);

OAI21x1_ASAP7_75t_SL g968 ( 
.A1(n_919),
.A2(n_27),
.B(n_28),
.Y(n_968)
);

AO31x2_ASAP7_75t_L g969 ( 
.A1(n_861),
.A2(n_680),
.A3(n_678),
.B(n_31),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_914),
.B(n_29),
.Y(n_970)
);

NOR2xp67_ASAP7_75t_L g971 ( 
.A(n_923),
.B(n_132),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_905),
.B(n_30),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_929),
.Y(n_973)
);

INVxp67_ASAP7_75t_SL g974 ( 
.A(n_833),
.Y(n_974)
);

OAI21x1_ASAP7_75t_L g975 ( 
.A1(n_866),
.A2(n_876),
.B(n_867),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_876),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_878),
.A2(n_680),
.B(n_133),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_840),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_922),
.A2(n_136),
.B(n_135),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_927),
.A2(n_138),
.B(n_137),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_860),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_869),
.B(n_35),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_909),
.A2(n_141),
.B(n_139),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_925),
.A2(n_148),
.B(n_145),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_894),
.A2(n_150),
.B(n_149),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_913),
.A2(n_153),
.B(n_151),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_845),
.B(n_35),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_901),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_926),
.B(n_36),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_926),
.B(n_36),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_834),
.B(n_37),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_910),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_833),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_858),
.B(n_38),
.Y(n_994)
);

AND3x4_ASAP7_75t_L g995 ( 
.A(n_864),
.B(n_39),
.C(n_40),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_889),
.A2(n_159),
.B(n_155),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_872),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_901),
.B(n_39),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_831),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_883),
.B(n_41),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_890),
.A2(n_163),
.B(n_161),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_921),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_SL g1003 ( 
.A1(n_893),
.A2(n_167),
.B(n_164),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_870),
.B(n_841),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_882),
.A2(n_169),
.B(n_168),
.Y(n_1005)
);

BUFx10_ASAP7_75t_L g1006 ( 
.A(n_868),
.Y(n_1006)
);

NAND2x1p5_ASAP7_75t_L g1007 ( 
.A(n_874),
.B(n_41),
.Y(n_1007)
);

AND2x2_ASAP7_75t_SL g1008 ( 
.A(n_848),
.B(n_42),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_859),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_842),
.B(n_43),
.Y(n_1010)
);

AO31x2_ASAP7_75t_L g1011 ( 
.A1(n_851),
.A2(n_46),
.A3(n_44),
.B(n_45),
.Y(n_1011)
);

AOI21x1_ASAP7_75t_L g1012 ( 
.A1(n_852),
.A2(n_171),
.B(n_170),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_930),
.B(n_44),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_884),
.B(n_871),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_891),
.A2(n_173),
.B(n_172),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_915),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_SL g1017 ( 
.A1(n_877),
.A2(n_48),
.B(n_49),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_886),
.B(n_50),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_885),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_837),
.A2(n_176),
.B(n_175),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_863),
.B(n_51),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_900),
.B(n_52),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_859),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_903),
.B(n_887),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_875),
.B(n_54),
.Y(n_1025)
);

AOI21x1_ASAP7_75t_L g1026 ( 
.A1(n_875),
.A2(n_178),
.B(n_177),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_873),
.A2(n_181),
.B(n_179),
.Y(n_1027)
);

AOI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_839),
.A2(n_55),
.B(n_56),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_833),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_839),
.B(n_55),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_892),
.A2(n_185),
.B(n_182),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_917),
.B(n_56),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_892),
.A2(n_189),
.B(n_187),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_844),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_833),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_SL g1036 ( 
.A1(n_924),
.A2(n_58),
.B(n_60),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_917),
.B(n_61),
.Y(n_1037)
);

OAI22x1_ASAP7_75t_L g1038 ( 
.A1(n_849),
.A2(n_66),
.B1(n_62),
.B2(n_64),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_839),
.B(n_62),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_843),
.A2(n_192),
.B(n_191),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_835),
.A2(n_196),
.B(n_193),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_L g1042 ( 
.A(n_839),
.B(n_67),
.C(n_68),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_892),
.A2(n_199),
.B(n_198),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_844),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_839),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_833),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_836),
.B(n_70),
.Y(n_1047)
);

AO31x2_ASAP7_75t_L g1048 ( 
.A1(n_880),
.A2(n_73),
.A3(n_71),
.B(n_72),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_835),
.A2(n_208),
.B(n_203),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_892),
.A2(n_211),
.B(n_210),
.Y(n_1050)
);

O2A1O1Ixp5_ASAP7_75t_L g1051 ( 
.A1(n_899),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_835),
.A2(n_214),
.B(n_213),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_838),
.Y(n_1053)
);

AOI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_839),
.A2(n_74),
.B(n_75),
.Y(n_1054)
);

OAI21x1_ASAP7_75t_L g1055 ( 
.A1(n_835),
.A2(n_218),
.B(n_217),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_843),
.A2(n_220),
.B(n_219),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_835),
.A2(n_224),
.B(n_223),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_L g1058 ( 
.A1(n_839),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.C(n_80),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_843),
.A2(n_226),
.B(n_225),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_836),
.B(n_76),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_833),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_892),
.A2(n_228),
.B(n_227),
.Y(n_1062)
);

AOI211x1_ASAP7_75t_L g1063 ( 
.A1(n_830),
.A2(n_77),
.B(n_78),
.C(n_82),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_836),
.B(n_83),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_843),
.A2(n_230),
.B(n_229),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_917),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_881),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_843),
.A2(n_233),
.B(n_232),
.Y(n_1068)
);

BUFx4f_ASAP7_75t_SL g1069 ( 
.A(n_917),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_892),
.A2(n_235),
.B(n_234),
.Y(n_1070)
);

OA22x2_ASAP7_75t_L g1071 ( 
.A1(n_836),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_918),
.A2(n_237),
.B(n_236),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_SL g1073 ( 
.A(n_874),
.B(n_238),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_850),
.Y(n_1074)
);

OAI22x1_ASAP7_75t_L g1075 ( 
.A1(n_849),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_881),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_843),
.A2(n_244),
.B(n_243),
.Y(n_1077)
);

NAND3xp33_ASAP7_75t_SL g1078 ( 
.A(n_839),
.B(n_92),
.C(n_93),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_843),
.A2(n_246),
.B(n_245),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_839),
.B(n_94),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_836),
.B(n_94),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_L g1082 ( 
.A1(n_899),
.A2(n_95),
.B(n_96),
.C(n_97),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_960),
.B(n_96),
.Y(n_1083)
);

BUFx2_ASAP7_75t_R g1084 ( 
.A(n_997),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_961),
.B(n_97),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1067),
.Y(n_1086)
);

AO21x2_ASAP7_75t_L g1087 ( 
.A1(n_932),
.A2(n_249),
.B(n_248),
.Y(n_1087)
);

AO21x2_ASAP7_75t_L g1088 ( 
.A1(n_1040),
.A2(n_252),
.B(n_251),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1067),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_937),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1076),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_SL g1092 ( 
.A1(n_1036),
.A2(n_98),
.B(n_99),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1076),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_959),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_941),
.B(n_98),
.Y(n_1095)
);

CKINVDCx6p67_ASAP7_75t_R g1096 ( 
.A(n_1066),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_966),
.A2(n_100),
.B(n_101),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1006),
.B(n_102),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_999),
.Y(n_1099)
);

AO21x2_ASAP7_75t_L g1100 ( 
.A1(n_1056),
.A2(n_256),
.B(n_254),
.Y(n_1100)
);

NAND2x1p5_ASAP7_75t_L g1101 ( 
.A(n_1053),
.B(n_257),
.Y(n_1101)
);

AO21x1_ASAP7_75t_SL g1102 ( 
.A1(n_1030),
.A2(n_103),
.B(n_104),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_999),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1008),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_935),
.A2(n_1039),
.B1(n_1080),
.B2(n_948),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_947),
.A2(n_351),
.A3(n_442),
.B(n_441),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_1074),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_956),
.A2(n_105),
.B(n_108),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1002),
.Y(n_1109)
);

AND2x4_ASAP7_75t_L g1110 ( 
.A(n_1066),
.B(n_108),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_940),
.Y(n_1111)
);

NOR2xp67_ASAP7_75t_SL g1112 ( 
.A(n_967),
.B(n_109),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_998),
.B(n_110),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1006),
.B(n_258),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_949),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_998),
.B(n_260),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_976),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1047),
.B(n_261),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_933),
.A2(n_262),
.B(n_263),
.Y(n_1119)
);

AO21x2_ASAP7_75t_L g1120 ( 
.A1(n_1059),
.A2(n_267),
.B(n_268),
.Y(n_1120)
);

OAI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_970),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.C(n_272),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_992),
.A2(n_273),
.B1(n_276),
.B2(n_279),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_951),
.B(n_280),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_1069),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_972),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_939),
.B(n_284),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1004),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_SL g1128 ( 
.A1(n_1073),
.A2(n_292),
.B(n_293),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_1066),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1041),
.A2(n_294),
.B(n_297),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_1065),
.A2(n_298),
.B(n_299),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_1060),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_964),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_964),
.Y(n_1134)
);

AO21x2_ASAP7_75t_L g1135 ( 
.A1(n_1068),
.A2(n_302),
.B(n_303),
.Y(n_1135)
);

BUFx4f_ASAP7_75t_SL g1136 ( 
.A(n_967),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1049),
.A2(n_304),
.B(n_306),
.Y(n_1137)
);

BUFx12f_ASAP7_75t_L g1138 ( 
.A(n_1032),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1052),
.A2(n_308),
.B(n_309),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_988),
.B(n_310),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1064),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1081),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_973),
.B(n_312),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_958),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_964),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_975),
.Y(n_1146)
);

CKINVDCx11_ASAP7_75t_R g1147 ( 
.A(n_1032),
.Y(n_1147)
);

OA21x2_ASAP7_75t_L g1148 ( 
.A1(n_1077),
.A2(n_313),
.B(n_314),
.Y(n_1148)
);

AO21x2_ASAP7_75t_L g1149 ( 
.A1(n_1079),
.A2(n_320),
.B(n_321),
.Y(n_1149)
);

BUFx2_ASAP7_75t_R g1150 ( 
.A(n_965),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1037),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_993),
.B(n_325),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1037),
.Y(n_1153)
);

OA21x2_ASAP7_75t_L g1154 ( 
.A1(n_1055),
.A2(n_328),
.B(n_329),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1057),
.A2(n_330),
.B(n_331),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_SL g1156 ( 
.A1(n_1073),
.A2(n_1022),
.B(n_986),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_945),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_942),
.B(n_332),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_989),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_990),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1072),
.A2(n_333),
.B(n_334),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_982),
.B(n_335),
.Y(n_1162)
);

INVxp67_ASAP7_75t_SL g1163 ( 
.A(n_1029),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_991),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1001),
.A2(n_336),
.B(n_338),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_SL g1166 ( 
.A1(n_1000),
.A2(n_339),
.B(n_340),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_934),
.Y(n_1167)
);

AO21x2_ASAP7_75t_L g1168 ( 
.A1(n_944),
.A2(n_341),
.B(n_343),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1014),
.B(n_345),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1010),
.B(n_346),
.Y(n_1170)
);

BUFx2_ASAP7_75t_SL g1171 ( 
.A(n_971),
.Y(n_1171)
);

NAND3xp33_ASAP7_75t_L g1172 ( 
.A(n_1028),
.B(n_347),
.C(n_348),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_1025),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_1029),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1029),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1023),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_954),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1061),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_955),
.A2(n_352),
.A3(n_354),
.B(n_355),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_957),
.A2(n_357),
.B(n_362),
.Y(n_1180)
);

INVx6_ASAP7_75t_L g1181 ( 
.A(n_952),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1061),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1071),
.B(n_443),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1061),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1031),
.A2(n_363),
.B(n_365),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_993),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_969),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1033),
.A2(n_366),
.B(n_367),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_969),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_994),
.A2(n_931),
.B(n_1013),
.Y(n_1190)
);

AO21x2_ASAP7_75t_L g1191 ( 
.A1(n_963),
.A2(n_368),
.B(n_369),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1043),
.A2(n_371),
.B(n_372),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1021),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1050),
.A2(n_1070),
.B(n_1062),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1015),
.A2(n_373),
.A3(n_374),
.B(n_375),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_977),
.A2(n_377),
.B(n_378),
.Y(n_1196)
);

OA21x2_ASAP7_75t_L g1197 ( 
.A1(n_1005),
.A2(n_384),
.B(n_385),
.Y(n_1197)
);

NOR2xp67_ASAP7_75t_L g1198 ( 
.A(n_1035),
.B(n_388),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1046),
.B(n_389),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1018),
.B(n_390),
.Y(n_1200)
);

OAI21xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1058),
.A2(n_391),
.B(n_392),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1038),
.B(n_393),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1011),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_979),
.A2(n_394),
.B(n_395),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_980),
.A2(n_396),
.B(n_397),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_1007),
.B(n_398),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1024),
.B(n_399),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1046),
.Y(n_1208)
);

NOR2xp67_ASAP7_75t_L g1209 ( 
.A(n_1042),
.B(n_400),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1012),
.A2(n_401),
.B(n_404),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1075),
.B(n_405),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_983),
.A2(n_406),
.B(n_407),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_984),
.A2(n_408),
.B(n_412),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_996),
.A2(n_414),
.B(n_415),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1051),
.A2(n_418),
.B(n_420),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_962),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1026),
.A2(n_421),
.B(n_422),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_987),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_985),
.A2(n_425),
.B(n_426),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_950),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_974),
.B(n_427),
.Y(n_1221)
);

AO21x2_ASAP7_75t_L g1222 ( 
.A1(n_938),
.A2(n_428),
.B(n_429),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_SL g1223 ( 
.A1(n_953),
.A2(n_433),
.B1(n_434),
.B2(n_435),
.Y(n_1223)
);

INVx6_ASAP7_75t_L g1224 ( 
.A(n_995),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1009),
.B(n_436),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_936),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_946),
.A2(n_437),
.B(n_438),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1020),
.A2(n_439),
.B(n_440),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_962),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1027),
.A2(n_1082),
.B(n_1003),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1048),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1078),
.B(n_1054),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1017),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_968),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1048),
.Y(n_1235)
);

BUFx2_ASAP7_75t_R g1236 ( 
.A(n_1063),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_978),
.A2(n_943),
.B(n_1016),
.Y(n_1237)
);

AOI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1156),
.A2(n_1034),
.B(n_1044),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1109),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1097),
.A2(n_1201),
.B(n_1105),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1125),
.B(n_981),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1109),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1099),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1099),
.Y(n_1244)
);

AO21x2_ASAP7_75t_L g1245 ( 
.A1(n_1187),
.A2(n_1019),
.B(n_1045),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1103),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1134),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1103),
.Y(n_1248)
);

AOI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1146),
.A2(n_1194),
.B(n_1189),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_SL g1250 ( 
.A1(n_1220),
.A2(n_1181),
.B1(n_1211),
.B2(n_1202),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1094),
.B(n_1086),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1086),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1089),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1090),
.Y(n_1254)
);

CKINVDCx6p67_ASAP7_75t_R g1255 ( 
.A(n_1124),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1138),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1091),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1091),
.Y(n_1258)
);

CKINVDCx12_ASAP7_75t_R g1259 ( 
.A(n_1116),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1094),
.B(n_1093),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1093),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1117),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1141),
.B(n_1125),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1151),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1111),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1117),
.Y(n_1266)
);

AO21x1_ASAP7_75t_L g1267 ( 
.A1(n_1232),
.A2(n_1108),
.B(n_1190),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1104),
.A2(n_1183),
.B1(n_1193),
.B2(n_1144),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1136),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1174),
.Y(n_1270)
);

AOI221xp5_ASAP7_75t_L g1271 ( 
.A1(n_1095),
.A2(n_1098),
.B1(n_1201),
.B2(n_1164),
.C(n_1083),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1176),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1144),
.A2(n_1173),
.B1(n_1142),
.B2(n_1181),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1115),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1116),
.A2(n_1236),
.B1(n_1223),
.B2(n_1123),
.Y(n_1275)
);

OR2x6_ASAP7_75t_L g1276 ( 
.A(n_1153),
.B(n_1140),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_1174),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1237),
.A2(n_1160),
.B(n_1159),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1096),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1143),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1178),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1143),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1152),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1223),
.A2(n_1118),
.B1(n_1162),
.B2(n_1159),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1182),
.B(n_1184),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1225),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1224),
.A2(n_1113),
.B1(n_1157),
.B2(n_1110),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1175),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1203),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1203),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1180),
.A2(n_1165),
.B(n_1155),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1177),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1110),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1160),
.Y(n_1294)
);

NAND2x1p5_ASAP7_75t_L g1295 ( 
.A(n_1145),
.B(n_1186),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1186),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1130),
.A2(n_1137),
.B(n_1139),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1208),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1147),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1132),
.B(n_1150),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1085),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1162),
.A2(n_1224),
.B1(n_1222),
.B2(n_1206),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1215),
.A2(n_1126),
.B(n_1158),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1231),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1235),
.A2(n_1216),
.B(n_1230),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1167),
.B(n_1084),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1087),
.A2(n_1088),
.B(n_1135),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1107),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1133),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1218),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1163),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1226),
.B(n_1129),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1101),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1229),
.A2(n_1119),
.B(n_1210),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1234),
.B(n_1233),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1172),
.A2(n_1209),
.B(n_1200),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1206),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1106),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1112),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1209),
.A2(n_1170),
.B1(n_1148),
.B2(n_1131),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1199),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1092),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1102),
.B(n_1114),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1198),
.B(n_1207),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1221),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1106),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1198),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1171),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1229),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1172),
.A2(n_1169),
.B(n_1219),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1191),
.Y(n_1331)
);

NAND2x1p5_ASAP7_75t_L g1332 ( 
.A(n_1228),
.B(n_1148),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1127),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1212),
.A2(n_1213),
.B(n_1161),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1166),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1204),
.A2(n_1205),
.B(n_1192),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1185),
.A2(n_1188),
.B(n_1214),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1222),
.A2(n_1087),
.B1(n_1088),
.B2(n_1100),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1179),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1128),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1121),
.A2(n_1122),
.B1(n_1197),
.B2(n_1154),
.Y(n_1341)
);

OR2x6_ASAP7_75t_L g1342 ( 
.A(n_1217),
.B(n_1227),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1195),
.Y(n_1343)
);

CKINVDCx14_ASAP7_75t_R g1344 ( 
.A(n_1168),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1168),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1100),
.B(n_1120),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1263),
.B(n_1120),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1301),
.B(n_1135),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1273),
.B(n_1149),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1251),
.B(n_1260),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1273),
.B(n_1149),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1239),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1242),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1287),
.B(n_1154),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1252),
.Y(n_1355)
);

AO22x1_ASAP7_75t_L g1356 ( 
.A1(n_1275),
.A2(n_1284),
.B1(n_1333),
.B2(n_1240),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1252),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1287),
.B(n_1265),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1275),
.A2(n_1196),
.B1(n_1284),
.B2(n_1240),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1251),
.B(n_1260),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1253),
.B(n_1265),
.Y(n_1361)
);

BUFx12f_ASAP7_75t_L g1362 ( 
.A(n_1279),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1253),
.B(n_1254),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1264),
.B(n_1300),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1300),
.B(n_1250),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1268),
.A2(n_1271),
.B1(n_1250),
.B2(n_1267),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1271),
.A2(n_1268),
.B1(n_1302),
.B2(n_1283),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1281),
.B(n_1293),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1243),
.B(n_1244),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1288),
.B(n_1276),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1315),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1276),
.B(n_1294),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1259),
.A2(n_1276),
.B1(n_1317),
.B2(n_1241),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1302),
.A2(n_1241),
.B1(n_1344),
.B2(n_1323),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1262),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1246),
.B(n_1248),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1266),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1344),
.A2(n_1280),
.B1(n_1282),
.B2(n_1245),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1309),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1272),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1269),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1306),
.B(n_1308),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1311),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1292),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1286),
.A2(n_1261),
.B1(n_1258),
.B2(n_1257),
.Y(n_1385)
);

CKINVDCx11_ASAP7_75t_R g1386 ( 
.A(n_1255),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1285),
.B(n_1310),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1289),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1310),
.B(n_1256),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1298),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1292),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1290),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1299),
.B(n_1312),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1279),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1278),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1245),
.A2(n_1303),
.B1(n_1320),
.B2(n_1316),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1247),
.B(n_1279),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1322),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1325),
.B(n_1329),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1328),
.B(n_1319),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1274),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1313),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1304),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1321),
.B(n_1296),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1270),
.B(n_1277),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1303),
.A2(n_1320),
.B1(n_1316),
.B2(n_1338),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1305),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1321),
.Y(n_1408)
);

INVx5_ASAP7_75t_L g1409 ( 
.A(n_1296),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1249),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1327),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1295),
.B(n_1238),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1335),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1340),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1329),
.B(n_1324),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1324),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1346),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1357),
.B(n_1363),
.Y(n_1418)
);

OAI222xp33_ASAP7_75t_L g1419 ( 
.A1(n_1366),
.A2(n_1338),
.B1(n_1341),
.B2(n_1339),
.C1(n_1343),
.C2(n_1345),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1352),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1366),
.A2(n_1367),
.B1(n_1359),
.B2(n_1365),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1398),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1355),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1350),
.B(n_1330),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1367),
.A2(n_1307),
.B1(n_1318),
.B2(n_1326),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1357),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1353),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1355),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1360),
.B(n_1330),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1375),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1409),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1412),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1413),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1361),
.B(n_1341),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_SL g1435 ( 
.A(n_1362),
.B(n_1331),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1407),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1399),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1377),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1380),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1347),
.B(n_1332),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1348),
.B(n_1349),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1369),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1399),
.B(n_1416),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1351),
.B(n_1332),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1406),
.B(n_1342),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1406),
.B(n_1342),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1388),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1396),
.B(n_1314),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1392),
.Y(n_1449)
);

NOR2xp67_ASAP7_75t_L g1450 ( 
.A(n_1381),
.B(n_1336),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1369),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1403),
.B(n_1337),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1403),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1396),
.B(n_1395),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1390),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1415),
.B(n_1334),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1409),
.B(n_1291),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1354),
.B(n_1297),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1390),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1376),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1376),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1455),
.B(n_1381),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1432),
.B(n_1370),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1441),
.B(n_1359),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1418),
.B(n_1459),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1432),
.B(n_1372),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1447),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1452),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1436),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1447),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1441),
.B(n_1410),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1445),
.B(n_1410),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1445),
.B(n_1417),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1426),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1418),
.B(n_1460),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1449),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1446),
.B(n_1374),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1426),
.B(n_1379),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1460),
.B(n_1356),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1449),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1421),
.A2(n_1385),
.B(n_1414),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1461),
.B(n_1379),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1422),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1422),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1433),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1454),
.B(n_1374),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1428),
.B(n_1423),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1428),
.B(n_1383),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1442),
.B(n_1401),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1454),
.B(n_1458),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1451),
.B(n_1386),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1432),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1461),
.B(n_1383),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1453),
.B(n_1358),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1483),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1475),
.B(n_1424),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1492),
.A2(n_1457),
.B(n_1419),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1483),
.Y(n_1498)
);

NAND2x2_ASAP7_75t_L g1499 ( 
.A(n_1465),
.B(n_1429),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1469),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1490),
.B(n_1434),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1490),
.B(n_1420),
.Y(n_1502)
);

OAI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1464),
.A2(n_1400),
.B(n_1458),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1463),
.B(n_1440),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1484),
.Y(n_1505)
);

INVxp67_ASAP7_75t_SL g1506 ( 
.A(n_1487),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1487),
.B(n_1437),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1485),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1467),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1463),
.B(n_1444),
.Y(n_1510)
);

NAND2x1p5_ASAP7_75t_L g1511 ( 
.A(n_1488),
.B(n_1431),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1471),
.B(n_1437),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1474),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1492),
.A2(n_1385),
.B(n_1448),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1481),
.A2(n_1450),
.B(n_1373),
.Y(n_1515)
);

NOR3x1_ASAP7_75t_L g1516 ( 
.A(n_1494),
.B(n_1474),
.C(n_1479),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1464),
.B(n_1427),
.Y(n_1517)
);

AOI32xp33_ASAP7_75t_L g1518 ( 
.A1(n_1503),
.A2(n_1486),
.A3(n_1477),
.B1(n_1506),
.B2(n_1472),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1495),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1496),
.B(n_1386),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1504),
.B(n_1471),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1498),
.Y(n_1522)
);

OAI33xp33_ASAP7_75t_L g1523 ( 
.A1(n_1517),
.A2(n_1482),
.A3(n_1493),
.B1(n_1488),
.B2(n_1478),
.B3(n_1480),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1501),
.B(n_1506),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1505),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1508),
.B(n_1470),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1509),
.B(n_1476),
.Y(n_1527)
);

NOR2x1_ASAP7_75t_L g1528 ( 
.A(n_1507),
.B(n_1491),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1502),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1512),
.Y(n_1530)
);

OAI322xp33_ASAP7_75t_L g1531 ( 
.A1(n_1514),
.A2(n_1497),
.A3(n_1478),
.B1(n_1489),
.B2(n_1430),
.C1(n_1439),
.C2(n_1438),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1515),
.A2(n_1486),
.B1(n_1477),
.B2(n_1443),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1500),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1533),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1519),
.Y(n_1535)
);

NOR3xp33_ASAP7_75t_L g1536 ( 
.A(n_1531),
.B(n_1462),
.C(n_1497),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1522),
.Y(n_1537)
);

AO22x1_ASAP7_75t_L g1538 ( 
.A1(n_1528),
.A2(n_1516),
.B1(n_1510),
.B2(n_1466),
.Y(n_1538)
);

OAI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1532),
.A2(n_1499),
.B1(n_1514),
.B2(n_1378),
.C(n_1425),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1523),
.A2(n_1499),
.B1(n_1444),
.B2(n_1473),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1526),
.Y(n_1541)
);

OAI21xp33_ASAP7_75t_L g1542 ( 
.A1(n_1536),
.A2(n_1518),
.B(n_1524),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1541),
.B(n_1529),
.Y(n_1543)
);

OAI211xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1535),
.A2(n_1520),
.B(n_1526),
.C(n_1527),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1539),
.A2(n_1527),
.B(n_1525),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1537),
.A2(n_1513),
.B(n_1530),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1542),
.B(n_1540),
.Y(n_1547)
);

O2A1O1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1545),
.A2(n_1544),
.B(n_1539),
.C(n_1546),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1543),
.A2(n_1538),
.B(n_1513),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1542),
.B(n_1521),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1542),
.A2(n_1382),
.B1(n_1534),
.B2(n_1364),
.Y(n_1551)
);

NAND4xp25_ASAP7_75t_L g1552 ( 
.A(n_1542),
.B(n_1404),
.C(n_1393),
.D(n_1468),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1548),
.B(n_1549),
.Y(n_1553)
);

NOR3xp33_ASAP7_75t_L g1554 ( 
.A(n_1547),
.B(n_1394),
.C(n_1389),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1550),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1555),
.Y(n_1556)
);

NOR3xp33_ASAP7_75t_L g1557 ( 
.A(n_1553),
.B(n_1552),
.C(n_1551),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1556),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1558),
.Y(n_1559)
);

NOR3xp33_ASAP7_75t_L g1560 ( 
.A(n_1559),
.B(n_1557),
.C(n_1554),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1560),
.A2(n_1404),
.B(n_1397),
.Y(n_1561)
);

AOI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1561),
.A2(n_1402),
.B1(n_1411),
.B2(n_1384),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1562),
.A2(n_1402),
.B1(n_1511),
.B2(n_1391),
.Y(n_1563)
);

XNOR2xp5_ASAP7_75t_L g1564 ( 
.A(n_1563),
.B(n_1387),
.Y(n_1564)
);

AOI21xp33_ASAP7_75t_SL g1565 ( 
.A1(n_1564),
.A2(n_1408),
.B(n_1368),
.Y(n_1565)
);

XNOR2xp5_ASAP7_75t_L g1566 ( 
.A(n_1565),
.B(n_1371),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1566),
.A2(n_1435),
.B1(n_1405),
.B2(n_1456),
.Y(n_1567)
);


endmodule