module fake_jpeg_28870_n_122 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_122);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_33),
.Y(n_55)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_41),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.C(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_35),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_13),
.B1(n_24),
.B2(n_26),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_52),
.B1(n_57),
.B2(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_18),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_27),
.C(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_27),
.A2(n_15),
.B1(n_22),
.B2(n_17),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_16),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_31),
.B1(n_40),
.B2(n_35),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_67),
.B1(n_54),
.B2(n_55),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_45),
.B1(n_58),
.B2(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_35),
.C(n_36),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_9),
.Y(n_74)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_55),
.A3(n_10),
.B1(n_4),
.B2(n_6),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_56),
.B1(n_58),
.B2(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_60),
.B1(n_73),
.B2(n_67),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_79),
.A2(n_66),
.B1(n_63),
.B2(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_85),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_67),
.B1(n_61),
.B2(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_93),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_79),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_79),
.B1(n_80),
.B2(n_84),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

OAI322xp33_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_95),
.A3(n_75),
.B1(n_87),
.B2(n_82),
.C1(n_89),
.C2(n_79),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_107),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_93),
.B(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_76),
.B1(n_85),
.B2(n_78),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_102),
.C(n_96),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_112),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_99),
.C(n_76),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_105),
.B1(n_98),
.B2(n_106),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_7),
.C(n_11),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_3),
.B(n_117),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_115),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_115),
.Y(n_122)
);


endmodule