module fake_netlist_6_4698_n_4591 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_443, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4591);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4591;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_700;
wire n_3783;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_4504;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_783;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4285;
wire n_4134;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_1009;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_4578;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_461;
wire n_1371;
wire n_1285;
wire n_873;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_4213;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_4531;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_2247;
wire n_544;
wire n_1711;
wire n_1078;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_522;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_4555;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_4308;
wire n_658;
wire n_616;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3737;
wire n_3624;
wire n_3077;
wire n_3979;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_4563;
wire n_493;
wire n_3107;
wire n_4556;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_4142;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4255;
wire n_4403;
wire n_4071;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_4549;
wire n_4575;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_1986;
wire n_699;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_813;
wire n_2080;
wire n_1909;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_3910;
wire n_1699;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_4507;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4581;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4377;
wire n_4158;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_4544;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_966;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_764;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4337;
wire n_4161;
wire n_4130;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_882;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_4526;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1950;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1664;
wire n_1722;
wire n_612;
wire n_4585;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2749;
wire n_2008;
wire n_3346;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_2254;
wire n_3298;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_4427;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4386;
wire n_4485;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_4523;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_816;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_2994;
wire n_1750;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_4552;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_825;
wire n_728;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_4510;
wire n_696;
wire n_1515;
wire n_4473;
wire n_961;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_4589;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_4560;
wire n_590;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1033;
wire n_462;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_595;
wire n_627;
wire n_1767;
wire n_3253;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3337;
wire n_3450;
wire n_3431;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_4588;
wire n_585;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3614;
wire n_840;
wire n_2913;
wire n_3421;
wire n_874;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_2535;
wire n_1880;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_4576;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_4389;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4540;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4240;
wire n_3491;
wire n_4156;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3353;
wire n_3150;
wire n_3018;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_765;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_4058;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3348;
wire n_3229;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_4481;
wire n_1246;
wire n_4528;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4587;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_4525;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4541;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4551;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_777;
wire n_4459;
wire n_1299;
wire n_4545;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3325;
wire n_3203;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_458;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_4455;
wire n_4453;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_4514;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4564;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_2424;
wire n_1604;
wire n_1284;
wire n_2296;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_4487;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1774;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_2354;
wire n_2682;
wire n_1475;
wire n_3103;
wire n_3032;
wire n_3638;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_3393;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_2442;
wire n_3627;
wire n_3451;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_1418;
wire n_1250;
wire n_958;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3641;
wire n_767;
wire n_3591;
wire n_1837;
wire n_600;
wire n_964;
wire n_831;
wire n_1314;
wire n_2788;
wire n_2218;
wire n_4533;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3909;
wire n_3944;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2357;
wire n_2025;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_4584;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_4430;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_4428;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4204;
wire n_4261;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_4570;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4056;
wire n_1617;
wire n_4034;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_4355;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_3016;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3688;
wire n_3566;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_1129;
wire n_3870;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_4470;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_4546;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_4583;
wire n_465;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4252;
wire n_4357;
wire n_4067;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4509;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_4374;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3276;
wire n_1934;
wire n_3250;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_4582;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_4420;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_4574;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_4405;
wire n_610;
wire n_4304;
wire n_4413;
wire n_4234;
wire n_1403;
wire n_1669;
wire n_4558;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_468;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_466;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_1818;
wire n_1108;
wire n_710;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_3042;
wire n_1356;
wire n_1589;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_3249;
wire n_1320;
wire n_2716;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_4590;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4192;
wire n_4109;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4038;
wire n_2790;
wire n_4131;
wire n_4565;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_4567;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_4554;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_4586;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2373;
wire n_1472;
wire n_2050;
wire n_2120;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_662;
wire n_3501;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_4515;
wire n_3845;
wire n_2017;
wire n_1682;
wire n_4516;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_4547;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_2760;
wire n_1979;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_4548;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_456;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_4553;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_482;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_4209;
wire n_4279;
wire n_2871;
wire n_4135;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_4561;
wire n_804;
wire n_4461;
wire n_464;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4571;
wire n_4343;
wire n_2835;
wire n_4530;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_3074;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_652;
wire n_2154;
wire n_2727;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3932;
wire n_3762;
wire n_3469;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_4524;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_4469;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_4572;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_4493;
wire n_2695;
wire n_4269;
wire n_3818;
wire n_4035;
wire n_743;
wire n_766;
wire n_3124;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_2888;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_4539;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_4421;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_1742;
wire n_3190;
wire n_4505;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_4542;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_4462;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_4536;
wire n_4543;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4173;
wire n_2752;
wire n_4324;
wire n_3135;
wire n_4157;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_4550;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_4534;
wire n_3846;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_4408;
wire n_4577;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_4439;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_3231;
wire n_4083;
wire n_4494;
wire n_1554;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_2380;
wire n_769;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_4579;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_2149;
wire n_1754;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_4557;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_4432;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_4568;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_4569;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_4559;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_4373;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2465;
wire n_1112;
wire n_2275;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_4521;
wire n_2444;
wire n_1215;
wire n_839;
wire n_2437;
wire n_2743;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_709;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4313;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_492;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_4532;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_2666;
wire n_4105;
wire n_1851;
wire n_1585;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_4486;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1362;
wire n_1156;
wire n_4259;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_4353;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_4529;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_4537;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4351;
wire n_4346;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_4396;
wire n_1244;
wire n_1685;
wire n_4508;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2478;
wire n_1619;
wire n_2303;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4460;
wire n_1133;
wire n_4108;
wire n_635;
wire n_1194;
wire n_3374;
wire n_4429;
wire n_4506;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_4538;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_553;
wire n_849;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_467;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_4580;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4522;
wire n_4148;
wire n_571;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_2280;
wire n_1888;
wire n_1557;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_640;
wire n_1322;
wire n_4129;
wire n_4457;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_4500;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_457;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_4566;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_4482;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_4426;
wire n_531;
wire n_827;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_4030;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_8),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_225),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_102),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_19),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_196),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_70),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_113),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_348),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_104),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_225),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_183),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_140),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_162),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_419),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_140),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_260),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_109),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_263),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_58),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_146),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_274),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_135),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_182),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_392),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_252),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_222),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_308),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_166),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_150),
.Y(n_486)
);

BUFx5_ASAP7_75t_L g487 ( 
.A(n_378),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_430),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_146),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_191),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_445),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_415),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_407),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_88),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_414),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_199),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_20),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_194),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_449),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_328),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_398),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_432),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_93),
.Y(n_503)
);

BUFx5_ASAP7_75t_L g504 ( 
.A(n_292),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_50),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_61),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_304),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_145),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_388),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_114),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_237),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_135),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_106),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_429),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_224),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_261),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_105),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_380),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_61),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_340),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_169),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_381),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_385),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_374),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_79),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_371),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_370),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_356),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_64),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_300),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_114),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_80),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_173),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_102),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_138),
.Y(n_535)
);

BUFx5_ASAP7_75t_L g536 ( 
.A(n_365),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_310),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_412),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_360),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_279),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_364),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_324),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_69),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_119),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_168),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_81),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_16),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_433),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_20),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_187),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_418),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_159),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_99),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_437),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_32),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_311),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_142),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_184),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_188),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_83),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_332),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_382),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_451),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_131),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_139),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_54),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_202),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_448),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_387),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_367),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_416),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_244),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_272),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_105),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_282),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_27),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_410),
.Y(n_577)
);

BUFx10_ASAP7_75t_L g578 ( 
.A(n_397),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_226),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_10),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_238),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_377),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_127),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_99),
.Y(n_584)
);

CKINVDCx14_ASAP7_75t_R g585 ( 
.A(n_2),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_40),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_349),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_76),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_217),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_231),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_50),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_81),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_368),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_131),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_323),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_257),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_232),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_447),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_243),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_100),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_48),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_446),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_280),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_72),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_4),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_30),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_49),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_286),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_178),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_89),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_157),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_186),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_420),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_106),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_329),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_425),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_394),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_234),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_142),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_90),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_362),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_422),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_17),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_315),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_212),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_267),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_201),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_201),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_423),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_27),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_92),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_137),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_74),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_337),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_53),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_177),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_386),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_316),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_438),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_74),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_14),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_8),
.Y(n_642)
);

CKINVDCx16_ASAP7_75t_R g643 ( 
.A(n_453),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_43),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_357),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_33),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_151),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_247),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_346),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_171),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_455),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_111),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_117),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_22),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_271),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_177),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_314),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_265),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_91),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_393),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_191),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_170),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_440),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_288),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_335),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_334),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_56),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_390),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_79),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_236),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_442),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_65),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_47),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_109),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_167),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_224),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_251),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_352),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_45),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_269),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_120),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_93),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_125),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_284),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_431),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_208),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_150),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_400),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_421),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_233),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_144),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_319),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_1),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_355),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_444),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_69),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_338),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_435),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_426),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_436),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_246),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_270),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_318),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_226),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_294),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_341),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_283),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_199),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_411),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_71),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_22),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_285),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_259),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_373),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_313),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_67),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_103),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_94),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_47),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_452),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_25),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_278),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_53),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_454),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_434),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_117),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_342),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_44),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_443),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_31),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_104),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_428),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_89),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_427),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_194),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_26),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_218),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_375),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_214),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_185),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_186),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_9),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_10),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_148),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_65),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_424),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_170),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_309),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_213),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_71),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_208),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_125),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_254),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_195),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_111),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_145),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_138),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_63),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_159),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_46),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_160),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_82),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_200),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_220),
.Y(n_764)
);

BUFx10_ASAP7_75t_L g765 ( 
.A(n_130),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_376),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_391),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_214),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_158),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_441),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_130),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_221),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_212),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_57),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_450),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_42),
.Y(n_776)
);

BUFx10_ASAP7_75t_L g777 ( 
.A(n_51),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_401),
.Y(n_778)
);

CKINVDCx14_ASAP7_75t_R g779 ( 
.A(n_49),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_121),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_41),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_7),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_6),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_157),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_78),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_175),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_76),
.Y(n_787)
);

CKINVDCx16_ASAP7_75t_R g788 ( 
.A(n_525),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_693),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_514),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_693),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_693),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_456),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_467),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_516),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_606),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_460),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_460),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_468),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_606),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_468),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_782),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_545),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_518),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_523),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_734),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_524),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_545),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_537),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_708),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_480),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_585),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_606),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_779),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_490),
.Y(n_815)
);

CKINVDCx16_ASAP7_75t_R g816 ( 
.A(n_643),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_708),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_733),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_733),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_508),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_752),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_513),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_549),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_510),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_752),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_566),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_512),
.Y(n_827)
);

BUFx10_ASAP7_75t_L g828 ( 
.A(n_640),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_606),
.Y(n_829)
);

BUFx10_ASAP7_75t_L g830 ( 
.A(n_606),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_719),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_567),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_669),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_719),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_719),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_719),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_515),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_593),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_519),
.Y(n_839)
);

BUFx5_ASAP7_75t_L g840 ( 
.A(n_469),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_521),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_593),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_719),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_780),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_780),
.Y(n_845)
);

BUFx5_ASAP7_75t_L g846 ( 
.A(n_477),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_538),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_780),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_735),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_747),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_780),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_541),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_734),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_542),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_457),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_780),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_459),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_487),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_548),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_551),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_561),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_734),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_462),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_563),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_730),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_734),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_568),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_457),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_569),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_487),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_570),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_575),
.Y(n_872)
);

BUFx10_ASAP7_75t_L g873 ( 
.A(n_472),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_465),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_577),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_581),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_582),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_587),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_730),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_466),
.Y(n_880)
);

CKINVDCx14_ASAP7_75t_R g881 ( 
.A(n_530),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_608),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_730),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_624),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_473),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_487),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_626),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_483),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_485),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_634),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_497),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_503),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_487),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_517),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_529),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_637),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_639),
.Y(n_897)
);

CKINVDCx16_ASAP7_75t_R g898 ( 
.A(n_765),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_648),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_458),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_533),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_535),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_651),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_560),
.Y(n_904)
);

CKINVDCx16_ASAP7_75t_R g905 ( 
.A(n_765),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_565),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_660),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_664),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_558),
.B(n_0),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_734),
.Y(n_910)
);

NOR2xp67_ASAP7_75t_L g911 ( 
.A(n_558),
.B(n_0),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_666),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_487),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_670),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_576),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_603),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_579),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_671),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_588),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_678),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_680),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_684),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_765),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_688),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_724),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_592),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_738),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_594),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_609),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_614),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_625),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_777),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_531),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_630),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_635),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_746),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_642),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_487),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_487),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_652),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_653),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_656),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_532),
.Y(n_943)
);

INVxp67_ASAP7_75t_SL g944 ( 
.A(n_540),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_534),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_661),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_766),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_487),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_767),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_672),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_674),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_675),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_598),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_679),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_686),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_691),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_458),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_704),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_716),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_718),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_504),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_663),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_685),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_705),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_602),
.B(n_1),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_726),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_603),
.Y(n_967)
);

CKINVDCx16_ASAP7_75t_R g968 ( 
.A(n_777),
.Y(n_968)
);

CKINVDCx11_ASAP7_75t_R g969 ( 
.A(n_777),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_736),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_707),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_740),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_475),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_742),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_744),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_573),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_750),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_754),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_727),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_543),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_771),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_776),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_786),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_482),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_504),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_484),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_461),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_544),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_505),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_479),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_461),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_464),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_546),
.Y(n_993)
);

INVxp67_ASAP7_75t_SL g994 ( 
.A(n_658),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_488),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_573),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_547),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_550),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_552),
.Y(n_999)
);

BUFx5_ASAP7_75t_L g1000 ( 
.A(n_502),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_504),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_511),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_520),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_479),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_464),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_553),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_522),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_526),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_632),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_527),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_554),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_556),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_555),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_787),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_571),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_572),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_785),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_590),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_595),
.Y(n_1019)
);

NOR2xp67_ASAP7_75t_L g1020 ( 
.A(n_632),
.B(n_2),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_596),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_573),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_599),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_613),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_471),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_557),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_615),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_618),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_621),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_559),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_629),
.Y(n_1031)
);

INVxp33_ASAP7_75t_L g1032 ( 
.A(n_650),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_638),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_785),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_564),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_657),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_665),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_471),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_668),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_476),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_574),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_580),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_476),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_689),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_583),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_690),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_695),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_584),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_586),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_700),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_589),
.Y(n_1051)
);

NOR2xp67_ASAP7_75t_L g1052 ( 
.A(n_650),
.B(n_3),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_701),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_591),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_712),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_725),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_748),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_753),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_770),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_645),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_645),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_600),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_478),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_655),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_655),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_697),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_697),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_706),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_601),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_578),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_604),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_706),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_681),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_478),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_605),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_607),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_681),
.B(n_3),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_743),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_743),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_472),
.Y(n_1080)
);

CKINVDCx14_ASAP7_75t_R g1081 ( 
.A(n_578),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_597),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_610),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_611),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_778),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_597),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_616),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_616),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_486),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_617),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_617),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_612),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_504),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_619),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_504),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_620),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_623),
.Y(n_1097)
);

INVxp67_ASAP7_75t_L g1098 ( 
.A(n_784),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_627),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_628),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_631),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_633),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_649),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_636),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_486),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_504),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_649),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_677),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_504),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_641),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_677),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_578),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_644),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_646),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_647),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_654),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_694),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_659),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_694),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_662),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_667),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_673),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_504),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_676),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_682),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_683),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_489),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_687),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_536),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_536),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_489),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_536),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_737),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_739),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_741),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_463),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_494),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_745),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_749),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_494),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_536),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_751),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_755),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_756),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_757),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_509),
.B(n_4),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_758),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_759),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_760),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_463),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_761),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_973),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_790),
.Y(n_1153)
);

INVxp33_ASAP7_75t_L g1154 ( 
.A(n_1025),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_795),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_829),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_831),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_804),
.Y(n_1158)
);

INVxp33_ASAP7_75t_SL g1159 ( 
.A(n_812),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_989),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_793),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_835),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_836),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_R g1164 ( 
.A(n_953),
.B(n_470),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_793),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_843),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_844),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_845),
.Y(n_1168)
);

INVxp67_ASAP7_75t_SL g1169 ( 
.A(n_916),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_805),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_916),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_807),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_848),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_851),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_856),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_916),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_990),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_990),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1014),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_990),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_990),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1004),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_809),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_794),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1004),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_916),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_806),
.Y(n_1187)
);

CKINVDCx16_ASAP7_75t_R g1188 ( 
.A(n_788),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_962),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_963),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_964),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_847),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_1089),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_967),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_852),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_1081),
.Y(n_1196)
);

HB1xp67_ASAP7_75t_L g1197 ( 
.A(n_980),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_796),
.Y(n_1198)
);

CKINVDCx14_ASAP7_75t_R g1199 ( 
.A(n_1081),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1004),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1004),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_789),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_825),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_881),
.B(n_528),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_791),
.Y(n_1205)
);

INVxp33_ASAP7_75t_SL g1206 ( 
.A(n_812),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_796),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_854),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_792),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_988),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_967),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_794),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_993),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_859),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_815),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_967),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_815),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_967),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_800),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_800),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_860),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_822),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_861),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_813),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_813),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_864),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_867),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_830),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_869),
.Y(n_1229)
);

INVxp33_ASAP7_75t_SL g1230 ( 
.A(n_814),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_834),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_834),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_871),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_830),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_971),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_830),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_984),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_986),
.Y(n_1238)
);

NOR2xp67_ASAP7_75t_L g1239 ( 
.A(n_1017),
.B(n_470),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_838),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_995),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1002),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1003),
.Y(n_1243)
);

INVxp67_ASAP7_75t_L g1244 ( 
.A(n_883),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1007),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_872),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_806),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_806),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_875),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_876),
.Y(n_1250)
);

INVxp33_ASAP7_75t_SL g1251 ( 
.A(n_814),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_877),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_878),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_882),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_822),
.Y(n_1255)
);

XNOR2x1_ASAP7_75t_L g1256 ( 
.A(n_811),
.B(n_496),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_884),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1008),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1010),
.Y(n_1259)
);

NOR2xp67_ASAP7_75t_L g1260 ( 
.A(n_1034),
.B(n_474),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1011),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_881),
.B(n_539),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1012),
.Y(n_1263)
);

CKINVDCx5p33_ASAP7_75t_R g1264 ( 
.A(n_887),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_890),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_823),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_806),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_997),
.Y(n_1268)
);

INVxp33_ASAP7_75t_L g1269 ( 
.A(n_1120),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1035),
.B(n_1076),
.Y(n_1270)
);

NOR2xp67_ASAP7_75t_L g1271 ( 
.A(n_1098),
.B(n_474),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_823),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_896),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1015),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_853),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1016),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1018),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_832),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1019),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_897),
.Y(n_1280)
);

CKINVDCx20_ASAP7_75t_R g1281 ( 
.A(n_832),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1084),
.B(n_562),
.Y(n_1282)
);

BUFx2_ASAP7_75t_SL g1283 ( 
.A(n_855),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_833),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_899),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1021),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1104),
.B(n_692),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_833),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_838),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_903),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_907),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_908),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_849),
.Y(n_1293)
);

NOR2xp67_ASAP7_75t_L g1294 ( 
.A(n_912),
.B(n_481),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1023),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_849),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_998),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1024),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1027),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_914),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_853),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1136),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_918),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1028),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1029),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_850),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_976),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1031),
.Y(n_1308)
);

INVxp33_ASAP7_75t_SL g1309 ( 
.A(n_965),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_976),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1033),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1036),
.Y(n_1312)
);

BUFx3_ASAP7_75t_L g1313 ( 
.A(n_842),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_850),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_920),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1037),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_921),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_969),
.Y(n_1318)
);

CKINVDCx20_ASAP7_75t_R g1319 ( 
.A(n_969),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1039),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_922),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1044),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_853),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_855),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1136),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1046),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1047),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_924),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1050),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1053),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1055),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1056),
.Y(n_1332)
);

INVxp33_ASAP7_75t_SL g1333 ( 
.A(n_925),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1057),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1138),
.B(n_722),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1058),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_999),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_927),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1059),
.Y(n_1339)
);

INVxp33_ASAP7_75t_SL g1340 ( 
.A(n_936),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1006),
.Y(n_1341)
);

INVxp67_ASAP7_75t_SL g1342 ( 
.A(n_1150),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_996),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_947),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_857),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_868),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_853),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_863),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_874),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_949),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_979),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1013),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1026),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_802),
.B(n_762),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_868),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1030),
.B(n_481),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_880),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1041),
.Y(n_1358)
);

INVxp67_ASAP7_75t_SL g1359 ( 
.A(n_1150),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_885),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_888),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_889),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_891),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_996),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_892),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1042),
.B(n_491),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_894),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_895),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_900),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_900),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_862),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_901),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_957),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_902),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_904),
.Y(n_1375)
);

CKINVDCx16_ASAP7_75t_R g1376 ( 
.A(n_1112),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1045),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_906),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_915),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_862),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_842),
.B(n_763),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_862),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_957),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_898),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_987),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_862),
.Y(n_1386)
);

CKINVDCx16_ASAP7_75t_R g1387 ( 
.A(n_905),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_917),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_919),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_816),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_926),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1048),
.Y(n_1392)
);

INVxp67_ASAP7_75t_SL g1393 ( 
.A(n_1122),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1049),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_928),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_929),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_930),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_987),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_991),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1051),
.B(n_491),
.Y(n_1400)
);

BUFx2_ASAP7_75t_L g1401 ( 
.A(n_991),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1022),
.Y(n_1402)
);

CKINVDCx16_ASAP7_75t_R g1403 ( 
.A(n_968),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1080),
.B(n_492),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1054),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1062),
.B(n_492),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1115),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_992),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1116),
.Y(n_1409)
);

BUFx2_ASAP7_75t_SL g1410 ( 
.A(n_992),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1118),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1121),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1125),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_931),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_934),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_935),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1005),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1126),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1005),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1134),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1142),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1038),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1038),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_937),
.Y(n_1424)
);

INVxp33_ASAP7_75t_L g1425 ( 
.A(n_1124),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_940),
.Y(n_1426)
);

INVxp67_ASAP7_75t_SL g1427 ( 
.A(n_1128),
.Y(n_1427)
);

CKINVDCx20_ASAP7_75t_R g1428 ( 
.A(n_1040),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1144),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_866),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1147),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_941),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1040),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_820),
.Y(n_1434)
);

INVxp33_ASAP7_75t_L g1435 ( 
.A(n_1133),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_942),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_1043),
.Y(n_1437)
);

INVxp67_ASAP7_75t_L g1438 ( 
.A(n_1022),
.Y(n_1438)
);

NOR2xp67_ASAP7_75t_L g1439 ( 
.A(n_820),
.B(n_493),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_824),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1043),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_824),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1063),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_946),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1063),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_827),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_827),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_950),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_866),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_951),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_837),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_837),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_839),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_839),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_841),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_952),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1074),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1198),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1282),
.B(n_1085),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1179),
.Y(n_1460)
);

BUFx8_ASAP7_75t_L g1461 ( 
.A(n_1401),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1345),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1348),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1198),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1349),
.Y(n_1465)
);

OAI22x1_ASAP7_75t_R g1466 ( 
.A1(n_1318),
.A2(n_1105),
.B1(n_1127),
.B2(n_1074),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1207),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1269),
.B(n_841),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1323),
.Y(n_1469)
);

BUFx8_ASAP7_75t_L g1470 ( 
.A(n_1441),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1207),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1287),
.B(n_1335),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1323),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1231),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1323),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1231),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1169),
.B(n_840),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1323),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1270),
.B(n_944),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1171),
.B(n_840),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1357),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1194),
.Y(n_1482)
);

OAI22x1_ASAP7_75t_R g1483 ( 
.A1(n_1318),
.A2(n_1127),
.B1(n_1131),
.B2(n_1105),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1360),
.Y(n_1484)
);

NOR2x1_ASAP7_75t_L g1485 ( 
.A(n_1228),
.B(n_1070),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1219),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1194),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1187),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1177),
.A2(n_1061),
.B(n_1060),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1187),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1361),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1362),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1161),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1152),
.B(n_826),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1220),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1363),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1224),
.Y(n_1497)
);

CKINVDCx11_ASAP7_75t_R g1498 ( 
.A(n_1319),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1160),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1225),
.Y(n_1500)
);

AND2x6_ASAP7_75t_L g1501 ( 
.A(n_1404),
.B(n_1135),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1365),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1178),
.A2(n_1065),
.B(n_1064),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1309),
.B(n_933),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1202),
.B(n_1151),
.Y(n_1505)
);

CKINVDCx16_ASAP7_75t_R g1506 ( 
.A(n_1188),
.Y(n_1506)
);

AND2x2_ASAP7_75t_SL g1507 ( 
.A(n_1204),
.B(n_1146),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1367),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1164),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1232),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1368),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1187),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1309),
.A2(n_994),
.B1(n_943),
.B2(n_945),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1248),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1372),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1374),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1161),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1375),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1240),
.B(n_1082),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1378),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1240),
.B(n_1289),
.Y(n_1521)
);

CKINVDCx6p67_ASAP7_75t_R g1522 ( 
.A(n_1196),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1351),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1247),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1248),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1244),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1267),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1289),
.B(n_1086),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1379),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1267),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1256),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1388),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1247),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1389),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1203),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1247),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1275),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1313),
.B(n_1087),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1205),
.B(n_1149),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1176),
.B(n_840),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1186),
.B(n_840),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1425),
.B(n_933),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1313),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1391),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1395),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1239),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1275),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1262),
.A2(n_945),
.B1(n_1069),
.B2(n_943),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1393),
.B(n_840),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1234),
.A2(n_870),
.B(n_858),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1386),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1301),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1396),
.Y(n_1553)
);

INVx5_ASAP7_75t_L g1554 ( 
.A(n_1386),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1397),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1435),
.B(n_1069),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1386),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1449),
.Y(n_1558)
);

AND2x2_ASAP7_75t_SL g1559 ( 
.A(n_1356),
.B(n_1077),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1427),
.B(n_1071),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1414),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1449),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1165),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1301),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1415),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1416),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1193),
.A2(n_1071),
.B1(n_1083),
.B2(n_1075),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1347),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1347),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1371),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1424),
.Y(n_1571)
);

INVx3_ASAP7_75t_L g1572 ( 
.A(n_1449),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1371),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1302),
.B(n_1325),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1380),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1211),
.B(n_1088),
.Y(n_1576)
);

NAND2xp33_ASAP7_75t_L g1577 ( 
.A(n_1381),
.B(n_536),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1342),
.B(n_1075),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1380),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1426),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1359),
.B(n_840),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1432),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1382),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1382),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1430),
.Y(n_1585)
);

AND2x6_ASAP7_75t_L g1586 ( 
.A(n_1404),
.B(n_1139),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1209),
.B(n_1148),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1216),
.B(n_840),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1436),
.Y(n_1589)
);

BUFx12f_ASAP7_75t_L g1590 ( 
.A(n_1390),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1430),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1218),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_L g1593 ( 
.A(n_1237),
.B(n_536),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1156),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1199),
.B(n_1083),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1404),
.Y(n_1596)
);

INVx6_ASAP7_75t_L g1597 ( 
.A(n_1228),
.Y(n_1597)
);

OA21x2_ASAP7_75t_L g1598 ( 
.A1(n_1180),
.A2(n_1067),
.B(n_1066),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1366),
.B(n_1092),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1157),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1189),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1181),
.Y(n_1602)
);

INVx4_ASAP7_75t_L g1603 ( 
.A(n_1182),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1444),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1448),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1450),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1456),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1189),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1190),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1238),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1241),
.B(n_1090),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1354),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1185),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1307),
.B(n_1092),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1242),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1162),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1163),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1243),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1245),
.B(n_1143),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1166),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1258),
.Y(n_1621)
);

BUFx6f_ASAP7_75t_L g1622 ( 
.A(n_1200),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1259),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1167),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1261),
.B(n_1091),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1201),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1168),
.Y(n_1627)
);

OA21x2_ASAP7_75t_L g1628 ( 
.A1(n_1173),
.A2(n_1072),
.B(n_1068),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1174),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1263),
.B(n_1145),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1175),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1274),
.Y(n_1632)
);

AND2x2_ASAP7_75t_SL g1633 ( 
.A(n_1400),
.B(n_1103),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1236),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1276),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1277),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1279),
.B(n_1107),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1439),
.B(n_1094),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1256),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1286),
.B(n_1108),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1295),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1298),
.Y(n_1642)
);

INVx5_ASAP7_75t_L g1643 ( 
.A(n_1376),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1299),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1304),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1305),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1308),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1311),
.B(n_1111),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1294),
.B(n_846),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1312),
.B(n_1032),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1316),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1406),
.A2(n_1094),
.B1(n_1097),
.B2(n_1096),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1310),
.B(n_1096),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1320),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1260),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1322),
.B(n_1117),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1271),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1326),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1190),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1327),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1329),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1343),
.B(n_846),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1330),
.A2(n_870),
.B(n_858),
.Y(n_1663)
);

INVx4_ASAP7_75t_L g1664 ( 
.A(n_1153),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1331),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1333),
.A2(n_1099),
.B1(n_1100),
.B2(n_1097),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1191),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1332),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1333),
.A2(n_1100),
.B1(n_1101),
.B2(n_1099),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1334),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1336),
.B(n_1119),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1339),
.B(n_1032),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1364),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1402),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1438),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1324),
.A2(n_1137),
.B1(n_1140),
.B2(n_1131),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1197),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1210),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1213),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1353),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1155),
.B(n_846),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1268),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1297),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1337),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1341),
.Y(n_1685)
);

AND2x6_ASAP7_75t_L g1686 ( 
.A(n_1340),
.B(n_886),
.Y(n_1686)
);

CKINVDCx6p67_ASAP7_75t_R g1687 ( 
.A(n_1319),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1158),
.B(n_846),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1352),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1170),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1154),
.B(n_797),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1172),
.Y(n_1692)
);

OAI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1394),
.A2(n_893),
.B(n_886),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1411),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1183),
.B(n_954),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1340),
.A2(n_1101),
.B1(n_1110),
.B2(n_1102),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1192),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1195),
.B(n_846),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1208),
.B(n_798),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1214),
.B(n_799),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1191),
.Y(n_1701)
);

NAND2xp33_ASAP7_75t_L g1702 ( 
.A(n_1358),
.B(n_536),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1377),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1221),
.A2(n_1110),
.B1(n_1113),
.B2(n_1102),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1223),
.A2(n_1113),
.B1(n_1114),
.B2(n_1137),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1226),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1227),
.B(n_846),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1229),
.Y(n_1708)
);

OAI22x1_ASAP7_75t_R g1709 ( 
.A1(n_1165),
.A2(n_1140),
.B1(n_498),
.B2(n_506),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1407),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1233),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1246),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1249),
.B(n_955),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1250),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1434),
.Y(n_1715)
);

INVx1_ASAP7_75t_SL g1716 ( 
.A(n_1283),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1252),
.Y(n_1717)
);

BUFx6f_ASAP7_75t_L g1718 ( 
.A(n_1253),
.Y(n_1718)
);

OA21x2_ASAP7_75t_L g1719 ( 
.A1(n_1254),
.A2(n_913),
.B(n_893),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1257),
.A2(n_1114),
.B1(n_1070),
.B2(n_879),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1264),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1265),
.B(n_956),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1440),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1273),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1280),
.B(n_846),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1285),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1290),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1235),
.Y(n_1728)
);

OA21x2_ASAP7_75t_L g1729 ( 
.A1(n_1291),
.A2(n_938),
.B(n_913),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1292),
.B(n_1000),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1300),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1303),
.B(n_1000),
.Y(n_1732)
);

OA21x2_ASAP7_75t_L g1733 ( 
.A1(n_1315),
.A2(n_939),
.B(n_938),
.Y(n_1733)
);

OA21x2_ASAP7_75t_L g1734 ( 
.A1(n_1317),
.A2(n_948),
.B(n_939),
.Y(n_1734)
);

BUFx6f_ASAP7_75t_L g1735 ( 
.A(n_1321),
.Y(n_1735)
);

NOR2x1_ASAP7_75t_L g1736 ( 
.A(n_1410),
.B(n_801),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1328),
.Y(n_1737)
);

INVx6_ASAP7_75t_L g1738 ( 
.A(n_1384),
.Y(n_1738)
);

AND2x6_ASAP7_75t_L g1739 ( 
.A(n_1159),
.B(n_948),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1235),
.Y(n_1740)
);

OA21x2_ASAP7_75t_L g1741 ( 
.A1(n_1338),
.A2(n_985),
.B(n_961),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1344),
.B(n_803),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1350),
.A2(n_1412),
.B1(n_1413),
.B2(n_1409),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1418),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1420),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1421),
.B(n_958),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1429),
.B(n_1000),
.Y(n_1747)
);

INVx6_ASAP7_75t_L g1748 ( 
.A(n_1643),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1663),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1550),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1482),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1472),
.B(n_1392),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1576),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1576),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1663),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1576),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1636),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1636),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1458),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1642),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1642),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1654),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1458),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1499),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1460),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1464),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1654),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1459),
.B(n_1431),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1573),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1550),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1559),
.B(n_1392),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1660),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1660),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1644),
.B(n_1000),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1479),
.B(n_1405),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1464),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1521),
.B(n_959),
.Y(n_1777)
);

NAND2x1p5_ASAP7_75t_L g1778 ( 
.A(n_1596),
.B(n_866),
.Y(n_1778)
);

NAND2x1_ASAP7_75t_L g1779 ( 
.A(n_1686),
.B(n_1533),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1661),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1661),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1670),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1559),
.B(n_1574),
.Y(n_1783)
);

BUFx2_ASAP7_75t_L g1784 ( 
.A(n_1460),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1482),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1670),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1462),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1650),
.B(n_1405),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1467),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1463),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_L g1791 ( 
.A1(n_1693),
.A2(n_985),
.B(n_961),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1465),
.Y(n_1792)
);

OAI21x1_ASAP7_75t_L g1793 ( 
.A1(n_1693),
.A2(n_1093),
.B(n_1001),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1481),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1484),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1491),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1492),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1494),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1467),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1633),
.B(n_1442),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1496),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1502),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1508),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1521),
.B(n_960),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1471),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1596),
.B(n_1446),
.Y(n_1806)
);

NAND2xp33_ASAP7_75t_SL g1807 ( 
.A(n_1612),
.B(n_1447),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1471),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1650),
.B(n_1451),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1526),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1511),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1644),
.B(n_1000),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1474),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1493),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1515),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1581),
.B(n_1452),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1516),
.Y(n_1817)
);

AND3x1_ASAP7_75t_L g1818 ( 
.A(n_1513),
.B(n_1705),
.C(n_1567),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1518),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1474),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1476),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1644),
.B(n_1000),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1520),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1476),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1573),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1482),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1493),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1549),
.B(n_1453),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1529),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1482),
.Y(n_1830)
);

BUFx3_ASAP7_75t_L g1831 ( 
.A(n_1521),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1633),
.B(n_1454),
.Y(n_1832)
);

BUFx8_ASAP7_75t_L g1833 ( 
.A(n_1590),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1489),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1532),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1646),
.B(n_1000),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1489),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1534),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_L g1839 ( 
.A1(n_1533),
.A2(n_1093),
.B(n_1001),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1573),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1544),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1487),
.Y(n_1842)
);

CKINVDCx8_ASAP7_75t_R g1843 ( 
.A(n_1506),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1560),
.B(n_1578),
.C(n_1653),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1545),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1517),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1553),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1646),
.B(n_1681),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1599),
.B(n_1455),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1555),
.Y(n_1850)
);

INVxp67_ASAP7_75t_L g1851 ( 
.A(n_1672),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1561),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1646),
.B(n_873),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1565),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1543),
.B(n_966),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1566),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1571),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1543),
.B(n_970),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1597),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1688),
.B(n_873),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1489),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1503),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1698),
.B(n_873),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1573),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1691),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1707),
.B(n_1159),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1517),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1580),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1582),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1503),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1589),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1604),
.Y(n_1872)
);

AND2x4_ASAP7_75t_L g1873 ( 
.A(n_1665),
.B(n_972),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1503),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1598),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1507),
.B(n_1206),
.Y(n_1876)
);

BUFx8_ASAP7_75t_L g1877 ( 
.A(n_1590),
.Y(n_1877)
);

BUFx2_ASAP7_75t_L g1878 ( 
.A(n_1563),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1598),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1628),
.Y(n_1880)
);

OA21x2_ASAP7_75t_L g1881 ( 
.A1(n_1588),
.A2(n_1106),
.B(n_1095),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1605),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1725),
.B(n_1206),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1606),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1598),
.Y(n_1885)
);

OA21x2_ASAP7_75t_L g1886 ( 
.A1(n_1477),
.A2(n_1106),
.B(n_1095),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1607),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1610),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1730),
.B(n_1230),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1615),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1618),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1628),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1621),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1623),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1628),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1732),
.B(n_1230),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1635),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1641),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1563),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1486),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1647),
.Y(n_1901)
);

BUFx6f_ASAP7_75t_L g1902 ( 
.A(n_1487),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1486),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1672),
.B(n_1387),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1495),
.Y(n_1905)
);

OA21x2_ASAP7_75t_L g1906 ( 
.A1(n_1480),
.A2(n_1123),
.B(n_1109),
.Y(n_1906)
);

OAI22xp33_ASAP7_75t_SL g1907 ( 
.A1(n_1504),
.A2(n_923),
.B1(n_932),
.B2(n_865),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1747),
.B(n_1251),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1651),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1507),
.B(n_1251),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1495),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1658),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1668),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1611),
.Y(n_1914)
);

INVx3_ASAP7_75t_L g1915 ( 
.A(n_1514),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1627),
.B(n_493),
.Y(n_1916)
);

BUFx6f_ASAP7_75t_L g1917 ( 
.A(n_1487),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1497),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1487),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1611),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1468),
.B(n_1403),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1514),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1611),
.Y(n_1923)
);

BUFx6f_ASAP7_75t_L g1924 ( 
.A(n_1632),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1625),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1625),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1625),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1665),
.B(n_974),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1637),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1637),
.Y(n_1930)
);

NAND3xp33_ASAP7_75t_L g1931 ( 
.A(n_1560),
.B(n_810),
.C(n_808),
.Y(n_1931)
);

AND2x6_ASAP7_75t_L g1932 ( 
.A(n_1619),
.B(n_1109),
.Y(n_1932)
);

INVx1_ASAP7_75t_SL g1933 ( 
.A(n_1691),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1497),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1632),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1627),
.B(n_495),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1637),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1468),
.B(n_828),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1640),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1640),
.Y(n_1940)
);

NAND3xp33_ASAP7_75t_L g1941 ( 
.A(n_1578),
.B(n_1653),
.C(n_1599),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1612),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1640),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1542),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1535),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1648),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1648),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1500),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1500),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1510),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1510),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1648),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1525),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1656),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1656),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1699),
.Y(n_1956)
);

INVxp67_ASAP7_75t_L g1957 ( 
.A(n_1542),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1656),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1632),
.B(n_536),
.Y(n_1959)
);

INVxp67_ASAP7_75t_L g1960 ( 
.A(n_1556),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1556),
.B(n_828),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1671),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1671),
.Y(n_1963)
);

HB1xp67_ASAP7_75t_L g1964 ( 
.A(n_1673),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1525),
.Y(n_1965)
);

INVx4_ASAP7_75t_L g1966 ( 
.A(n_1488),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1671),
.Y(n_1967)
);

INVxp67_ASAP7_75t_L g1968 ( 
.A(n_1614),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1594),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1627),
.B(n_495),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1594),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1527),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1662),
.B(n_499),
.Y(n_1973)
);

BUFx2_ASAP7_75t_L g1974 ( 
.A(n_1699),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1600),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1600),
.Y(n_1976)
);

BUFx3_ASAP7_75t_L g1977 ( 
.A(n_1597),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1616),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1527),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1616),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1617),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1632),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_L g1983 ( 
.A(n_1645),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1645),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1530),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1530),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1617),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1739),
.A2(n_1390),
.B1(n_500),
.B2(n_501),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1645),
.B(n_499),
.Y(n_1989)
);

AND2x2_ASAP7_75t_SL g1990 ( 
.A(n_1577),
.B(n_1702),
.Y(n_1990)
);

INVxp67_ASAP7_75t_L g1991 ( 
.A(n_1505),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1537),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1501),
.B(n_500),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1537),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1620),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1547),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1501),
.B(n_501),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1689),
.B(n_828),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1645),
.B(n_507),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1547),
.Y(n_2000)
);

OA21x2_ASAP7_75t_L g2001 ( 
.A1(n_1540),
.A2(n_1129),
.B(n_1123),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1620),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1689),
.B(n_817),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1501),
.B(n_507),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1624),
.Y(n_2005)
);

INVx6_ASAP7_75t_L g2006 ( 
.A(n_1643),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1552),
.Y(n_2007)
);

OA21x2_ASAP7_75t_L g2008 ( 
.A1(n_1541),
.A2(n_1130),
.B(n_1129),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1519),
.B(n_975),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1519),
.B(n_977),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1552),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1624),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1629),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1473),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1473),
.Y(n_2015)
);

BUFx6f_ASAP7_75t_L g2016 ( 
.A(n_1473),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1629),
.Y(n_2017)
);

AND2x6_ASAP7_75t_L g2018 ( 
.A(n_1619),
.B(n_1130),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1631),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1631),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1673),
.B(n_818),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1564),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1675),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1519),
.B(n_978),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1473),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1564),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1528),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1478),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1528),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_1568),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1528),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1538),
.Y(n_2032)
);

INVx3_ASAP7_75t_L g2033 ( 
.A(n_1568),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1538),
.Y(n_2034)
);

AND2x6_ASAP7_75t_L g2035 ( 
.A(n_1630),
.B(n_1132),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1675),
.B(n_622),
.Y(n_2036)
);

HB1xp67_ASAP7_75t_L g2037 ( 
.A(n_1630),
.Y(n_2037)
);

INVx3_ASAP7_75t_L g2038 ( 
.A(n_1569),
.Y(n_2038)
);

BUFx6f_ASAP7_75t_L g2039 ( 
.A(n_1478),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1538),
.Y(n_2040)
);

BUFx8_ASAP7_75t_L g2041 ( 
.A(n_1659),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1569),
.Y(n_2042)
);

BUFx6f_ASAP7_75t_L g2043 ( 
.A(n_1478),
.Y(n_2043)
);

HB1xp67_ASAP7_75t_L g2044 ( 
.A(n_1505),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_SL g2045 ( 
.A1(n_1676),
.A2(n_1346),
.B1(n_1355),
.B2(n_1324),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1570),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1570),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1990),
.B(n_1690),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1759),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1759),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1763),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1933),
.B(n_1700),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1865),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1990),
.A2(n_1577),
.B1(n_1729),
.B2(n_1719),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1900),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1900),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1783),
.B(n_1690),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_L g2058 ( 
.A(n_2014),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1775),
.B(n_2037),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1763),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1783),
.B(n_1686),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1903),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1798),
.B(n_1531),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2037),
.B(n_1700),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1903),
.Y(n_2065)
);

NAND3xp33_ASAP7_75t_L g2066 ( 
.A(n_1941),
.B(n_1548),
.C(n_1652),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1944),
.B(n_1957),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1944),
.B(n_1686),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1766),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1905),
.Y(n_2070)
);

OR2x6_ASAP7_75t_L g2071 ( 
.A(n_1765),
.B(n_1738),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1766),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1776),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_1844),
.A2(n_1501),
.B1(n_1586),
.B2(n_1686),
.Y(n_2074)
);

INVx3_ASAP7_75t_L g2075 ( 
.A(n_1831),
.Y(n_2075)
);

AOI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_1851),
.A2(n_1501),
.B1(n_1586),
.B2(n_1686),
.Y(n_2076)
);

NAND2xp33_ASAP7_75t_SL g2077 ( 
.A(n_1866),
.B(n_1690),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_1957),
.B(n_1960),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2044),
.B(n_1742),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1905),
.Y(n_2080)
);

NOR2x1p5_ASAP7_75t_L g2081 ( 
.A(n_1768),
.B(n_1522),
.Y(n_2081)
);

INVx11_ASAP7_75t_L g2082 ( 
.A(n_1833),
.Y(n_2082)
);

NOR2x1p5_ASAP7_75t_L g2083 ( 
.A(n_1883),
.B(n_1522),
.Y(n_2083)
);

INVx2_ASAP7_75t_SL g2084 ( 
.A(n_1945),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1960),
.B(n_1739),
.Y(n_2085)
);

INVxp67_ASAP7_75t_SL g2086 ( 
.A(n_2014),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1776),
.Y(n_2087)
);

BUFx3_ASAP7_75t_L g2088 ( 
.A(n_1859),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1789),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1911),
.Y(n_2090)
);

NAND2xp33_ASAP7_75t_L g2091 ( 
.A(n_1932),
.B(n_1586),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1911),
.Y(n_2092)
);

OR2x2_ASAP7_75t_L g2093 ( 
.A(n_1956),
.B(n_1639),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_1831),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1789),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_1859),
.Y(n_2096)
);

BUFx6f_ASAP7_75t_L g2097 ( 
.A(n_2014),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1924),
.B(n_1690),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_SL g2099 ( 
.A(n_1784),
.B(n_1523),
.Y(n_2099)
);

INVxp33_ASAP7_75t_L g2100 ( 
.A(n_1998),
.Y(n_2100)
);

OAI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_1851),
.A2(n_1684),
.B1(n_1694),
.B2(n_1677),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1924),
.B(n_1692),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1918),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1918),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1799),
.Y(n_2105)
);

HB1xp67_ASAP7_75t_L g2106 ( 
.A(n_1865),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2044),
.B(n_1742),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_1991),
.B(n_1964),
.Y(n_2108)
);

INVx2_ASAP7_75t_SL g2109 ( 
.A(n_1942),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1934),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1934),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_1977),
.B(n_1634),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1948),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1948),
.Y(n_2114)
);

INVx2_ASAP7_75t_SL g2115 ( 
.A(n_2003),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1924),
.B(n_1692),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1949),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1924),
.B(n_1692),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1799),
.Y(n_2119)
);

BUFx6f_ASAP7_75t_L g2120 ( 
.A(n_2014),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1949),
.Y(n_2121)
);

INVx5_ASAP7_75t_L g2122 ( 
.A(n_1932),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1968),
.B(n_1504),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1991),
.B(n_1739),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1950),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1964),
.B(n_1739),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2023),
.B(n_1739),
.Y(n_2127)
);

OR2x6_ASAP7_75t_L g2128 ( 
.A(n_1827),
.B(n_1738),
.Y(n_2128)
);

CKINVDCx20_ASAP7_75t_R g2129 ( 
.A(n_1843),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1788),
.B(n_1695),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1805),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1950),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_1855),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1951),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1843),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1805),
.Y(n_2136)
);

INVx2_ASAP7_75t_SL g2137 ( 
.A(n_1855),
.Y(n_2137)
);

BUFx12f_ASAP7_75t_L g2138 ( 
.A(n_1833),
.Y(n_2138)
);

BUFx4f_ASAP7_75t_L g2139 ( 
.A(n_1748),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2023),
.B(n_1586),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1951),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_1977),
.B(n_1634),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_1968),
.B(n_1680),
.Y(n_2143)
);

INVx1_ASAP7_75t_SL g2144 ( 
.A(n_1904),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1889),
.B(n_1586),
.Y(n_2145)
);

OR2x6_ASAP7_75t_L g2146 ( 
.A(n_1867),
.B(n_1738),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1757),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_1751),
.Y(n_2148)
);

OR2x6_ASAP7_75t_L g2149 ( 
.A(n_1878),
.B(n_1692),
.Y(n_2149)
);

BUFx2_ASAP7_75t_L g2150 ( 
.A(n_1764),
.Y(n_2150)
);

INVx4_ASAP7_75t_L g2151 ( 
.A(n_1748),
.Y(n_2151)
);

INVx2_ASAP7_75t_SL g2152 ( 
.A(n_1855),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1758),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_1752),
.B(n_1680),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1808),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1760),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_1833),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_1751),
.Y(n_2158)
);

AND2x6_ASAP7_75t_L g2159 ( 
.A(n_1892),
.B(n_1711),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_1752),
.B(n_1680),
.Y(n_2160)
);

INVx2_ASAP7_75t_SL g2161 ( 
.A(n_1858),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_1935),
.B(n_1711),
.Y(n_2162)
);

INVx2_ASAP7_75t_SL g2163 ( 
.A(n_1858),
.Y(n_2163)
);

INVx3_ASAP7_75t_L g2164 ( 
.A(n_1751),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1808),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1761),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1896),
.B(n_1546),
.Y(n_2167)
);

BUFx6f_ASAP7_75t_L g2168 ( 
.A(n_2015),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_1892),
.A2(n_1719),
.B1(n_1733),
.B2(n_1729),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1813),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1935),
.B(n_1711),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1762),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1813),
.Y(n_2173)
);

BUFx6f_ASAP7_75t_L g2174 ( 
.A(n_2015),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_1751),
.Y(n_2175)
);

AND3x2_ASAP7_75t_L g2176 ( 
.A(n_1849),
.B(n_1728),
.C(n_1667),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1785),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1935),
.B(n_1711),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1820),
.Y(n_2179)
);

OR2x6_ASAP7_75t_L g2180 ( 
.A(n_1764),
.B(n_1718),
.Y(n_2180)
);

INVx4_ASAP7_75t_L g2181 ( 
.A(n_1748),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1908),
.B(n_1655),
.Y(n_2182)
);

BUFx3_ASAP7_75t_L g2183 ( 
.A(n_2006),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1820),
.Y(n_2184)
);

NAND2xp33_ASAP7_75t_L g2185 ( 
.A(n_1932),
.B(n_1718),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1767),
.Y(n_2186)
);

INVx1_ASAP7_75t_SL g2187 ( 
.A(n_1809),
.Y(n_2187)
);

AOI22xp33_ASAP7_75t_L g2188 ( 
.A1(n_1895),
.A2(n_1719),
.B1(n_1733),
.B2(n_1729),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1821),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_1849),
.B(n_1703),
.Y(n_2190)
);

BUFx4f_ASAP7_75t_L g2191 ( 
.A(n_2006),
.Y(n_2191)
);

INVx2_ASAP7_75t_SL g2192 ( 
.A(n_1858),
.Y(n_2192)
);

INVx4_ASAP7_75t_L g2193 ( 
.A(n_2006),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1860),
.B(n_1657),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1821),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1772),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1824),
.Y(n_2197)
);

INVx4_ASAP7_75t_L g2198 ( 
.A(n_1935),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1824),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1773),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_1982),
.B(n_1718),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1780),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1938),
.B(n_1695),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1863),
.B(n_1539),
.Y(n_2204)
);

BUFx3_ASAP7_75t_L g2205 ( 
.A(n_2041),
.Y(n_2205)
);

INVx2_ASAP7_75t_SL g2206 ( 
.A(n_2021),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1781),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_1877),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_1974),
.B(n_1703),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1953),
.Y(n_2210)
);

BUFx6f_ASAP7_75t_L g2211 ( 
.A(n_2015),
.Y(n_2211)
);

INVx3_ASAP7_75t_L g2212 ( 
.A(n_1785),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1782),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_SL g2214 ( 
.A(n_2009),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_1982),
.B(n_1718),
.Y(n_2215)
);

OR2x6_ASAP7_75t_L g2216 ( 
.A(n_2045),
.B(n_1727),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1786),
.Y(n_2217)
);

INVx3_ASAP7_75t_L g2218 ( 
.A(n_1785),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1982),
.B(n_1727),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_1771),
.A2(n_1702),
.B1(n_1638),
.B2(n_1695),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1969),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_1800),
.B(n_1832),
.Y(n_2222)
);

INVx5_ASAP7_75t_L g2223 ( 
.A(n_1932),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_L g2224 ( 
.A(n_1800),
.B(n_1703),
.Y(n_2224)
);

INVxp33_ASAP7_75t_L g2225 ( 
.A(n_1961),
.Y(n_2225)
);

INVxp33_ASAP7_75t_L g2226 ( 
.A(n_2036),
.Y(n_2226)
);

INVxp67_ASAP7_75t_SL g2227 ( 
.A(n_2015),
.Y(n_2227)
);

INVxp67_ASAP7_75t_L g2228 ( 
.A(n_2036),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1971),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1953),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1848),
.B(n_1539),
.Y(n_2231)
);

XOR2xp5_ASAP7_75t_L g2232 ( 
.A(n_1818),
.B(n_1184),
.Y(n_2232)
);

NAND2xp33_ASAP7_75t_SL g2233 ( 
.A(n_1771),
.B(n_1727),
.Y(n_2233)
);

INVx5_ASAP7_75t_L g2234 ( 
.A(n_1932),
.Y(n_2234)
);

INVx4_ASAP7_75t_L g2235 ( 
.A(n_1982),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1965),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_1810),
.B(n_1713),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1975),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1976),
.B(n_1587),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_1785),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_1832),
.B(n_1876),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1965),
.Y(n_2242)
);

AND2x6_ASAP7_75t_L g2243 ( 
.A(n_1895),
.B(n_1727),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_1777),
.B(n_1587),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1978),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1876),
.B(n_1910),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1980),
.B(n_1733),
.Y(n_2247)
);

INVx1_ASAP7_75t_SL g2248 ( 
.A(n_1814),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1985),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_1910),
.B(n_1710),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1985),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1981),
.B(n_1734),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_1810),
.B(n_1713),
.Y(n_2253)
);

AND3x1_ASAP7_75t_L g2254 ( 
.A(n_1921),
.B(n_1696),
.C(n_1720),
.Y(n_2254)
);

BUFx10_ASAP7_75t_L g2255 ( 
.A(n_1777),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1987),
.B(n_1734),
.Y(n_2256)
);

BUFx10_ASAP7_75t_L g2257 ( 
.A(n_1777),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1986),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1995),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1986),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1992),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1992),
.Y(n_2262)
);

AOI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_2018),
.A2(n_1734),
.B1(n_1741),
.B2(n_1593),
.Y(n_2263)
);

AND2x6_ASAP7_75t_L g2264 ( 
.A(n_1834),
.B(n_1735),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1996),
.Y(n_2265)
);

BUFx3_ASAP7_75t_L g2266 ( 
.A(n_2041),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2002),
.B(n_1741),
.Y(n_2267)
);

INVx4_ASAP7_75t_SL g2268 ( 
.A(n_2018),
.Y(n_2268)
);

NAND2xp33_ASAP7_75t_L g2269 ( 
.A(n_2018),
.B(n_2035),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2005),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_1846),
.Y(n_2271)
);

BUFx3_ASAP7_75t_L g2272 ( 
.A(n_2041),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2012),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_1983),
.B(n_1735),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2013),
.B(n_1741),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2017),
.B(n_2019),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2020),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_1983),
.B(n_1735),
.Y(n_2278)
);

AOI22xp33_ASAP7_75t_L g2279 ( 
.A1(n_2018),
.A2(n_1593),
.B1(n_911),
.B2(n_1020),
.Y(n_2279)
);

OAI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_1914),
.A2(n_1712),
.B1(n_1714),
.B2(n_1706),
.Y(n_2280)
);

AND2x6_ASAP7_75t_L g2281 ( 
.A(n_1834),
.B(n_1837),
.Y(n_2281)
);

INVx2_ASAP7_75t_SL g2282 ( 
.A(n_1804),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1787),
.Y(n_2283)
);

OAI22xp33_ASAP7_75t_L g2284 ( 
.A1(n_1920),
.A2(n_1925),
.B1(n_1926),
.B2(n_1923),
.Y(n_2284)
);

INVx4_ASAP7_75t_L g2285 ( 
.A(n_1983),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_1996),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1790),
.Y(n_2287)
);

BUFx3_ASAP7_75t_L g2288 ( 
.A(n_1877),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1792),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2007),
.Y(n_2290)
);

CKINVDCx5p33_ASAP7_75t_R g2291 ( 
.A(n_1877),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2007),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_1873),
.B(n_1713),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_1828),
.B(n_1710),
.Y(n_2294)
);

CKINVDCx5p33_ASAP7_75t_R g2295 ( 
.A(n_1899),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_2011),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1794),
.Y(n_2297)
);

CKINVDCx20_ASAP7_75t_R g2298 ( 
.A(n_1807),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2011),
.Y(n_2299)
);

BUFx10_ASAP7_75t_L g2300 ( 
.A(n_1804),
.Y(n_2300)
);

OR2x6_ASAP7_75t_L g2301 ( 
.A(n_1806),
.B(n_1735),
.Y(n_2301)
);

INVx1_ASAP7_75t_SL g2302 ( 
.A(n_1807),
.Y(n_2302)
);

INVx5_ASAP7_75t_L g2303 ( 
.A(n_2018),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2022),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1795),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2022),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2026),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_1983),
.B(n_1710),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_1984),
.B(n_1706),
.Y(n_2309)
);

INVx1_ASAP7_75t_SL g2310 ( 
.A(n_1804),
.Y(n_2310)
);

AOI22xp33_ASAP7_75t_L g2311 ( 
.A1(n_2035),
.A2(n_1880),
.B1(n_1861),
.B2(n_1862),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1796),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1797),
.B(n_1674),
.Y(n_2313)
);

NOR2x1p5_ASAP7_75t_L g2314 ( 
.A(n_1927),
.B(n_1664),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1801),
.Y(n_2315)
);

NOR2x1p5_ASAP7_75t_L g2316 ( 
.A(n_1929),
.B(n_1664),
.Y(n_2316)
);

BUFx3_ASAP7_75t_L g2317 ( 
.A(n_2027),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2026),
.Y(n_2318)
);

AOI21x1_ASAP7_75t_L g2319 ( 
.A1(n_1774),
.A2(n_1822),
.B(n_1812),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2042),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1802),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_1984),
.B(n_1712),
.Y(n_2322)
);

OR2x2_ASAP7_75t_L g2323 ( 
.A(n_2009),
.B(n_1740),
.Y(n_2323)
);

INVx2_ASAP7_75t_SL g2324 ( 
.A(n_1873),
.Y(n_2324)
);

BUFx6f_ASAP7_75t_L g2325 ( 
.A(n_2016),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1803),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2042),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2046),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2046),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1811),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1815),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1817),
.B(n_1722),
.Y(n_2332)
);

NAND2xp33_ASAP7_75t_SL g2333 ( 
.A(n_1779),
.B(n_1714),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2047),
.Y(n_2334)
);

INVx4_ASAP7_75t_L g2335 ( 
.A(n_1984),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2047),
.Y(n_2336)
);

BUFx8_ASAP7_75t_SL g2337 ( 
.A(n_2009),
.Y(n_2337)
);

INVx3_ASAP7_75t_L g2338 ( 
.A(n_1826),
.Y(n_2338)
);

AOI22xp33_ASAP7_75t_L g2339 ( 
.A1(n_2035),
.A2(n_1052),
.B1(n_909),
.B2(n_1575),
.Y(n_2339)
);

NAND2xp33_ASAP7_75t_R g2340 ( 
.A(n_1886),
.B(n_1601),
.Y(n_2340)
);

INVx1_ASAP7_75t_SL g2341 ( 
.A(n_1873),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1819),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_1984),
.B(n_1724),
.Y(n_2343)
);

CKINVDCx5p33_ASAP7_75t_R g2344 ( 
.A(n_1806),
.Y(n_2344)
);

NOR3xp33_ASAP7_75t_L g2345 ( 
.A(n_1907),
.B(n_1704),
.C(n_1669),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_1853),
.B(n_1724),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_1749),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1823),
.Y(n_2348)
);

BUFx3_ASAP7_75t_L g2349 ( 
.A(n_2029),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_1836),
.B(n_1726),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_2222),
.B(n_1601),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2190),
.B(n_1828),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2222),
.B(n_1608),
.Y(n_2353)
);

NOR2xp67_ASAP7_75t_L g2354 ( 
.A(n_2084),
.B(n_1664),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2231),
.B(n_2035),
.Y(n_2355)
);

BUFx5_ASAP7_75t_L g2356 ( 
.A(n_2281),
.Y(n_2356)
);

INVxp67_ASAP7_75t_L g2357 ( 
.A(n_2150),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2049),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2226),
.B(n_1608),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2067),
.B(n_2035),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2067),
.B(n_1816),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2078),
.B(n_1816),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_2190),
.B(n_1726),
.Y(n_2363)
);

CKINVDCx20_ASAP7_75t_R g2364 ( 
.A(n_2129),
.Y(n_2364)
);

INVx4_ASAP7_75t_L g2365 ( 
.A(n_2139),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2055),
.Y(n_2366)
);

OR2x2_ASAP7_75t_L g2367 ( 
.A(n_2063),
.B(n_1609),
.Y(n_2367)
);

NOR3xp33_ASAP7_75t_L g2368 ( 
.A(n_2066),
.B(n_1666),
.C(n_1638),
.Y(n_2368)
);

INVx2_ASAP7_75t_SL g2369 ( 
.A(n_2109),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2049),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2078),
.B(n_1880),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2228),
.B(n_1829),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2056),
.Y(n_2373)
);

NAND2xp33_ASAP7_75t_SL g2374 ( 
.A(n_2226),
.B(n_1731),
.Y(n_2374)
);

NOR3xp33_ASAP7_75t_L g2375 ( 
.A(n_2224),
.B(n_1723),
.C(n_1715),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2062),
.Y(n_2376)
);

INVxp67_ASAP7_75t_L g2377 ( 
.A(n_2093),
.Y(n_2377)
);

BUFx6f_ASAP7_75t_L g2378 ( 
.A(n_2058),
.Y(n_2378)
);

INVx2_ASAP7_75t_SL g2379 ( 
.A(n_2271),
.Y(n_2379)
);

INVx2_ASAP7_75t_SL g2380 ( 
.A(n_2071),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_2058),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2059),
.B(n_1677),
.Y(n_2382)
);

BUFx6f_ASAP7_75t_L g2383 ( 
.A(n_2058),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2228),
.B(n_1835),
.Y(n_2384)
);

BUFx6f_ASAP7_75t_SL g2385 ( 
.A(n_2288),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2065),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2204),
.B(n_1838),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2050),
.Y(n_2388)
);

NOR2xp33_ASAP7_75t_L g2389 ( 
.A(n_2167),
.B(n_1609),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_2058),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2070),
.Y(n_2391)
);

NAND2x1_ASAP7_75t_L g2392 ( 
.A(n_2198),
.B(n_1966),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2182),
.B(n_1701),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_2224),
.B(n_1731),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2050),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_2225),
.B(n_1701),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2060),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_SL g2398 ( 
.A(n_2203),
.B(n_1737),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2241),
.B(n_1841),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2060),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2241),
.B(n_2108),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2073),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2073),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2087),
.Y(n_2404)
);

BUFx6f_ASAP7_75t_L g2405 ( 
.A(n_2097),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2143),
.B(n_1845),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2143),
.B(n_1847),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_2151),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_SL g2409 ( 
.A(n_2154),
.B(n_1737),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2080),
.Y(n_2410)
);

NOR2x1p5_ASAP7_75t_L g2411 ( 
.A(n_2288),
.B(n_1744),
.Y(n_2411)
);

NOR2xp33_ASAP7_75t_L g2412 ( 
.A(n_2225),
.B(n_1523),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2090),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2092),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2087),
.Y(n_2415)
);

NAND3xp33_ASAP7_75t_L g2416 ( 
.A(n_2345),
.B(n_2123),
.C(n_2246),
.Y(n_2416)
);

NOR3xp33_ASAP7_75t_L g2417 ( 
.A(n_2130),
.B(n_1679),
.C(n_1678),
.Y(n_2417)
);

INVx1_ASAP7_75t_SL g2418 ( 
.A(n_2144),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2154),
.B(n_1745),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2160),
.B(n_1850),
.Y(n_2420)
);

INVx2_ASAP7_75t_SL g2421 ( 
.A(n_2071),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2103),
.Y(n_2422)
);

INVxp33_ASAP7_75t_L g2423 ( 
.A(n_2099),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2187),
.B(n_1509),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2246),
.B(n_1852),
.Y(n_2425)
);

NOR3xp33_ASAP7_75t_L g2426 ( 
.A(n_2160),
.B(n_1683),
.C(n_1682),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2095),
.Y(n_2427)
);

NAND2xp33_ASAP7_75t_L g2428 ( 
.A(n_2159),
.B(n_1509),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2095),
.Y(n_2429)
);

AO221x1_ASAP7_75t_L g2430 ( 
.A1(n_2280),
.A2(n_1708),
.B1(n_1721),
.B2(n_1717),
.C(n_1697),
.Y(n_2430)
);

INVx4_ASAP7_75t_L g2431 ( 
.A(n_2139),
.Y(n_2431)
);

OR2x2_ASAP7_75t_L g2432 ( 
.A(n_2248),
.B(n_1684),
.Y(n_2432)
);

INVxp33_ASAP7_75t_L g2433 ( 
.A(n_2237),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2105),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2123),
.B(n_1854),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_2194),
.B(n_1745),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2048),
.B(n_1856),
.Y(n_2437)
);

INVxp33_ASAP7_75t_L g2438 ( 
.A(n_2253),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2048),
.B(n_1857),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2294),
.B(n_1868),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2105),
.Y(n_2441)
);

AO221x1_ASAP7_75t_L g2442 ( 
.A1(n_2284),
.A2(n_1685),
.B1(n_1694),
.B2(n_1709),
.C(n_1466),
.Y(n_2442)
);

NAND3xp33_ASAP7_75t_L g2443 ( 
.A(n_2345),
.B(n_1743),
.C(n_1988),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2294),
.B(n_1869),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2104),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_2244),
.B(n_1744),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2119),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2110),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2119),
.Y(n_2449)
);

NOR2xp33_ASAP7_75t_L g2450 ( 
.A(n_2100),
.B(n_1346),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2111),
.Y(n_2451)
);

BUFx5_ASAP7_75t_L g2452 ( 
.A(n_2281),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2052),
.B(n_1871),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2131),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2131),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2100),
.B(n_1355),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2136),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2250),
.B(n_1872),
.Y(n_2458)
);

INVxp67_ASAP7_75t_L g2459 ( 
.A(n_2053),
.Y(n_2459)
);

INVxp67_ASAP7_75t_L g2460 ( 
.A(n_2053),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2136),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2199),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_2209),
.B(n_1369),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2113),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2250),
.B(n_1882),
.Y(n_2465)
);

INVxp33_ASAP7_75t_L g2466 ( 
.A(n_2323),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_R g2467 ( 
.A(n_2135),
.B(n_1184),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2239),
.B(n_1884),
.Y(n_2468)
);

NOR3xp33_ASAP7_75t_L g2469 ( 
.A(n_2332),
.B(n_1716),
.C(n_1736),
.Y(n_2469)
);

INVxp67_ASAP7_75t_L g2470 ( 
.A(n_2106),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2199),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2114),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2117),
.Y(n_2473)
);

OR2x6_ASAP7_75t_L g2474 ( 
.A(n_2071),
.B(n_1597),
.Y(n_2474)
);

OR2x2_ASAP7_75t_L g2475 ( 
.A(n_2064),
.B(n_1722),
.Y(n_2475)
);

NOR3xp33_ASAP7_75t_L g2476 ( 
.A(n_2209),
.B(n_1595),
.C(n_1931),
.Y(n_2476)
);

BUFx2_ASAP7_75t_L g2477 ( 
.A(n_2295),
.Y(n_2477)
);

AOI221xp5_ASAP7_75t_L g2478 ( 
.A1(n_2254),
.A2(n_506),
.B1(n_696),
.B2(n_498),
.C(n_496),
.Y(n_2478)
);

A2O1A1Ixp33_ASAP7_75t_L g2479 ( 
.A1(n_2220),
.A2(n_1937),
.B(n_1939),
.C(n_1930),
.Y(n_2479)
);

NOR2xp33_ASAP7_75t_L g2480 ( 
.A(n_2115),
.B(n_1369),
.Y(n_2480)
);

AND2x6_ASAP7_75t_L g2481 ( 
.A(n_2074),
.B(n_2076),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2121),
.Y(n_2482)
);

INVx5_ASAP7_75t_L g2483 ( 
.A(n_2159),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2079),
.B(n_1887),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2107),
.B(n_1888),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2125),
.Y(n_2486)
);

NOR2xp33_ASAP7_75t_L g2487 ( 
.A(n_2344),
.B(n_1370),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2210),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2210),
.Y(n_2489)
);

OR2x2_ASAP7_75t_L g2490 ( 
.A(n_2106),
.B(n_1722),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2057),
.B(n_1890),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2057),
.B(n_1370),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2206),
.B(n_1891),
.Y(n_2493)
);

NAND2xp33_ASAP7_75t_L g2494 ( 
.A(n_2159),
.B(n_1993),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2132),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2230),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2341),
.B(n_1373),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2283),
.B(n_1893),
.Y(n_2498)
);

NAND2xp33_ASAP7_75t_L g2499 ( 
.A(n_2159),
.B(n_1997),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2244),
.B(n_1746),
.Y(n_2500)
);

XOR2xp5_ASAP7_75t_L g2501 ( 
.A(n_2232),
.B(n_1212),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2293),
.B(n_1746),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2134),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2230),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2141),
.Y(n_2505)
);

INVxp67_ASAP7_75t_L g2506 ( 
.A(n_2128),
.Y(n_2506)
);

AND2x2_ASAP7_75t_SL g2507 ( 
.A(n_2185),
.B(n_1483),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_2101),
.B(n_1746),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2287),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2236),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2236),
.Y(n_2511)
);

NOR2xp67_ASAP7_75t_L g2512 ( 
.A(n_2313),
.B(n_1643),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2289),
.B(n_1894),
.Y(n_2513)
);

NOR2xp33_ASAP7_75t_L g2514 ( 
.A(n_2302),
.B(n_1373),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2310),
.B(n_1383),
.Y(n_2515)
);

AOI221xp5_ASAP7_75t_L g2516 ( 
.A1(n_2101),
.A2(n_711),
.B1(n_717),
.B2(n_710),
.C(n_696),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_2097),
.Y(n_2517)
);

BUFx3_ASAP7_75t_L g2518 ( 
.A(n_2128),
.Y(n_2518)
);

AND2x6_ASAP7_75t_SL g2519 ( 
.A(n_2128),
.B(n_1498),
.Y(n_2519)
);

NOR3xp33_ASAP7_75t_L g2520 ( 
.A(n_2324),
.B(n_1485),
.C(n_1498),
.Y(n_2520)
);

NOR2xp67_ASAP7_75t_L g2521 ( 
.A(n_2297),
.B(n_1643),
.Y(n_2521)
);

NOR3xp33_ASAP7_75t_L g2522 ( 
.A(n_2282),
.B(n_1943),
.C(n_1940),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2305),
.B(n_1897),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2312),
.B(n_1898),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2315),
.B(n_1901),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2321),
.B(n_1909),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_2133),
.B(n_1643),
.Y(n_2527)
);

NOR3xp33_ASAP7_75t_L g2528 ( 
.A(n_2233),
.B(n_1947),
.C(n_1946),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2326),
.B(n_1912),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2330),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2331),
.B(n_1913),
.Y(n_2531)
);

OR2x2_ASAP7_75t_L g2532 ( 
.A(n_2146),
.B(n_2031),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2342),
.B(n_1928),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2348),
.B(n_1928),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2242),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2346),
.B(n_1928),
.Y(n_2536)
);

INVxp67_ASAP7_75t_SL g2537 ( 
.A(n_2311),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2061),
.B(n_1837),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2242),
.Y(n_2539)
);

OR2x6_ASAP7_75t_L g2540 ( 
.A(n_2146),
.B(n_2149),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2085),
.B(n_1861),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2068),
.B(n_1862),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2249),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2249),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2258),
.Y(n_2545)
);

NOR2xp67_ASAP7_75t_L g2546 ( 
.A(n_2137),
.B(n_2032),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_SL g2547 ( 
.A(n_2152),
.B(n_2010),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2281),
.B(n_1870),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2258),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2281),
.B(n_1870),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2260),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2260),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2261),
.Y(n_2553)
);

CKINVDCx20_ASAP7_75t_R g2554 ( 
.A(n_2337),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_SL g2555 ( 
.A(n_2161),
.B(n_2010),
.Y(n_2555)
);

INVx2_ASAP7_75t_SL g2556 ( 
.A(n_2146),
.Y(n_2556)
);

INVx1_ASAP7_75t_SL g2557 ( 
.A(n_2180),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2281),
.B(n_1874),
.Y(n_2558)
);

OR2x2_ASAP7_75t_L g2559 ( 
.A(n_2163),
.B(n_2034),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2124),
.B(n_1874),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2054),
.B(n_1875),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_2097),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2261),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2262),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_SL g2565 ( 
.A(n_2192),
.B(n_2010),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2262),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_SL g2567 ( 
.A(n_2112),
.B(n_2024),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2112),
.B(n_2024),
.Y(n_2568)
);

INVx1_ASAP7_75t_SL g2569 ( 
.A(n_2180),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2054),
.B(n_1875),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_SL g2571 ( 
.A(n_2142),
.B(n_2024),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2265),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_2346),
.B(n_1383),
.Y(n_2573)
);

INVx2_ASAP7_75t_SL g2574 ( 
.A(n_2180),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_SL g2575 ( 
.A(n_2142),
.B(n_1952),
.Y(n_2575)
);

OR2x2_ASAP7_75t_SL g2576 ( 
.A(n_2216),
.B(n_1385),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2301),
.B(n_1385),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2265),
.B(n_1879),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2286),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2286),
.Y(n_2580)
);

AND2x6_ASAP7_75t_SL g2581 ( 
.A(n_2149),
.B(n_2216),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2290),
.B(n_1879),
.Y(n_2582)
);

BUFx3_ASAP7_75t_L g2583 ( 
.A(n_2149),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2301),
.B(n_1398),
.Y(n_2584)
);

NAND2xp33_ASAP7_75t_L g2585 ( 
.A(n_2159),
.B(n_2004),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2290),
.B(n_1885),
.Y(n_2586)
);

INVxp67_ASAP7_75t_L g2587 ( 
.A(n_2337),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2301),
.B(n_1398),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2327),
.B(n_1885),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2088),
.B(n_1399),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_SL g2591 ( 
.A(n_2191),
.B(n_1954),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2088),
.B(n_1399),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2327),
.B(n_1955),
.Y(n_2593)
);

AND3x1_ASAP7_75t_L g2594 ( 
.A(n_2147),
.B(n_1962),
.C(n_1958),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2096),
.B(n_1408),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2328),
.B(n_1963),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2317),
.B(n_1967),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2509),
.Y(n_2598)
);

AOI22xp33_ASAP7_75t_L g2599 ( 
.A1(n_2416),
.A2(n_2233),
.B1(n_2216),
.B2(n_2077),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2530),
.Y(n_2600)
);

BUFx3_ASAP7_75t_L g2601 ( 
.A(n_2379),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2358),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2366),
.Y(n_2603)
);

OAI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2351),
.A2(n_2311),
.B1(n_2191),
.B2(n_2223),
.Y(n_2604)
);

INVxp67_ASAP7_75t_L g2605 ( 
.A(n_2382),
.Y(n_2605)
);

NAND3xp33_ASAP7_75t_L g2606 ( 
.A(n_2353),
.B(n_1470),
.C(n_1461),
.Y(n_2606)
);

INVxp67_ASAP7_75t_L g2607 ( 
.A(n_2432),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2373),
.Y(n_2608)
);

AOI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2368),
.A2(n_2077),
.B1(n_2156),
.B2(n_2153),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2492),
.B(n_2096),
.Y(n_2610)
);

NAND2x1_ASAP7_75t_L g2611 ( 
.A(n_2408),
.B(n_2198),
.Y(n_2611)
);

OR2x2_ASAP7_75t_L g2612 ( 
.A(n_2367),
.B(n_2040),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2376),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2401),
.B(n_2349),
.Y(n_2614)
);

OR2x2_ASAP7_75t_L g2615 ( 
.A(n_2475),
.B(n_2166),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_SL g2616 ( 
.A(n_2389),
.B(n_2255),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2436),
.B(n_2349),
.Y(n_2617)
);

NOR2xp33_ASAP7_75t_L g2618 ( 
.A(n_2393),
.B(n_1408),
.Y(n_2618)
);

O2A1O1Ixp33_ASAP7_75t_L g2619 ( 
.A1(n_2361),
.A2(n_2284),
.B(n_1999),
.C(n_1989),
.Y(n_2619)
);

INVx2_ASAP7_75t_SL g2620 ( 
.A(n_2369),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2399),
.B(n_2317),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2502),
.B(n_2255),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2370),
.Y(n_2623)
);

OAI221xp5_ASAP7_75t_L g2624 ( 
.A1(n_2478),
.A2(n_2279),
.B1(n_1753),
.B2(n_1756),
.C(n_1754),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2388),
.Y(n_2625)
);

AOI21xp5_ASAP7_75t_L g2626 ( 
.A1(n_2494),
.A2(n_2091),
.B(n_2263),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2361),
.B(n_2172),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_L g2628 ( 
.A(n_2362),
.B(n_2298),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2386),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2391),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2362),
.B(n_2186),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2410),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2395),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2413),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2435),
.B(n_2196),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2359),
.B(n_2257),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2397),
.Y(n_2637)
);

AOI22xp5_ASAP7_75t_L g2638 ( 
.A1(n_2463),
.A2(n_1419),
.B1(n_1422),
.B2(n_1417),
.Y(n_2638)
);

NOR3xp33_ASAP7_75t_L g2639 ( 
.A(n_2443),
.B(n_2145),
.C(n_1999),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2435),
.B(n_2200),
.Y(n_2640)
);

NOR3xp33_ASAP7_75t_L g2641 ( 
.A(n_2375),
.B(n_1989),
.C(n_2350),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2400),
.Y(n_2642)
);

NAND2xp33_ASAP7_75t_L g2643 ( 
.A(n_2483),
.B(n_2243),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2414),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2387),
.B(n_2202),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2402),
.Y(n_2646)
);

NOR2xp33_ASAP7_75t_L g2647 ( 
.A(n_2433),
.B(n_1417),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_SL g2648 ( 
.A(n_2365),
.B(n_1212),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2425),
.B(n_2468),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2450),
.A2(n_1422),
.B1(n_1423),
.B2(n_1419),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2422),
.Y(n_2651)
);

AOI22xp33_ASAP7_75t_L g2652 ( 
.A1(n_2508),
.A2(n_2213),
.B1(n_2217),
.B2(n_2207),
.Y(n_2652)
);

INVx2_ASAP7_75t_SL g2653 ( 
.A(n_2518),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2425),
.B(n_2221),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2445),
.Y(n_2655)
);

NOR2xp33_ASAP7_75t_L g2656 ( 
.A(n_2438),
.B(n_1423),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2403),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2484),
.B(n_2229),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2485),
.B(n_2238),
.Y(n_2659)
);

AND2x4_ASAP7_75t_L g2660 ( 
.A(n_2365),
.B(n_2314),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_L g2661 ( 
.A(n_2424),
.B(n_1428),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_2466),
.B(n_1428),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2404),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2377),
.B(n_1433),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2453),
.B(n_2245),
.Y(n_2665)
);

AOI22xp33_ASAP7_75t_L g2666 ( 
.A1(n_2430),
.A2(n_2270),
.B1(n_2273),
.B2(n_2259),
.Y(n_2666)
);

AOI21xp5_ASAP7_75t_L g2667 ( 
.A1(n_2499),
.A2(n_2263),
.B(n_2269),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2352),
.B(n_2277),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2415),
.Y(n_2669)
);

OAI22xp5_ASAP7_75t_SL g2670 ( 
.A1(n_2576),
.A2(n_1437),
.B1(n_1443),
.B2(n_1433),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2427),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2429),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2372),
.B(n_2126),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2357),
.B(n_1437),
.Y(n_2674)
);

AOI22xp5_ASAP7_75t_L g2675 ( 
.A1(n_2456),
.A2(n_1445),
.B1(n_1457),
.B2(n_1443),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2448),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2372),
.B(n_2127),
.Y(n_2677)
);

NOR2xp33_ASAP7_75t_L g2678 ( 
.A(n_2423),
.B(n_1445),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2451),
.Y(n_2679)
);

AOI22xp33_ASAP7_75t_L g2680 ( 
.A1(n_2442),
.A2(n_2276),
.B1(n_2350),
.B2(n_2279),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2464),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2434),
.Y(n_2682)
);

AOI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2585),
.A2(n_2188),
.B(n_2169),
.Y(n_2683)
);

INVx8_ASAP7_75t_L g2684 ( 
.A(n_2540),
.Y(n_2684)
);

INVx4_ASAP7_75t_L g2685 ( 
.A(n_2431),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2440),
.B(n_2075),
.Y(n_2686)
);

AOI22xp33_ASAP7_75t_L g2687 ( 
.A1(n_2440),
.A2(n_2316),
.B1(n_2094),
.B2(n_2075),
.Y(n_2687)
);

NOR2xp33_ASAP7_75t_L g2688 ( 
.A(n_2514),
.B(n_1457),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2472),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2444),
.B(n_2094),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2473),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2444),
.B(n_1916),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2441),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2447),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_L g2695 ( 
.A(n_2573),
.B(n_1215),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2449),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2482),
.Y(n_2697)
);

OAI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2537),
.A2(n_2122),
.B1(n_2234),
.B2(n_2223),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2454),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_L g2700 ( 
.A(n_2418),
.B(n_1215),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2384),
.B(n_1936),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2486),
.Y(n_2702)
);

AOI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2480),
.A2(n_1222),
.B1(n_1255),
.B2(n_1217),
.Y(n_2703)
);

AND2x6_ASAP7_75t_SL g2704 ( 
.A(n_2487),
.B(n_2082),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2455),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2457),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_SL g2707 ( 
.A(n_2418),
.B(n_2257),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2461),
.Y(n_2708)
);

AOI21xp5_ASAP7_75t_L g2709 ( 
.A1(n_2363),
.A2(n_2188),
.B(n_2169),
.Y(n_2709)
);

NOR3xp33_ASAP7_75t_L g2710 ( 
.A(n_2396),
.B(n_1970),
.C(n_2140),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2406),
.B(n_2098),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2462),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_L g2713 ( 
.A(n_2497),
.B(n_1217),
.Y(n_2713)
);

NOR2xp33_ASAP7_75t_L g2714 ( 
.A(n_2515),
.B(n_1222),
.Y(n_2714)
);

AOI21xp5_ASAP7_75t_L g2715 ( 
.A1(n_2561),
.A2(n_2223),
.B(n_2122),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_L g2716 ( 
.A(n_2412),
.B(n_1255),
.Y(n_2716)
);

INVxp67_ASAP7_75t_SL g2717 ( 
.A(n_2561),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2471),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2477),
.B(n_2300),
.Y(n_2719)
);

AOI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2570),
.A2(n_2223),
.B(n_2122),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2488),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2407),
.B(n_2098),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2490),
.B(n_2300),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2495),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2420),
.B(n_2102),
.Y(n_2725)
);

CKINVDCx5p33_ASAP7_75t_R g2726 ( 
.A(n_2467),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2489),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2496),
.Y(n_2728)
);

HB1xp67_ASAP7_75t_L g2729 ( 
.A(n_2459),
.Y(n_2729)
);

AOI22x1_ASAP7_75t_L g2730 ( 
.A1(n_2503),
.A2(n_2051),
.B1(n_2072),
.B2(n_2069),
.Y(n_2730)
);

AND2x6_ASAP7_75t_SL g2731 ( 
.A(n_2590),
.B(n_1687),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2458),
.B(n_2102),
.Y(n_2732)
);

NOR2xp67_ASAP7_75t_L g2733 ( 
.A(n_2354),
.B(n_2138),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2465),
.B(n_2116),
.Y(n_2734)
);

AOI22xp33_ASAP7_75t_L g2735 ( 
.A1(n_2481),
.A2(n_2374),
.B1(n_2426),
.B2(n_2476),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_L g2736 ( 
.A(n_2498),
.B(n_2116),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2394),
.B(n_1266),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_L g2738 ( 
.A(n_2460),
.B(n_1266),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2470),
.B(n_1272),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_SL g2740 ( 
.A(n_2417),
.B(n_2122),
.Y(n_2740)
);

BUFx8_ASAP7_75t_L g2741 ( 
.A(n_2385),
.Y(n_2741)
);

HB1xp67_ASAP7_75t_L g2742 ( 
.A(n_2548),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2513),
.B(n_2118),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2505),
.Y(n_2744)
);

A2O1A1Ixp33_ASAP7_75t_L g2745 ( 
.A1(n_2409),
.A2(n_2333),
.B(n_2309),
.C(n_2322),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2504),
.Y(n_2746)
);

AOI22xp33_ASAP7_75t_L g2747 ( 
.A1(n_2481),
.A2(n_2162),
.B1(n_2171),
.B2(n_2118),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2469),
.B(n_2234),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2510),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2511),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2535),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2523),
.B(n_2524),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_SL g2753 ( 
.A(n_2507),
.B(n_2234),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2543),
.Y(n_2754)
);

OR2x6_ASAP7_75t_L g2755 ( 
.A(n_2540),
.B(n_2205),
.Y(n_2755)
);

O2A1O1Ixp5_ASAP7_75t_L g2756 ( 
.A1(n_2419),
.A2(n_2308),
.B(n_2322),
.C(n_2309),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2525),
.B(n_2162),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2526),
.B(n_2171),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2398),
.B(n_1272),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_2592),
.B(n_1278),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2529),
.B(n_2531),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_SL g2762 ( 
.A(n_2431),
.B(n_2595),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_SL g2763 ( 
.A(n_2533),
.B(n_2234),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_SL g2764 ( 
.A(n_2364),
.B(n_1278),
.Y(n_2764)
);

INVx4_ASAP7_75t_L g2765 ( 
.A(n_2378),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2534),
.B(n_2178),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2437),
.B(n_2178),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2437),
.B(n_2201),
.Y(n_2768)
);

AND2x2_ASAP7_75t_SL g2769 ( 
.A(n_2594),
.B(n_2151),
.Y(n_2769)
);

INVxp33_ASAP7_75t_L g2770 ( 
.A(n_2577),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_L g2771 ( 
.A(n_2493),
.B(n_2439),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_SL g2772 ( 
.A(n_2597),
.B(n_2303),
.Y(n_2772)
);

AOI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_2481),
.A2(n_2215),
.B1(n_2219),
.B2(n_2201),
.Y(n_2773)
);

AND2x6_ASAP7_75t_L g2774 ( 
.A(n_2408),
.B(n_2347),
.Y(n_2774)
);

HB1xp67_ASAP7_75t_L g2775 ( 
.A(n_2548),
.Y(n_2775)
);

INVxp67_ASAP7_75t_L g2776 ( 
.A(n_2532),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2439),
.B(n_2371),
.Y(n_2777)
);

NOR2xp33_ASAP7_75t_L g2778 ( 
.A(n_2501),
.B(n_1281),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2544),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_L g2780 ( 
.A1(n_2481),
.A2(n_2219),
.B1(n_2274),
.B2(n_2215),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2371),
.B(n_2274),
.Y(n_2781)
);

BUFx3_ASAP7_75t_L g2782 ( 
.A(n_2583),
.Y(n_2782)
);

INVx3_ASAP7_75t_L g2783 ( 
.A(n_2378),
.Y(n_2783)
);

NOR2xp33_ASAP7_75t_L g2784 ( 
.A(n_2500),
.B(n_1281),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2491),
.B(n_2278),
.Y(n_2785)
);

AOI22xp33_ASAP7_75t_L g2786 ( 
.A1(n_2528),
.A2(n_2278),
.B1(n_2343),
.B2(n_2308),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_2584),
.B(n_2303),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2549),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2553),
.Y(n_2789)
);

BUFx5_ASAP7_75t_L g2790 ( 
.A(n_2539),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2567),
.B(n_2568),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2571),
.B(n_1973),
.Y(n_2792)
);

NOR2xp67_ASAP7_75t_L g2793 ( 
.A(n_2587),
.B(n_2157),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2588),
.B(n_2083),
.Y(n_2794)
);

INVx4_ASAP7_75t_L g2795 ( 
.A(n_2685),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2771),
.B(n_2516),
.Y(n_2796)
);

NOR3xp33_ASAP7_75t_L g2797 ( 
.A(n_2618),
.B(n_2446),
.C(n_2520),
.Y(n_2797)
);

OAI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2628),
.A2(n_2540),
.B1(n_2569),
.B2(n_2557),
.Y(n_2798)
);

INVxp33_ASAP7_75t_L g2799 ( 
.A(n_2700),
.Y(n_2799)
);

AOI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2643),
.A2(n_2483),
.B(n_2303),
.Y(n_2800)
);

AND2x4_ASAP7_75t_L g2801 ( 
.A(n_2685),
.B(n_2660),
.Y(n_2801)
);

AOI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2628),
.A2(n_2522),
.B1(n_2536),
.B2(n_2360),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2771),
.B(n_2176),
.Y(n_2803)
);

AOI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2626),
.A2(n_2483),
.B(n_2303),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2713),
.B(n_1284),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2626),
.A2(n_2483),
.B(n_2570),
.Y(n_2806)
);

AOI21xp5_ASAP7_75t_L g2807 ( 
.A1(n_2667),
.A2(n_2479),
.B(n_2355),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2649),
.B(n_2176),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2598),
.Y(n_2809)
);

AND2x4_ASAP7_75t_L g2810 ( 
.A(n_2660),
.B(n_2380),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2752),
.B(n_2559),
.Y(n_2811)
);

INVx4_ASAP7_75t_L g2812 ( 
.A(n_2684),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_L g2813 ( 
.A(n_2714),
.B(n_1284),
.Y(n_2813)
);

OAI22xp5_ASAP7_75t_L g2814 ( 
.A1(n_2661),
.A2(n_2557),
.B1(n_2569),
.B2(n_2474),
.Y(n_2814)
);

AOI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2667),
.A2(n_2355),
.B(n_2428),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2761),
.B(n_2506),
.Y(n_2816)
);

AO21x1_ASAP7_75t_L g2817 ( 
.A1(n_2619),
.A2(n_2360),
.B(n_2343),
.Y(n_2817)
);

AOI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2683),
.A2(n_2333),
.B(n_2538),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2701),
.B(n_2645),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2600),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2605),
.B(n_2614),
.Y(n_2821)
);

AOI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2683),
.A2(n_2538),
.B(n_2227),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2605),
.B(n_2575),
.Y(n_2823)
);

AOI21xp5_ASAP7_75t_L g2824 ( 
.A1(n_2692),
.A2(n_2227),
.B(n_2086),
.Y(n_2824)
);

AOI22xp5_ASAP7_75t_L g2825 ( 
.A1(n_2695),
.A2(n_1293),
.B1(n_1296),
.B2(n_1288),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_SL g2826 ( 
.A(n_2617),
.B(n_2512),
.Y(n_2826)
);

AOI21xp5_ASAP7_75t_L g2827 ( 
.A1(n_2709),
.A2(n_2086),
.B(n_2550),
.Y(n_2827)
);

AOI21xp5_ASAP7_75t_L g2828 ( 
.A1(n_2709),
.A2(n_2604),
.B(n_2715),
.Y(n_2828)
);

A2O1A1Ixp33_ASAP7_75t_L g2829 ( 
.A1(n_2619),
.A2(n_2546),
.B(n_2521),
.C(n_2547),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2665),
.B(n_2556),
.Y(n_2830)
);

NOR2xp33_ASAP7_75t_L g2831 ( 
.A(n_2716),
.B(n_1288),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2770),
.B(n_1293),
.Y(n_2832)
);

OAI21xp33_ASAP7_75t_L g2833 ( 
.A1(n_2735),
.A2(n_1306),
.B(n_1296),
.Y(n_2833)
);

OAI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2639),
.A2(n_2527),
.B(n_2339),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2607),
.B(n_2555),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2622),
.B(n_2421),
.Y(n_2836)
);

OAI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2639),
.A2(n_2339),
.B(n_2565),
.Y(n_2837)
);

OAI21xp5_ASAP7_75t_L g2838 ( 
.A1(n_2641),
.A2(n_2591),
.B(n_2593),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2602),
.Y(n_2839)
);

NAND2x1_ASAP7_75t_L g2840 ( 
.A(n_2774),
.B(n_2235),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2607),
.B(n_2563),
.Y(n_2841)
);

NAND2xp33_ASAP7_75t_L g2842 ( 
.A(n_2735),
.B(n_2243),
.Y(n_2842)
);

AOI21xp5_ASAP7_75t_L g2843 ( 
.A1(n_2715),
.A2(n_2558),
.B(n_2550),
.Y(n_2843)
);

AOI21xp5_ASAP7_75t_L g2844 ( 
.A1(n_2720),
.A2(n_2558),
.B(n_2542),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2603),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_2688),
.B(n_1306),
.Y(n_2846)
);

AOI21xp5_ASAP7_75t_L g2847 ( 
.A1(n_2720),
.A2(n_2542),
.B(n_2541),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2623),
.Y(n_2848)
);

OAI21xp5_ASAP7_75t_L g2849 ( 
.A1(n_2641),
.A2(n_2710),
.B(n_2792),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2625),
.Y(n_2850)
);

AOI21x1_ASAP7_75t_L g2851 ( 
.A1(n_2748),
.A2(n_2541),
.B(n_2560),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2633),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2627),
.B(n_2631),
.Y(n_2853)
);

AOI22xp5_ASAP7_75t_L g2854 ( 
.A1(n_2737),
.A2(n_1314),
.B1(n_2214),
.B2(n_2411),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2668),
.A2(n_2560),
.B(n_2252),
.Y(n_2855)
);

NOR2xp67_ASAP7_75t_L g2856 ( 
.A(n_2620),
.B(n_2574),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2610),
.B(n_2474),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2608),
.Y(n_2858)
);

NOR2xp33_ASAP7_75t_L g2859 ( 
.A(n_2662),
.B(n_1314),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2755),
.B(n_2474),
.Y(n_2860)
);

AOI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2717),
.A2(n_2256),
.B(n_2247),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2658),
.B(n_2572),
.Y(n_2862)
);

AOI21xp5_ASAP7_75t_L g2863 ( 
.A1(n_2717),
.A2(n_2275),
.B(n_2267),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2613),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2659),
.B(n_2579),
.Y(n_2865)
);

OAI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2599),
.A2(n_2081),
.B1(n_2266),
.B2(n_2205),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2621),
.B(n_2635),
.Y(n_2867)
);

AOI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2640),
.A2(n_2745),
.B(n_2654),
.Y(n_2868)
);

AOI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_2725),
.A2(n_2582),
.B(n_2578),
.Y(n_2869)
);

INVx4_ASAP7_75t_L g2870 ( 
.A(n_2684),
.Y(n_2870)
);

NOR2xp33_ASAP7_75t_L g2871 ( 
.A(n_2647),
.B(n_1687),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2673),
.B(n_2593),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2677),
.B(n_2596),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2629),
.Y(n_2874)
);

BUFx4f_ASAP7_75t_L g2875 ( 
.A(n_2684),
.Y(n_2875)
);

OAI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_2710),
.A2(n_2596),
.B(n_1959),
.Y(n_2876)
);

BUFx3_ASAP7_75t_L g2877 ( 
.A(n_2601),
.Y(n_2877)
);

NOR2xp67_ASAP7_75t_SL g2878 ( 
.A(n_2606),
.B(n_2266),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2732),
.A2(n_2582),
.B(n_2578),
.Y(n_2879)
);

AOI21xp5_ASAP7_75t_L g2880 ( 
.A1(n_2734),
.A2(n_2589),
.B(n_2586),
.Y(n_2880)
);

O2A1O1Ixp5_ASAP7_75t_L g2881 ( 
.A1(n_2740),
.A2(n_2319),
.B(n_1959),
.C(n_2392),
.Y(n_2881)
);

A2O1A1Ixp33_ASAP7_75t_L g2882 ( 
.A1(n_2599),
.A2(n_2551),
.B(n_2552),
.C(n_2545),
.Y(n_2882)
);

HB1xp67_ASAP7_75t_L g2883 ( 
.A(n_2729),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2637),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2615),
.B(n_2564),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2776),
.B(n_2566),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_L g2887 ( 
.A(n_2656),
.B(n_2581),
.Y(n_2887)
);

O2A1O1Ixp5_ASAP7_75t_L g2888 ( 
.A1(n_2616),
.A2(n_2580),
.B(n_2586),
.C(n_2589),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_SL g2889 ( 
.A(n_2648),
.B(n_1461),
.Y(n_2889)
);

AOI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2760),
.A2(n_2214),
.B1(n_1470),
.B2(n_1461),
.Y(n_2890)
);

INVx11_ASAP7_75t_L g2891 ( 
.A(n_2741),
.Y(n_2891)
);

AOI21xp5_ASAP7_75t_L g2892 ( 
.A1(n_2777),
.A2(n_2193),
.B(n_2181),
.Y(n_2892)
);

AOI21xp5_ASAP7_75t_L g2893 ( 
.A1(n_2711),
.A2(n_2193),
.B(n_2181),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2722),
.A2(n_2347),
.B(n_2285),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2642),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2776),
.B(n_2089),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2646),
.Y(n_2897)
);

OAI21xp33_ASAP7_75t_L g2898 ( 
.A1(n_2638),
.A2(n_821),
.B(n_819),
.Y(n_2898)
);

NOR2xp67_ASAP7_75t_L g2899 ( 
.A(n_2653),
.B(n_2272),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2723),
.B(n_981),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2703),
.B(n_1470),
.Y(n_2901)
);

BUFx6f_ASAP7_75t_L g2902 ( 
.A(n_2782),
.Y(n_2902)
);

BUFx12f_ASAP7_75t_L g2903 ( 
.A(n_2741),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_2764),
.B(n_2784),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2759),
.B(n_2155),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2742),
.B(n_2165),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2742),
.B(n_2170),
.Y(n_2907)
);

AO21x1_ASAP7_75t_L g2908 ( 
.A1(n_2686),
.A2(n_2340),
.B(n_1778),
.Y(n_2908)
);

AOI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2690),
.A2(n_2285),
.B(n_2235),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2630),
.Y(n_2910)
);

BUFx8_ASAP7_75t_L g2911 ( 
.A(n_2794),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2775),
.B(n_2729),
.Y(n_2912)
);

AOI21xp5_ASAP7_75t_L g2913 ( 
.A1(n_2698),
.A2(n_2335),
.B(n_2120),
.Y(n_2913)
);

OAI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2609),
.A2(n_1649),
.B(n_2243),
.Y(n_2914)
);

INVxp67_ASAP7_75t_L g2915 ( 
.A(n_2738),
.Y(n_2915)
);

OAI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2609),
.A2(n_2756),
.B(n_2666),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2657),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2632),
.Y(n_2918)
);

AOI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2736),
.A2(n_2335),
.B(n_2120),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2775),
.B(n_2173),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2743),
.A2(n_2120),
.B(n_2097),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2663),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2757),
.B(n_2179),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2758),
.B(n_2184),
.Y(n_2924)
);

OAI21xp5_ASAP7_75t_L g2925 ( 
.A1(n_2756),
.A2(n_2264),
.B(n_2243),
.Y(n_2925)
);

AND2x4_ASAP7_75t_L g2926 ( 
.A(n_2755),
.B(n_2183),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2755),
.B(n_2183),
.Y(n_2927)
);

OAI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2666),
.A2(n_2264),
.B(n_2243),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2634),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_L g2930 ( 
.A(n_2674),
.B(n_2208),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2767),
.B(n_2189),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2644),
.Y(n_2932)
);

AOI21xp5_ASAP7_75t_L g2933 ( 
.A1(n_2781),
.A2(n_2168),
.B(n_2120),
.Y(n_2933)
);

AOI21xp5_ASAP7_75t_L g2934 ( 
.A1(n_2785),
.A2(n_2768),
.B(n_2763),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2669),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2612),
.B(n_2195),
.Y(n_2936)
);

AOI21xp5_ASAP7_75t_L g2937 ( 
.A1(n_2766),
.A2(n_2174),
.B(n_2168),
.Y(n_2937)
);

A2O1A1Ixp33_ASAP7_75t_L g2938 ( 
.A1(n_2680),
.A2(n_1613),
.B(n_2272),
.C(n_2158),
.Y(n_2938)
);

OAI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2680),
.A2(n_2687),
.B1(n_2739),
.B2(n_2652),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2671),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2651),
.Y(n_2941)
);

BUFx6f_ASAP7_75t_L g2942 ( 
.A(n_2783),
.Y(n_2942)
);

AOI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2772),
.A2(n_2174),
.B(n_2168),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_SL g2944 ( 
.A(n_2650),
.B(n_2356),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2672),
.Y(n_2945)
);

INVx3_ASAP7_75t_L g2946 ( 
.A(n_2765),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_SL g2947 ( 
.A(n_2675),
.B(n_2356),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2762),
.B(n_2197),
.Y(n_2948)
);

INVx4_ASAP7_75t_L g2949 ( 
.A(n_2765),
.Y(n_2949)
);

BUFx2_ASAP7_75t_L g2950 ( 
.A(n_2783),
.Y(n_2950)
);

AOI21xp5_ASAP7_75t_L g2951 ( 
.A1(n_2787),
.A2(n_2174),
.B(n_2168),
.Y(n_2951)
);

HB1xp67_ASAP7_75t_L g2952 ( 
.A(n_2655),
.Y(n_2952)
);

AND2x4_ASAP7_75t_L g2953 ( 
.A(n_2733),
.B(n_2378),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2682),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_2791),
.B(n_2356),
.Y(n_2955)
);

A2O1A1Ixp33_ASAP7_75t_L g2956 ( 
.A1(n_2624),
.A2(n_1613),
.B(n_2158),
.C(n_2148),
.Y(n_2956)
);

AOI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2652),
.A2(n_2773),
.B(n_2747),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2664),
.B(n_2251),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2676),
.Y(n_2959)
);

INVx3_ASAP7_75t_L g2960 ( 
.A(n_2611),
.Y(n_2960)
);

AOI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2747),
.A2(n_2211),
.B(n_2174),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2636),
.B(n_2292),
.Y(n_2962)
);

AOI21xp5_ASAP7_75t_L g2963 ( 
.A1(n_2773),
.A2(n_2325),
.B(n_2211),
.Y(n_2963)
);

AO21x1_ASAP7_75t_L g2964 ( 
.A1(n_2753),
.A2(n_2340),
.B(n_1778),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2704),
.Y(n_2965)
);

AOI21xp5_ASAP7_75t_L g2966 ( 
.A1(n_2780),
.A2(n_2769),
.B(n_2786),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2678),
.B(n_2296),
.Y(n_2967)
);

AOI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2670),
.A2(n_2385),
.B1(n_768),
.B2(n_769),
.Y(n_2968)
);

NOR2xp33_ASAP7_75t_L g2969 ( 
.A(n_2778),
.B(n_2291),
.Y(n_2969)
);

OAI321xp33_ASAP7_75t_L g2970 ( 
.A1(n_2687),
.A2(n_983),
.A3(n_982),
.B1(n_1009),
.B2(n_1078),
.C(n_1073),
.Y(n_2970)
);

NOR2x1_ASAP7_75t_L g2971 ( 
.A(n_2719),
.B(n_2554),
.Y(n_2971)
);

OAI21xp33_ASAP7_75t_L g2972 ( 
.A1(n_2780),
.A2(n_711),
.B(n_710),
.Y(n_2972)
);

OAI22xp5_ASAP7_75t_L g2973 ( 
.A1(n_2786),
.A2(n_2681),
.B1(n_2689),
.B2(n_2679),
.Y(n_2973)
);

OAI21xp5_ASAP7_75t_L g2974 ( 
.A1(n_2769),
.A2(n_2264),
.B(n_2299),
.Y(n_2974)
);

HB1xp67_ASAP7_75t_L g2975 ( 
.A(n_2691),
.Y(n_2975)
);

INVx6_ASAP7_75t_L g2976 ( 
.A(n_2731),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2697),
.B(n_2304),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2702),
.B(n_2306),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2724),
.B(n_2307),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2744),
.B(n_2318),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2693),
.B(n_2320),
.Y(n_2981)
);

AOI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2730),
.A2(n_2325),
.B(n_2211),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2694),
.B(n_2328),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2696),
.B(n_2329),
.Y(n_2984)
);

AOI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2751),
.A2(n_2325),
.B(n_2211),
.Y(n_2985)
);

AOI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2754),
.A2(n_2325),
.B(n_1770),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2699),
.Y(n_2987)
);

BUFx6f_ASAP7_75t_L g2988 ( 
.A(n_2902),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2857),
.B(n_2915),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_2904),
.B(n_2900),
.Y(n_2990)
);

HB1xp67_ASAP7_75t_L g2991 ( 
.A(n_2883),
.Y(n_2991)
);

INVx6_ASAP7_75t_L g2992 ( 
.A(n_2911),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2839),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2848),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2821),
.B(n_2707),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2952),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_SL g2997 ( 
.A(n_2819),
.B(n_2726),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2975),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_L g2999 ( 
.A1(n_2833),
.A2(n_2793),
.B1(n_2264),
.B2(n_2779),
.Y(n_2999)
);

OR2x6_ASAP7_75t_L g3000 ( 
.A(n_2966),
.B(n_2957),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2853),
.B(n_2790),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2867),
.B(n_2790),
.Y(n_3002)
);

HB1xp67_ASAP7_75t_L g3003 ( 
.A(n_2912),
.Y(n_3003)
);

BUFx2_ASAP7_75t_L g3004 ( 
.A(n_2860),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2809),
.Y(n_3005)
);

BUFx6f_ASAP7_75t_L g3006 ( 
.A(n_2902),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2849),
.B(n_2790),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2868),
.B(n_2790),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2820),
.Y(n_3009)
);

INVx3_ASAP7_75t_L g3010 ( 
.A(n_2942),
.Y(n_3010)
);

AND2x2_ASAP7_75t_L g3011 ( 
.A(n_2860),
.B(n_2705),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2845),
.Y(n_3012)
);

INVxp67_ASAP7_75t_L g3013 ( 
.A(n_2832),
.Y(n_3013)
);

INVx3_ASAP7_75t_L g3014 ( 
.A(n_2942),
.Y(n_3014)
);

BUFx3_ASAP7_75t_L g3015 ( 
.A(n_2902),
.Y(n_3015)
);

INVx1_ASAP7_75t_SL g3016 ( 
.A(n_2950),
.Y(n_3016)
);

INVx3_ASAP7_75t_L g3017 ( 
.A(n_2942),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2858),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2864),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2811),
.B(n_2816),
.Y(n_3020)
);

BUFx2_ASAP7_75t_L g3021 ( 
.A(n_2926),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2836),
.B(n_2706),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2874),
.Y(n_3023)
);

BUFx2_ASAP7_75t_L g3024 ( 
.A(n_2926),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2796),
.B(n_2708),
.Y(n_3025)
);

OAI22xp5_ASAP7_75t_L g3026 ( 
.A1(n_2833),
.A2(n_721),
.B1(n_723),
.B2(n_717),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2797),
.B(n_2790),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2910),
.Y(n_3028)
);

CKINVDCx5p33_ASAP7_75t_R g3029 ( 
.A(n_2903),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2830),
.B(n_2712),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2836),
.B(n_2718),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2905),
.B(n_2721),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2799),
.B(n_2519),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2850),
.Y(n_3034)
);

NOR2xp33_ASAP7_75t_L g3035 ( 
.A(n_2805),
.B(n_2727),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2862),
.B(n_2728),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2852),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2918),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2929),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2932),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2872),
.B(n_2790),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_SL g3042 ( 
.A(n_2808),
.B(n_2746),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2873),
.B(n_2749),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2941),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_SL g3045 ( 
.A(n_2803),
.B(n_2750),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2877),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_2887),
.B(n_2788),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_SL g3048 ( 
.A(n_2802),
.B(n_2939),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2934),
.B(n_2789),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2973),
.B(n_2774),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2959),
.Y(n_3051)
);

BUFx6f_ASAP7_75t_L g3052 ( 
.A(n_2875),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2798),
.B(n_1079),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2813),
.B(n_622),
.Y(n_3054)
);

AND2x2_ASAP7_75t_SL g3055 ( 
.A(n_2842),
.B(n_2381),
.Y(n_3055)
);

AND3x1_ASAP7_75t_L g3056 ( 
.A(n_2901),
.B(n_2968),
.C(n_2854),
.Y(n_3056)
);

BUFx3_ASAP7_75t_L g3057 ( 
.A(n_2911),
.Y(n_3057)
);

INVx4_ASAP7_75t_L g3058 ( 
.A(n_2801),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2802),
.B(n_2774),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2886),
.Y(n_3060)
);

OAI21x1_ASAP7_75t_L g3061 ( 
.A1(n_2844),
.A2(n_1793),
.B(n_1791),
.Y(n_3061)
);

AND3x1_ASAP7_75t_SL g3062 ( 
.A(n_2968),
.B(n_723),
.C(n_721),
.Y(n_3062)
);

BUFx4f_ASAP7_75t_L g3063 ( 
.A(n_2965),
.Y(n_3063)
);

HB1xp67_ASAP7_75t_L g3064 ( 
.A(n_2835),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2841),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_SL g3066 ( 
.A(n_2854),
.B(n_2356),
.Y(n_3066)
);

INVx3_ASAP7_75t_L g3067 ( 
.A(n_2875),
.Y(n_3067)
);

INVx2_ASAP7_75t_SL g3068 ( 
.A(n_2891),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2838),
.B(n_2356),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2884),
.Y(n_3070)
);

NOR2xp33_ASAP7_75t_L g3071 ( 
.A(n_2846),
.B(n_698),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2895),
.Y(n_3072)
);

OR2x2_ASAP7_75t_L g3073 ( 
.A(n_2885),
.B(n_2329),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2967),
.B(n_698),
.Y(n_3074)
);

AND2x4_ASAP7_75t_L g3075 ( 
.A(n_2812),
.B(n_2381),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_L g3076 ( 
.A(n_2831),
.B(n_699),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2865),
.B(n_2774),
.Y(n_3077)
);

CKINVDCx5p33_ASAP7_75t_R g3078 ( 
.A(n_2965),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2936),
.B(n_2958),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2906),
.B(n_2774),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_2897),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2896),
.B(n_764),
.Y(n_3082)
);

CKINVDCx20_ASAP7_75t_R g3083 ( 
.A(n_2976),
.Y(n_3083)
);

INVx4_ASAP7_75t_L g3084 ( 
.A(n_2801),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2917),
.Y(n_3085)
);

INVx3_ASAP7_75t_L g3086 ( 
.A(n_2812),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2922),
.B(n_772),
.Y(n_3087)
);

BUFx4f_ASAP7_75t_L g3088 ( 
.A(n_2965),
.Y(n_3088)
);

NOR2x1p5_ASAP7_75t_L g3089 ( 
.A(n_2870),
.B(n_699),
.Y(n_3089)
);

BUFx4f_ASAP7_75t_L g3090 ( 
.A(n_2976),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2935),
.B(n_2334),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2940),
.Y(n_3092)
);

CKINVDCx5p33_ASAP7_75t_R g3093 ( 
.A(n_2930),
.Y(n_3093)
);

HB1xp67_ASAP7_75t_L g3094 ( 
.A(n_2907),
.Y(n_3094)
);

AND2x4_ASAP7_75t_L g3095 ( 
.A(n_2870),
.B(n_2381),
.Y(n_3095)
);

INVx3_ASAP7_75t_L g3096 ( 
.A(n_2927),
.Y(n_3096)
);

A2O1A1Ixp33_ASAP7_75t_L g3097 ( 
.A1(n_2972),
.A2(n_703),
.B(n_709),
.C(n_702),
.Y(n_3097)
);

INVxp67_ASAP7_75t_L g3098 ( 
.A(n_2859),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2945),
.Y(n_3099)
);

INVx4_ASAP7_75t_L g3100 ( 
.A(n_2795),
.Y(n_3100)
);

INVx1_ASAP7_75t_SL g3101 ( 
.A(n_2920),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2916),
.B(n_2334),
.Y(n_3102)
);

BUFx6f_ASAP7_75t_L g3103 ( 
.A(n_2810),
.Y(n_3103)
);

AND2x2_ASAP7_75t_L g3104 ( 
.A(n_2954),
.B(n_702),
.Y(n_3104)
);

INVxp33_ASAP7_75t_L g3105 ( 
.A(n_2969),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_L g3106 ( 
.A(n_2825),
.B(n_703),
.Y(n_3106)
);

NOR2x1_ASAP7_75t_L g3107 ( 
.A(n_2826),
.B(n_2148),
.Y(n_3107)
);

BUFx3_ASAP7_75t_L g3108 ( 
.A(n_2810),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2931),
.B(n_2336),
.Y(n_3109)
);

NOR2xp33_ASAP7_75t_L g3110 ( 
.A(n_2825),
.B(n_709),
.Y(n_3110)
);

BUFx6f_ASAP7_75t_L g3111 ( 
.A(n_2927),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2923),
.B(n_2336),
.Y(n_3112)
);

INVx2_ASAP7_75t_SL g3113 ( 
.A(n_2953),
.Y(n_3113)
);

CKINVDCx20_ASAP7_75t_R g3114 ( 
.A(n_2814),
.Y(n_3114)
);

AOI221x1_ASAP7_75t_L g3115 ( 
.A1(n_2938),
.A2(n_2405),
.B1(n_2517),
.B2(n_2390),
.C(n_2383),
.Y(n_3115)
);

BUFx6f_ASAP7_75t_L g3116 ( 
.A(n_2953),
.Y(n_3116)
);

INVx1_ASAP7_75t_SL g3117 ( 
.A(n_2962),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2987),
.B(n_713),
.Y(n_3118)
);

INVx2_ASAP7_75t_SL g3119 ( 
.A(n_2946),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2977),
.Y(n_3120)
);

BUFx6f_ASAP7_75t_L g3121 ( 
.A(n_2946),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2823),
.B(n_728),
.Y(n_3122)
);

INVx3_ASAP7_75t_L g3123 ( 
.A(n_2795),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2924),
.B(n_728),
.Y(n_3124)
);

HB1xp67_ASAP7_75t_L g3125 ( 
.A(n_2948),
.Y(n_3125)
);

BUFx3_ASAP7_75t_L g3126 ( 
.A(n_2949),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2978),
.B(n_731),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2979),
.B(n_731),
.Y(n_3128)
);

OR2x2_ASAP7_75t_L g3129 ( 
.A(n_2944),
.B(n_2947),
.Y(n_3129)
);

AO22x1_ASAP7_75t_L g3130 ( 
.A1(n_2971),
.A2(n_774),
.B1(n_781),
.B2(n_773),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2980),
.B(n_773),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2878),
.B(n_774),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2981),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2983),
.Y(n_3134)
);

HB1xp67_ASAP7_75t_L g3135 ( 
.A(n_2955),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2869),
.B(n_2264),
.Y(n_3136)
);

BUFx6f_ASAP7_75t_L g3137 ( 
.A(n_2949),
.Y(n_3137)
);

AOI221xp5_ASAP7_75t_L g3138 ( 
.A1(n_2898),
.A2(n_784),
.B1(n_783),
.B2(n_781),
.C(n_1009),
.Y(n_3138)
);

INVx3_ASAP7_75t_L g3139 ( 
.A(n_2960),
.Y(n_3139)
);

CKINVDCx20_ASAP7_75t_R g3140 ( 
.A(n_2889),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2879),
.B(n_2452),
.Y(n_3141)
);

AND3x1_ASAP7_75t_SL g3142 ( 
.A(n_2866),
.B(n_783),
.C(n_5),
.Y(n_3142)
);

BUFx3_ASAP7_75t_L g3143 ( 
.A(n_2871),
.Y(n_3143)
);

INVx5_ASAP7_75t_L g3144 ( 
.A(n_2960),
.Y(n_3144)
);

NOR2xp33_ASAP7_75t_L g3145 ( 
.A(n_2890),
.B(n_2856),
.Y(n_3145)
);

INVx2_ASAP7_75t_SL g3146 ( 
.A(n_2984),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2851),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2817),
.Y(n_3148)
);

AND2x4_ASAP7_75t_L g3149 ( 
.A(n_2899),
.B(n_2383),
.Y(n_3149)
);

AO22x1_ASAP7_75t_L g3150 ( 
.A1(n_2837),
.A2(n_714),
.B1(n_715),
.B2(n_713),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2824),
.B(n_714),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2888),
.Y(n_3152)
);

INVx1_ASAP7_75t_SL g3153 ( 
.A(n_2933),
.Y(n_3153)
);

BUFx4f_ASAP7_75t_L g3154 ( 
.A(n_2964),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2840),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2881),
.Y(n_3156)
);

NAND3xp33_ASAP7_75t_L g3157 ( 
.A(n_2834),
.B(n_720),
.C(n_715),
.Y(n_3157)
);

CKINVDCx5p33_ASAP7_75t_R g3158 ( 
.A(n_2951),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2876),
.Y(n_3159)
);

OAI22xp5_ASAP7_75t_L g3160 ( 
.A1(n_2882),
.A2(n_2390),
.B1(n_2405),
.B2(n_2383),
.Y(n_3160)
);

BUFx6f_ASAP7_75t_L g3161 ( 
.A(n_2961),
.Y(n_3161)
);

INVx3_ASAP7_75t_L g3162 ( 
.A(n_2985),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_SL g3163 ( 
.A(n_2829),
.B(n_2452),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2855),
.B(n_720),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2880),
.B(n_2807),
.Y(n_3165)
);

CKINVDCx5p33_ASAP7_75t_R g3166 ( 
.A(n_2919),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2974),
.Y(n_3167)
);

BUFx3_ASAP7_75t_L g3168 ( 
.A(n_2908),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2828),
.B(n_2452),
.Y(n_3169)
);

AND2x4_ASAP7_75t_L g3170 ( 
.A(n_2943),
.B(n_2390),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_2892),
.B(n_2452),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_SL g3172 ( 
.A(n_2893),
.B(n_2452),
.Y(n_3172)
);

INVx3_ASAP7_75t_L g3173 ( 
.A(n_2937),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2843),
.B(n_2847),
.Y(n_3174)
);

OR2x6_ASAP7_75t_L g3175 ( 
.A(n_2815),
.B(n_2405),
.Y(n_3175)
);

INVx3_ASAP7_75t_L g3176 ( 
.A(n_2921),
.Y(n_3176)
);

AND2x2_ASAP7_75t_L g3177 ( 
.A(n_2956),
.B(n_729),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_2970),
.B(n_729),
.Y(n_3178)
);

BUFx2_ASAP7_75t_L g3179 ( 
.A(n_2928),
.Y(n_3179)
);

HB1xp67_ASAP7_75t_L g3180 ( 
.A(n_2963),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2925),
.Y(n_3181)
);

INVx3_ASAP7_75t_L g3182 ( 
.A(n_2913),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2861),
.B(n_732),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2827),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2822),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_SL g3186 ( 
.A(n_2909),
.B(n_2517),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2806),
.Y(n_3187)
);

INVx2_ASAP7_75t_SL g3188 ( 
.A(n_2986),
.Y(n_3188)
);

INVx2_ASAP7_75t_SL g3189 ( 
.A(n_2800),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2996),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_3105),
.B(n_732),
.Y(n_3191)
);

BUFx12f_ASAP7_75t_L g3192 ( 
.A(n_3078),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_3098),
.B(n_775),
.Y(n_3193)
);

AOI21xp33_ASAP7_75t_L g3194 ( 
.A1(n_3157),
.A2(n_2914),
.B(n_2818),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2998),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_3013),
.B(n_775),
.Y(n_3196)
);

BUFx6f_ASAP7_75t_L g3197 ( 
.A(n_2988),
.Y(n_3197)
);

BUFx3_ASAP7_75t_L g3198 ( 
.A(n_3015),
.Y(n_3198)
);

HB1xp67_ASAP7_75t_L g3199 ( 
.A(n_2991),
.Y(n_3199)
);

BUFx6f_ASAP7_75t_L g3200 ( 
.A(n_2988),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_3165),
.A2(n_2863),
.B(n_2804),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3005),
.Y(n_3202)
);

BUFx6f_ASAP7_75t_L g3203 ( 
.A(n_2988),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_3003),
.B(n_3094),
.Y(n_3204)
);

AOI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_3174),
.A2(n_2982),
.B(n_2894),
.Y(n_3205)
);

NOR2xp33_ASAP7_75t_L g3206 ( 
.A(n_3093),
.B(n_5),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3101),
.B(n_6),
.Y(n_3207)
);

BUFx6f_ASAP7_75t_L g3208 ( 
.A(n_3006),
.Y(n_3208)
);

AOI22xp5_ASAP7_75t_L g3209 ( 
.A1(n_3056),
.A2(n_2268),
.B1(n_1603),
.B2(n_2175),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3009),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_3174),
.A2(n_1830),
.B(n_1826),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3012),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3018),
.Y(n_3213)
);

AOI21xp5_ASAP7_75t_L g3214 ( 
.A1(n_3008),
.A2(n_3048),
.B(n_3150),
.Y(n_3214)
);

NOR2x1_ASAP7_75t_SL g3215 ( 
.A(n_3000),
.B(n_2517),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_R g3216 ( 
.A(n_3029),
.B(n_2562),
.Y(n_3216)
);

AND2x4_ASAP7_75t_L g3217 ( 
.A(n_3019),
.B(n_2562),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_3101),
.B(n_7),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3023),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_3028),
.Y(n_3220)
);

OR2x2_ASAP7_75t_L g3221 ( 
.A(n_3000),
.B(n_1132),
.Y(n_3221)
);

BUFx6f_ASAP7_75t_L g3222 ( 
.A(n_3006),
.Y(n_3222)
);

HB1xp67_ASAP7_75t_L g3223 ( 
.A(n_3135),
.Y(n_3223)
);

CKINVDCx20_ASAP7_75t_R g3224 ( 
.A(n_3083),
.Y(n_3224)
);

BUFx4f_ASAP7_75t_SL g3225 ( 
.A(n_3057),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_3020),
.B(n_9),
.Y(n_3226)
);

CKINVDCx5p33_ASAP7_75t_R g3227 ( 
.A(n_3090),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_3038),
.Y(n_3228)
);

BUFx6f_ASAP7_75t_L g3229 ( 
.A(n_3006),
.Y(n_3229)
);

BUFx8_ASAP7_75t_L g3230 ( 
.A(n_3068),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_3064),
.B(n_11),
.Y(n_3231)
);

CKINVDCx5p33_ASAP7_75t_R g3232 ( 
.A(n_3090),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3117),
.B(n_11),
.Y(n_3233)
);

HB1xp67_ASAP7_75t_L g3234 ( 
.A(n_3125),
.Y(n_3234)
);

NOR2xp33_ASAP7_75t_L g3235 ( 
.A(n_2997),
.B(n_12),
.Y(n_3235)
);

NAND2x1_ASAP7_75t_L g3236 ( 
.A(n_3139),
.B(n_2562),
.Y(n_3236)
);

INVx4_ASAP7_75t_L g3237 ( 
.A(n_3137),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_3039),
.Y(n_3238)
);

O2A1O1Ixp33_ASAP7_75t_L g3239 ( 
.A1(n_3106),
.A2(n_2175),
.B(n_2177),
.C(n_2164),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_3117),
.B(n_12),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_3143),
.B(n_13),
.Y(n_3241)
);

HB1xp67_ASAP7_75t_L g3242 ( 
.A(n_3016),
.Y(n_3242)
);

OAI222xp33_ASAP7_75t_SL g3243 ( 
.A1(n_3056),
.A2(n_3100),
.B1(n_3058),
.B2(n_3084),
.C1(n_3088),
.C2(n_3063),
.Y(n_3243)
);

A2O1A1Ixp33_ASAP7_75t_L g3244 ( 
.A1(n_3157),
.A2(n_2164),
.B(n_2212),
.C(n_2177),
.Y(n_3244)
);

BUFx4f_ASAP7_75t_L g3245 ( 
.A(n_3052),
.Y(n_3245)
);

O2A1O1Ixp33_ASAP7_75t_L g3246 ( 
.A1(n_3110),
.A2(n_2218),
.B(n_2240),
.C(n_2212),
.Y(n_3246)
);

INVx1_ASAP7_75t_SL g3247 ( 
.A(n_3047),
.Y(n_3247)
);

INVx4_ASAP7_75t_L g3248 ( 
.A(n_3137),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_3008),
.A2(n_1830),
.B(n_1826),
.Y(n_3249)
);

NAND2x1p5_ASAP7_75t_L g3250 ( 
.A(n_3144),
.B(n_2338),
.Y(n_3250)
);

INVx1_ASAP7_75t_SL g3251 ( 
.A(n_2989),
.Y(n_3251)
);

BUFx12f_ASAP7_75t_L g3252 ( 
.A(n_3046),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_3040),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_3004),
.B(n_13),
.Y(n_3254)
);

AND2x4_ASAP7_75t_L g3255 ( 
.A(n_3044),
.B(n_2218),
.Y(n_3255)
);

A2O1A1Ixp33_ASAP7_75t_SL g3256 ( 
.A1(n_3145),
.A2(n_1141),
.B(n_1475),
.C(n_1469),
.Y(n_3256)
);

HAxp5_ASAP7_75t_L g3257 ( 
.A(n_3089),
.B(n_14),
.CON(n_3257),
.SN(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3051),
.Y(n_3258)
);

OR2x2_ASAP7_75t_L g3259 ( 
.A(n_3000),
.B(n_1141),
.Y(n_3259)
);

INVx3_ASAP7_75t_L g3260 ( 
.A(n_3121),
.Y(n_3260)
);

O2A1O1Ixp33_ASAP7_75t_L g3261 ( 
.A1(n_3026),
.A2(n_2338),
.B(n_2240),
.C(n_1922),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_3060),
.B(n_15),
.Y(n_3262)
);

NOR2xp33_ASAP7_75t_L g3263 ( 
.A(n_3035),
.B(n_15),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_3070),
.Y(n_3264)
);

INVx2_ASAP7_75t_SL g3265 ( 
.A(n_3046),
.Y(n_3265)
);

OAI22xp5_ASAP7_75t_L g3266 ( 
.A1(n_3114),
.A2(n_1825),
.B1(n_1840),
.B2(n_1769),
.Y(n_3266)
);

BUFx6f_ASAP7_75t_L g3267 ( 
.A(n_3046),
.Y(n_3267)
);

INVx3_ASAP7_75t_L g3268 ( 
.A(n_3121),
.Y(n_3268)
);

BUFx2_ASAP7_75t_L g3269 ( 
.A(n_3021),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3065),
.B(n_16),
.Y(n_3270)
);

BUFx3_ASAP7_75t_L g3271 ( 
.A(n_2992),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_3072),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3141),
.A2(n_1830),
.B(n_1826),
.Y(n_3273)
);

AOI22xp33_ASAP7_75t_L g3274 ( 
.A1(n_3066),
.A2(n_1603),
.B1(n_1842),
.B2(n_1830),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3085),
.Y(n_3275)
);

INVx3_ASAP7_75t_L g3276 ( 
.A(n_3121),
.Y(n_3276)
);

AOI22xp33_ASAP7_75t_L g3277 ( 
.A1(n_3179),
.A2(n_1603),
.B1(n_1902),
.B2(n_1842),
.Y(n_3277)
);

AND3x1_ASAP7_75t_SL g3278 ( 
.A(n_3138),
.B(n_3142),
.C(n_3062),
.Y(n_3278)
);

BUFx3_ASAP7_75t_L g3279 ( 
.A(n_2992),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3092),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3099),
.Y(n_3281)
);

INVx2_ASAP7_75t_SL g3282 ( 
.A(n_3063),
.Y(n_3282)
);

O2A1O1Ixp33_ASAP7_75t_L g3283 ( 
.A1(n_3026),
.A2(n_1922),
.B(n_1972),
.C(n_1915),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3079),
.B(n_17),
.Y(n_3284)
);

BUFx2_ASAP7_75t_L g3285 ( 
.A(n_3024),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3152),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2993),
.Y(n_3287)
);

O2A1O1Ixp33_ASAP7_75t_SL g3288 ( 
.A1(n_3045),
.A2(n_21),
.B(n_18),
.C(n_19),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_3141),
.A2(n_1902),
.B(n_1842),
.Y(n_3289)
);

INVx3_ASAP7_75t_L g3290 ( 
.A(n_3096),
.Y(n_3290)
);

INVx3_ASAP7_75t_L g3291 ( 
.A(n_3096),
.Y(n_3291)
);

AOI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_3164),
.A2(n_1902),
.B(n_1842),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_2994),
.Y(n_3293)
);

AO22x1_ASAP7_75t_L g3294 ( 
.A1(n_3166),
.A2(n_23),
.B1(n_18),
.B2(n_21),
.Y(n_3294)
);

OR2x6_ASAP7_75t_L g3295 ( 
.A(n_3058),
.B(n_1902),
.Y(n_3295)
);

A2O1A1Ixp33_ASAP7_75t_L g3296 ( 
.A1(n_3054),
.A2(n_1791),
.B(n_1793),
.C(n_1839),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3147),
.Y(n_3297)
);

O2A1O1Ixp5_ASAP7_75t_L g3298 ( 
.A1(n_3154),
.A2(n_3027),
.B(n_3163),
.C(n_3069),
.Y(n_3298)
);

BUFx12f_ASAP7_75t_L g3299 ( 
.A(n_3052),
.Y(n_3299)
);

NOR2xp33_ASAP7_75t_L g3300 ( 
.A(n_3071),
.B(n_23),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3007),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3007),
.Y(n_3302)
);

A2O1A1Ixp33_ASAP7_75t_L g3303 ( 
.A1(n_3076),
.A2(n_1839),
.B(n_1825),
.C(n_1769),
.Y(n_3303)
);

INVx3_ASAP7_75t_L g3304 ( 
.A(n_3111),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_3183),
.A2(n_1919),
.B(n_1917),
.Y(n_3305)
);

AOI21xp5_ASAP7_75t_L g3306 ( 
.A1(n_3171),
.A2(n_1919),
.B(n_1917),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3034),
.Y(n_3307)
);

INVx3_ASAP7_75t_L g3308 ( 
.A(n_3111),
.Y(n_3308)
);

OAI22xp5_ASAP7_75t_L g3309 ( 
.A1(n_2999),
.A2(n_1864),
.B1(n_1840),
.B2(n_1749),
.Y(n_3309)
);

OAI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_3140),
.A2(n_1864),
.B1(n_1755),
.B2(n_1917),
.Y(n_3310)
);

A2O1A1Ixp33_ASAP7_75t_L g3311 ( 
.A1(n_3154),
.A2(n_2038),
.B(n_1915),
.C(n_1979),
.Y(n_3311)
);

A2O1A1Ixp33_ASAP7_75t_L g3312 ( 
.A1(n_3178),
.A2(n_2038),
.B(n_1972),
.C(n_1994),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_2995),
.B(n_3120),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3002),
.B(n_24),
.Y(n_3314)
);

AOI222xp33_ASAP7_75t_L g3315 ( 
.A1(n_3130),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.C1(n_25),
.C2(n_28),
.Y(n_3315)
);

AND2x4_ASAP7_75t_L g3316 ( 
.A(n_3016),
.B(n_2268),
.Y(n_3316)
);

HB1xp67_ASAP7_75t_L g3317 ( 
.A(n_3129),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3002),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3172),
.A2(n_3169),
.B(n_3189),
.Y(n_3319)
);

OAI22x1_ASAP7_75t_L g3320 ( 
.A1(n_3159),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3049),
.Y(n_3321)
);

O2A1O1Ixp33_ASAP7_75t_L g3322 ( 
.A1(n_3097),
.A2(n_1994),
.B(n_2000),
.C(n_1979),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3037),
.Y(n_3323)
);

OAI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3055),
.A2(n_1755),
.B1(n_1919),
.B2(n_1917),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3081),
.Y(n_3325)
);

O2A1O1Ixp33_ASAP7_75t_L g3326 ( 
.A1(n_3132),
.A2(n_2030),
.B(n_2033),
.C(n_2000),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_2990),
.B(n_31),
.Y(n_3327)
);

OR2x6_ASAP7_75t_L g3328 ( 
.A(n_3084),
.B(n_1919),
.Y(n_3328)
);

INVx5_ASAP7_75t_L g3329 ( 
.A(n_3162),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3049),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3148),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3001),
.Y(n_3332)
);

NOR2xp33_ASAP7_75t_L g3333 ( 
.A(n_3033),
.B(n_32),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3001),
.B(n_33),
.Y(n_3334)
);

INVx2_ASAP7_75t_SL g3335 ( 
.A(n_3088),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_3169),
.A2(n_2268),
.B(n_2025),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_3022),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_3111),
.B(n_34),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3146),
.B(n_34),
.Y(n_3339)
);

HB1xp67_ASAP7_75t_L g3340 ( 
.A(n_3180),
.Y(n_3340)
);

NOR2xp33_ASAP7_75t_L g3341 ( 
.A(n_3108),
.B(n_35),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3041),
.Y(n_3342)
);

O2A1O1Ixp33_ASAP7_75t_L g3343 ( 
.A1(n_3042),
.A2(n_2033),
.B(n_2030),
.C(n_1579),
.Y(n_3343)
);

AOI221xp5_ASAP7_75t_L g3344 ( 
.A1(n_3122),
.A2(n_1585),
.B1(n_1591),
.B2(n_1579),
.C(n_1575),
.Y(n_3344)
);

A2O1A1Ixp33_ASAP7_75t_L g3345 ( 
.A1(n_3177),
.A2(n_2038),
.B(n_37),
.C(n_35),
.Y(n_3345)
);

A2O1A1Ixp33_ASAP7_75t_L g3346 ( 
.A1(n_3151),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_3346)
);

OAI22x1_ASAP7_75t_SL g3347 ( 
.A1(n_3158),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_3133),
.B(n_39),
.Y(n_3348)
);

NOR2xp33_ASAP7_75t_SL g3349 ( 
.A(n_3052),
.B(n_1966),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_3103),
.B(n_40),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3030),
.B(n_3032),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_SL g3352 ( 
.A(n_3067),
.B(n_1966),
.Y(n_3352)
);

A2O1A1Ixp33_ASAP7_75t_SL g3353 ( 
.A1(n_3182),
.A2(n_1475),
.B(n_1469),
.C(n_1583),
.Y(n_3353)
);

AND2x4_ASAP7_75t_L g3354 ( 
.A(n_3086),
.B(n_1585),
.Y(n_3354)
);

INVx6_ASAP7_75t_L g3355 ( 
.A(n_3116),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3041),
.B(n_41),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_3134),
.B(n_42),
.Y(n_3357)
);

OR2x2_ASAP7_75t_L g3358 ( 
.A(n_3187),
.B(n_1591),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3043),
.B(n_43),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3011),
.B(n_44),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3031),
.Y(n_3361)
);

AND2x6_ASAP7_75t_L g3362 ( 
.A(n_3059),
.B(n_1592),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3073),
.Y(n_3363)
);

INVx6_ASAP7_75t_L g3364 ( 
.A(n_3116),
.Y(n_3364)
);

O2A1O1Ixp33_ASAP7_75t_L g3365 ( 
.A1(n_3025),
.A2(n_1584),
.B(n_1583),
.C(n_1558),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3185),
.Y(n_3366)
);

AOI22xp33_ASAP7_75t_SL g3367 ( 
.A1(n_3059),
.A2(n_910),
.B1(n_866),
.B2(n_48),
.Y(n_3367)
);

O2A1O1Ixp5_ASAP7_75t_SL g3368 ( 
.A1(n_3173),
.A2(n_1770),
.B(n_1750),
.C(n_1584),
.Y(n_3368)
);

INVxp67_ASAP7_75t_L g3369 ( 
.A(n_3074),
.Y(n_3369)
);

HB1xp67_ASAP7_75t_L g3370 ( 
.A(n_3080),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3043),
.B(n_45),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3102),
.Y(n_3372)
);

BUFx6f_ASAP7_75t_L g3373 ( 
.A(n_3116),
.Y(n_3373)
);

A2O1A1Ixp33_ASAP7_75t_L g3374 ( 
.A1(n_3168),
.A2(n_3160),
.B(n_3050),
.C(n_3053),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3102),
.Y(n_3375)
);

AOI22xp33_ASAP7_75t_L g3376 ( 
.A1(n_3167),
.A2(n_1592),
.B1(n_1622),
.B2(n_1602),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3156),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_SL g3378 ( 
.A(n_3103),
.B(n_1592),
.Y(n_3378)
);

INVx3_ASAP7_75t_L g3379 ( 
.A(n_3137),
.Y(n_3379)
);

NAND3xp33_ASAP7_75t_L g3380 ( 
.A(n_3124),
.B(n_3082),
.C(n_3184),
.Y(n_3380)
);

AO31x2_ASAP7_75t_L g3381 ( 
.A1(n_3115),
.A2(n_1770),
.A3(n_1750),
.B(n_1886),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3010),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3181),
.Y(n_3383)
);

BUFx2_ASAP7_75t_L g3384 ( 
.A(n_3103),
.Y(n_3384)
);

AND2x4_ASAP7_75t_L g3385 ( 
.A(n_3086),
.B(n_228),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3153),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3153),
.Y(n_3387)
);

AOI22x1_ASAP7_75t_L g3388 ( 
.A1(n_3100),
.A2(n_910),
.B1(n_1592),
.B2(n_52),
.Y(n_3388)
);

AOI22xp33_ASAP7_75t_L g3389 ( 
.A1(n_3161),
.A2(n_1622),
.B1(n_1626),
.B2(n_1602),
.Y(n_3389)
);

NOR2xp33_ASAP7_75t_SL g3390 ( 
.A(n_3067),
.B(n_2016),
.Y(n_3390)
);

INVx3_ASAP7_75t_L g3391 ( 
.A(n_3139),
.Y(n_3391)
);

AOI22xp33_ASAP7_75t_L g3392 ( 
.A1(n_3161),
.A2(n_1622),
.B1(n_1626),
.B2(n_1602),
.Y(n_3392)
);

AOI21xp33_ASAP7_75t_L g3393 ( 
.A1(n_3188),
.A2(n_1906),
.B(n_1886),
.Y(n_3393)
);

A2O1A1Ixp33_ASAP7_75t_L g3394 ( 
.A1(n_3160),
.A2(n_52),
.B(n_46),
.C(n_51),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3080),
.Y(n_3395)
);

BUFx2_ASAP7_75t_L g3396 ( 
.A(n_3126),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3173),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3176),
.Y(n_3398)
);

NOR2xp33_ASAP7_75t_L g3399 ( 
.A(n_3127),
.B(n_54),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3010),
.Y(n_3400)
);

AOI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_3136),
.A2(n_2025),
.B(n_2016),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3176),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_3014),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3301),
.B(n_3161),
.Y(n_3404)
);

BUFx6f_ASAP7_75t_L g3405 ( 
.A(n_3267),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3220),
.Y(n_3406)
);

OAI22xp33_ASAP7_75t_L g3407 ( 
.A1(n_3214),
.A2(n_3050),
.B1(n_3175),
.B2(n_3077),
.Y(n_3407)
);

BUFx3_ASAP7_75t_L g3408 ( 
.A(n_3230),
.Y(n_3408)
);

O2A1O1Ixp33_ASAP7_75t_L g3409 ( 
.A1(n_3346),
.A2(n_3186),
.B(n_3131),
.C(n_3128),
.Y(n_3409)
);

INVx2_ASAP7_75t_SL g3410 ( 
.A(n_3267),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3202),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3210),
.Y(n_3412)
);

BUFx2_ASAP7_75t_L g3413 ( 
.A(n_3242),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_3201),
.A2(n_3136),
.B(n_3175),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_SL g3415 ( 
.A(n_3380),
.B(n_3144),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3369),
.B(n_3113),
.Y(n_3416)
);

INVx3_ASAP7_75t_SL g3417 ( 
.A(n_3227),
.Y(n_3417)
);

INVx1_ASAP7_75t_SL g3418 ( 
.A(n_3234),
.Y(n_3418)
);

INVx2_ASAP7_75t_SL g3419 ( 
.A(n_3267),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3228),
.Y(n_3420)
);

AND2x4_ASAP7_75t_SL g3421 ( 
.A(n_3224),
.B(n_3075),
.Y(n_3421)
);

AND2x2_ASAP7_75t_L g3422 ( 
.A(n_3317),
.B(n_3199),
.Y(n_3422)
);

BUFx6f_ASAP7_75t_L g3423 ( 
.A(n_3252),
.Y(n_3423)
);

AND2x4_ASAP7_75t_L g3424 ( 
.A(n_3223),
.B(n_3182),
.Y(n_3424)
);

INVx2_ASAP7_75t_SL g3425 ( 
.A(n_3198),
.Y(n_3425)
);

BUFx6f_ASAP7_75t_L g3426 ( 
.A(n_3197),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_3238),
.Y(n_3427)
);

INVx2_ASAP7_75t_SL g3428 ( 
.A(n_3265),
.Y(n_3428)
);

INVx3_ASAP7_75t_L g3429 ( 
.A(n_3237),
.Y(n_3429)
);

BUFx12f_ASAP7_75t_L g3430 ( 
.A(n_3232),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3253),
.Y(n_3431)
);

NOR2xp67_ASAP7_75t_SL g3432 ( 
.A(n_3192),
.B(n_3144),
.Y(n_3432)
);

HB1xp67_ASAP7_75t_L g3433 ( 
.A(n_3340),
.Y(n_3433)
);

AOI22xp5_ASAP7_75t_L g3434 ( 
.A1(n_3347),
.A2(n_3107),
.B1(n_3175),
.B2(n_3118),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_3251),
.B(n_3014),
.Y(n_3435)
);

A2O1A1Ixp33_ASAP7_75t_L g3436 ( 
.A1(n_3300),
.A2(n_3149),
.B(n_3104),
.C(n_3162),
.Y(n_3436)
);

BUFx2_ASAP7_75t_L g3437 ( 
.A(n_3269),
.Y(n_3437)
);

NOR2x1_ASAP7_75t_L g3438 ( 
.A(n_3286),
.B(n_3386),
.Y(n_3438)
);

AND2x4_ASAP7_75t_L g3439 ( 
.A(n_3395),
.B(n_3170),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_3212),
.Y(n_3440)
);

NOR2x1_ASAP7_75t_SL g3441 ( 
.A(n_3387),
.B(n_3155),
.Y(n_3441)
);

AND2x2_ASAP7_75t_L g3442 ( 
.A(n_3285),
.B(n_3017),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3213),
.Y(n_3443)
);

NOR2xp67_ASAP7_75t_L g3444 ( 
.A(n_3329),
.B(n_3123),
.Y(n_3444)
);

OAI21x1_ASAP7_75t_L g3445 ( 
.A1(n_3205),
.A2(n_3061),
.B(n_3109),
.Y(n_3445)
);

AND2x2_ASAP7_75t_L g3446 ( 
.A(n_3247),
.B(n_3017),
.Y(n_3446)
);

AOI22xp33_ASAP7_75t_L g3447 ( 
.A1(n_3333),
.A2(n_3170),
.B1(n_3087),
.B2(n_3119),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3219),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3258),
.Y(n_3449)
);

OAI22xp5_ASAP7_75t_L g3450 ( 
.A1(n_3394),
.A2(n_3036),
.B1(n_3112),
.B2(n_3109),
.Y(n_3450)
);

AOI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_3315),
.A2(n_3278),
.B1(n_3263),
.B2(n_3235),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3331),
.Y(n_3452)
);

HB1xp67_ASAP7_75t_L g3453 ( 
.A(n_3370),
.Y(n_3453)
);

INVx2_ASAP7_75t_L g3454 ( 
.A(n_3264),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_3230),
.Y(n_3455)
);

OR2x6_ASAP7_75t_L g3456 ( 
.A(n_3319),
.B(n_3155),
.Y(n_3456)
);

OR2x6_ASAP7_75t_L g3457 ( 
.A(n_3336),
.B(n_3155),
.Y(n_3457)
);

AOI21xp5_ASAP7_75t_L g3458 ( 
.A1(n_3194),
.A2(n_3112),
.B(n_3123),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3272),
.Y(n_3459)
);

INVx3_ASAP7_75t_L g3460 ( 
.A(n_3237),
.Y(n_3460)
);

INVx1_ASAP7_75t_SL g3461 ( 
.A(n_3204),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_L g3462 ( 
.A1(n_3206),
.A2(n_3095),
.B1(n_3075),
.B2(n_3149),
.Y(n_3462)
);

AND2x6_ASAP7_75t_L g3463 ( 
.A(n_3243),
.B(n_3095),
.Y(n_3463)
);

INVx2_ASAP7_75t_SL g3464 ( 
.A(n_3355),
.Y(n_3464)
);

BUFx6f_ASAP7_75t_L g3465 ( 
.A(n_3197),
.Y(n_3465)
);

AOI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_3292),
.A2(n_3091),
.B(n_2001),
.Y(n_3466)
);

INVxp67_ASAP7_75t_SL g3467 ( 
.A(n_3377),
.Y(n_3467)
);

A2O1A1Ixp33_ASAP7_75t_L g3468 ( 
.A1(n_3345),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_3468)
);

NAND3xp33_ASAP7_75t_L g3469 ( 
.A(n_3294),
.B(n_910),
.C(n_55),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3363),
.B(n_58),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3313),
.B(n_59),
.Y(n_3471)
);

OR2x6_ASAP7_75t_L g3472 ( 
.A(n_3401),
.B(n_3273),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3190),
.B(n_59),
.Y(n_3473)
);

BUFx6f_ASAP7_75t_L g3474 ( 
.A(n_3197),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3195),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3302),
.B(n_60),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3275),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3280),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_3342),
.B(n_60),
.Y(n_3479)
);

INVxp67_ASAP7_75t_SL g3480 ( 
.A(n_3321),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3281),
.Y(n_3481)
);

OAI22xp5_ASAP7_75t_L g3482 ( 
.A1(n_3367),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_3482)
);

INVx3_ASAP7_75t_L g3483 ( 
.A(n_3248),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3366),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3318),
.Y(n_3485)
);

HB1xp67_ASAP7_75t_L g3486 ( 
.A(n_3332),
.Y(n_3486)
);

AOI221xp5_ASAP7_75t_L g3487 ( 
.A1(n_3320),
.A2(n_67),
.B1(n_62),
.B2(n_66),
.C(n_68),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_3396),
.B(n_66),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3297),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3330),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3351),
.B(n_68),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3337),
.B(n_70),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_SL g3493 ( 
.A1(n_3388),
.A2(n_75),
.B1(n_72),
.B2(n_73),
.Y(n_3493)
);

HB1xp67_ASAP7_75t_L g3494 ( 
.A(n_3397),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3361),
.B(n_73),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3287),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3384),
.B(n_75),
.Y(n_3497)
);

INVx2_ASAP7_75t_SL g3498 ( 
.A(n_3355),
.Y(n_3498)
);

AOI222xp33_ASAP7_75t_L g3499 ( 
.A1(n_3399),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.C1(n_82),
.C2(n_83),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3293),
.Y(n_3500)
);

BUFx2_ASAP7_75t_L g3501 ( 
.A(n_3290),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3372),
.B(n_77),
.Y(n_3502)
);

HB1xp67_ASAP7_75t_L g3503 ( 
.A(n_3398),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3375),
.B(n_84),
.Y(n_3504)
);

INVxp67_ASAP7_75t_SL g3505 ( 
.A(n_3402),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3307),
.Y(n_3506)
);

NOR2xp33_ASAP7_75t_L g3507 ( 
.A(n_3191),
.B(n_3226),
.Y(n_3507)
);

NAND3xp33_ASAP7_75t_L g3508 ( 
.A(n_3241),
.B(n_910),
.C(n_84),
.Y(n_3508)
);

CKINVDCx5p33_ASAP7_75t_R g3509 ( 
.A(n_3225),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_3323),
.Y(n_3510)
);

BUFx3_ASAP7_75t_L g3511 ( 
.A(n_3271),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3305),
.A2(n_2001),
.B(n_1906),
.Y(n_3512)
);

BUFx6f_ASAP7_75t_L g3513 ( 
.A(n_3200),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_3303),
.A2(n_2001),
.B(n_1906),
.Y(n_3514)
);

INVx3_ASAP7_75t_L g3515 ( 
.A(n_3248),
.Y(n_3515)
);

INVx4_ASAP7_75t_L g3516 ( 
.A(n_3200),
.Y(n_3516)
);

AND2x2_ASAP7_75t_L g3517 ( 
.A(n_3290),
.B(n_85),
.Y(n_3517)
);

OR2x2_ASAP7_75t_L g3518 ( 
.A(n_3356),
.B(n_85),
.Y(n_3518)
);

INVx2_ASAP7_75t_SL g3519 ( 
.A(n_3364),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3314),
.B(n_86),
.Y(n_3520)
);

INVx6_ASAP7_75t_L g3521 ( 
.A(n_3299),
.Y(n_3521)
);

CKINVDCx20_ASAP7_75t_R g3522 ( 
.A(n_3279),
.Y(n_3522)
);

BUFx3_ASAP7_75t_L g3523 ( 
.A(n_3200),
.Y(n_3523)
);

OR2x2_ASAP7_75t_L g3524 ( 
.A(n_3334),
.B(n_3325),
.Y(n_3524)
);

OAI21x1_ASAP7_75t_L g3525 ( 
.A1(n_3211),
.A2(n_1750),
.B(n_2008),
.Y(n_3525)
);

BUFx2_ASAP7_75t_L g3526 ( 
.A(n_3291),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3383),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3358),
.Y(n_3528)
);

AND2x2_ASAP7_75t_L g3529 ( 
.A(n_3291),
.B(n_86),
.Y(n_3529)
);

BUFx6f_ASAP7_75t_L g3530 ( 
.A(n_3203),
.Y(n_3530)
);

INVx2_ASAP7_75t_SL g3531 ( 
.A(n_3364),
.Y(n_3531)
);

BUFx3_ASAP7_75t_L g3532 ( 
.A(n_3203),
.Y(n_3532)
);

AND2x2_ASAP7_75t_L g3533 ( 
.A(n_3304),
.B(n_87),
.Y(n_3533)
);

BUFx2_ASAP7_75t_L g3534 ( 
.A(n_3391),
.Y(n_3534)
);

INVx3_ASAP7_75t_L g3535 ( 
.A(n_3391),
.Y(n_3535)
);

AND2x2_ASAP7_75t_L g3536 ( 
.A(n_3304),
.B(n_87),
.Y(n_3536)
);

INVxp67_ASAP7_75t_L g3537 ( 
.A(n_3231),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3382),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3400),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3403),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3233),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3240),
.Y(n_3542)
);

AND2x4_ASAP7_75t_L g3543 ( 
.A(n_3329),
.B(n_88),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3359),
.B(n_90),
.Y(n_3544)
);

INVx3_ASAP7_75t_L g3545 ( 
.A(n_3379),
.Y(n_3545)
);

AND2x2_ASAP7_75t_SL g3546 ( 
.A(n_3245),
.B(n_91),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3371),
.B(n_92),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3207),
.Y(n_3548)
);

INVx2_ASAP7_75t_SL g3549 ( 
.A(n_3203),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3365),
.A2(n_2008),
.B(n_2016),
.Y(n_3550)
);

AND2x4_ASAP7_75t_L g3551 ( 
.A(n_3329),
.B(n_3308),
.Y(n_3551)
);

AOI22xp33_ASAP7_75t_L g3552 ( 
.A1(n_3362),
.A2(n_1622),
.B1(n_1626),
.B2(n_1602),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3308),
.B(n_3327),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3218),
.Y(n_3554)
);

OAI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3374),
.A2(n_2008),
.B(n_1881),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3217),
.Y(n_3556)
);

OR2x6_ASAP7_75t_L g3557 ( 
.A(n_3289),
.B(n_1626),
.Y(n_3557)
);

INVx1_ASAP7_75t_SL g3558 ( 
.A(n_3260),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3262),
.Y(n_3559)
);

INVx3_ASAP7_75t_L g3560 ( 
.A(n_3379),
.Y(n_3560)
);

CKINVDCx20_ASAP7_75t_R g3561 ( 
.A(n_3216),
.Y(n_3561)
);

AOI22xp33_ASAP7_75t_SL g3562 ( 
.A1(n_3215),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_3562)
);

CKINVDCx8_ASAP7_75t_R g3563 ( 
.A(n_3208),
.Y(n_3563)
);

INVx2_ASAP7_75t_SL g3564 ( 
.A(n_3208),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_3352),
.A2(n_2028),
.B(n_2025),
.Y(n_3565)
);

AND2x4_ASAP7_75t_L g3566 ( 
.A(n_3260),
.B(n_95),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_3322),
.A2(n_2028),
.B(n_2025),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3249),
.B(n_96),
.Y(n_3568)
);

O2A1O1Ixp5_ASAP7_75t_SL g3569 ( 
.A1(n_3268),
.A2(n_1584),
.B(n_1583),
.C(n_1475),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3284),
.B(n_97),
.Y(n_3570)
);

CKINVDCx5p33_ASAP7_75t_R g3571 ( 
.A(n_3208),
.Y(n_3571)
);

BUFx2_ASAP7_75t_L g3572 ( 
.A(n_3268),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3270),
.B(n_97),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3217),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_3348),
.Y(n_3575)
);

AO32x2_ASAP7_75t_L g3576 ( 
.A1(n_3428),
.A2(n_3324),
.A3(n_3310),
.B1(n_3309),
.B2(n_3266),
.Y(n_3576)
);

OAI21x1_ASAP7_75t_L g3577 ( 
.A1(n_3414),
.A2(n_3298),
.B(n_3306),
.Y(n_3577)
);

INVx3_ASAP7_75t_L g3578 ( 
.A(n_3429),
.Y(n_3578)
);

BUFx6f_ASAP7_75t_L g3579 ( 
.A(n_3408),
.Y(n_3579)
);

OR2x4_ASAP7_75t_L g3580 ( 
.A(n_3423),
.B(n_3507),
.Y(n_3580)
);

NAND2x1p5_ASAP7_75t_L g3581 ( 
.A(n_3438),
.B(n_3316),
.Y(n_3581)
);

AOI22xp5_ASAP7_75t_L g3582 ( 
.A1(n_3451),
.A2(n_3350),
.B1(n_3338),
.B2(n_3341),
.Y(n_3582)
);

AND2x4_ASAP7_75t_L g3583 ( 
.A(n_3424),
.B(n_3276),
.Y(n_3583)
);

OAI221xp5_ASAP7_75t_L g3584 ( 
.A1(n_3451),
.A2(n_3193),
.B1(n_3196),
.B2(n_3339),
.C(n_3357),
.Y(n_3584)
);

A2O1A1Ixp33_ASAP7_75t_L g3585 ( 
.A1(n_3469),
.A2(n_3282),
.B(n_3335),
.C(n_3254),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3452),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3411),
.Y(n_3587)
);

BUFx3_ASAP7_75t_L g3588 ( 
.A(n_3522),
.Y(n_3588)
);

AOI21x1_ASAP7_75t_L g3589 ( 
.A1(n_3432),
.A2(n_3378),
.B(n_3236),
.Y(n_3589)
);

NOR2x1_ASAP7_75t_R g3590 ( 
.A(n_3430),
.B(n_3385),
.Y(n_3590)
);

OAI21x1_ASAP7_75t_L g3591 ( 
.A1(n_3445),
.A2(n_3368),
.B(n_3259),
.Y(n_3591)
);

OR2x2_ASAP7_75t_L g3592 ( 
.A(n_3461),
.B(n_3221),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3412),
.Y(n_3593)
);

BUFx3_ASAP7_75t_L g3594 ( 
.A(n_3509),
.Y(n_3594)
);

OAI21x1_ASAP7_75t_L g3595 ( 
.A1(n_3438),
.A2(n_3246),
.B(n_3239),
.Y(n_3595)
);

AOI21xp5_ASAP7_75t_L g3596 ( 
.A1(n_3514),
.A2(n_3353),
.B(n_3256),
.Y(n_3596)
);

CKINVDCx5p33_ASAP7_75t_R g3597 ( 
.A(n_3455),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3448),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3449),
.Y(n_3599)
);

OAI21x1_ASAP7_75t_L g3600 ( 
.A1(n_3458),
.A2(n_3250),
.B(n_3261),
.Y(n_3600)
);

NAND2x1p5_ASAP7_75t_L g3601 ( 
.A(n_3444),
.B(n_3316),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3486),
.B(n_3480),
.Y(n_3602)
);

OAI21x1_ASAP7_75t_L g3603 ( 
.A1(n_3466),
.A2(n_3276),
.B(n_3274),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3485),
.Y(n_3604)
);

OAI21x1_ASAP7_75t_L g3605 ( 
.A1(n_3415),
.A2(n_3326),
.B(n_3209),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3413),
.Y(n_3606)
);

OAI21x1_ASAP7_75t_L g3607 ( 
.A1(n_3568),
.A2(n_3277),
.B(n_3376),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_L g3608 ( 
.A(n_3537),
.B(n_3360),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3461),
.B(n_3362),
.Y(n_3609)
);

NAND2x1p5_ASAP7_75t_L g3610 ( 
.A(n_3444),
.B(n_3373),
.Y(n_3610)
);

HB1xp67_ASAP7_75t_L g3611 ( 
.A(n_3453),
.Y(n_3611)
);

AOI22xp33_ASAP7_75t_L g3612 ( 
.A1(n_3499),
.A2(n_3362),
.B1(n_3385),
.B2(n_3373),
.Y(n_3612)
);

CKINVDCx11_ASAP7_75t_R g3613 ( 
.A(n_3417),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3467),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3490),
.B(n_3362),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3478),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3440),
.Y(n_3617)
);

BUFx2_ASAP7_75t_L g3618 ( 
.A(n_3551),
.Y(n_3618)
);

NOR4xp25_ASAP7_75t_L g3619 ( 
.A(n_3508),
.B(n_3288),
.C(n_3257),
.D(n_3244),
.Y(n_3619)
);

OAI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_3469),
.A2(n_3311),
.B(n_3312),
.Y(n_3620)
);

O2A1O1Ixp5_ASAP7_75t_L g3621 ( 
.A1(n_3508),
.A2(n_3255),
.B(n_3354),
.C(n_3296),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3443),
.Y(n_3622)
);

OAI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_3468),
.A2(n_3255),
.B(n_3390),
.Y(n_3623)
);

BUFx6f_ASAP7_75t_L g3624 ( 
.A(n_3405),
.Y(n_3624)
);

OAI21x1_ASAP7_75t_L g3625 ( 
.A1(n_3568),
.A2(n_3392),
.B(n_3389),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3437),
.Y(n_3626)
);

CKINVDCx5p33_ASAP7_75t_R g3627 ( 
.A(n_3561),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3433),
.B(n_3222),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3475),
.Y(n_3629)
);

NOR2x1_ASAP7_75t_SL g3630 ( 
.A(n_3456),
.B(n_3295),
.Y(n_3630)
);

AOI22xp33_ASAP7_75t_SL g3631 ( 
.A1(n_3546),
.A2(n_3373),
.B1(n_3229),
.B2(n_3222),
.Y(n_3631)
);

OAI21x1_ASAP7_75t_L g3632 ( 
.A1(n_3525),
.A2(n_3283),
.B(n_3343),
.Y(n_3632)
);

NAND3xp33_ASAP7_75t_SL g3633 ( 
.A(n_3434),
.B(n_3499),
.C(n_3436),
.Y(n_3633)
);

AND2x4_ASAP7_75t_L g3634 ( 
.A(n_3424),
.B(n_3222),
.Y(n_3634)
);

AOI22xp33_ASAP7_75t_L g3635 ( 
.A1(n_3482),
.A2(n_3354),
.B1(n_3229),
.B2(n_3344),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_3422),
.Y(n_3636)
);

HB1xp67_ASAP7_75t_L g3637 ( 
.A(n_3418),
.Y(n_3637)
);

OAI21x1_ASAP7_75t_L g3638 ( 
.A1(n_3512),
.A2(n_3381),
.B(n_1881),
.Y(n_3638)
);

OA21x2_ASAP7_75t_L g3639 ( 
.A1(n_3476),
.A2(n_3393),
.B(n_3381),
.Y(n_3639)
);

AOI21x1_ASAP7_75t_L g3640 ( 
.A1(n_3476),
.A2(n_3328),
.B(n_3295),
.Y(n_3640)
);

AOI221x1_ASAP7_75t_L g3641 ( 
.A1(n_3559),
.A2(n_3229),
.B1(n_3381),
.B2(n_101),
.C(n_103),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3481),
.Y(n_3642)
);

A2O1A1Ixp33_ASAP7_75t_L g3643 ( 
.A1(n_3434),
.A2(n_3487),
.B(n_3409),
.C(n_3482),
.Y(n_3643)
);

AO32x2_ASAP7_75t_L g3644 ( 
.A1(n_3450),
.A2(n_3328),
.A3(n_100),
.B1(n_101),
.B2(n_107),
.Y(n_3644)
);

HB1xp67_ASAP7_75t_L g3645 ( 
.A(n_3418),
.Y(n_3645)
);

AOI22xp33_ASAP7_75t_L g3646 ( 
.A1(n_3407),
.A2(n_3349),
.B1(n_1488),
.B2(n_1512),
.Y(n_3646)
);

INVx1_ASAP7_75t_SL g3647 ( 
.A(n_3534),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3496),
.B(n_98),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3406),
.Y(n_3649)
);

HB1xp67_ASAP7_75t_L g3650 ( 
.A(n_3494),
.Y(n_3650)
);

OAI22xp5_ASAP7_75t_L g3651 ( 
.A1(n_3493),
.A2(n_108),
.B1(n_98),
.B2(n_107),
.Y(n_3651)
);

AND2x4_ASAP7_75t_L g3652 ( 
.A(n_3439),
.B(n_108),
.Y(n_3652)
);

INVx2_ASAP7_75t_SL g3653 ( 
.A(n_3521),
.Y(n_3653)
);

AOI21x1_ASAP7_75t_L g3654 ( 
.A1(n_3479),
.A2(n_1881),
.B(n_110),
.Y(n_3654)
);

OAI21x1_ASAP7_75t_L g3655 ( 
.A1(n_3567),
.A2(n_1469),
.B(n_1533),
.Y(n_3655)
);

HB1xp67_ASAP7_75t_L g3656 ( 
.A(n_3503),
.Y(n_3656)
);

AOI22xp33_ASAP7_75t_L g3657 ( 
.A1(n_3463),
.A2(n_1488),
.B1(n_1512),
.B2(n_1490),
.Y(n_3657)
);

A2O1A1Ixp33_ASAP7_75t_L g3658 ( 
.A1(n_3471),
.A2(n_113),
.B(n_110),
.C(n_112),
.Y(n_3658)
);

INVx1_ASAP7_75t_SL g3659 ( 
.A(n_3501),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3420),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3538),
.Y(n_3661)
);

OAI21x1_ASAP7_75t_L g3662 ( 
.A1(n_3404),
.A2(n_1572),
.B(n_1558),
.Y(n_3662)
);

HB1xp67_ASAP7_75t_L g3663 ( 
.A(n_3524),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_L g3664 ( 
.A1(n_3463),
.A2(n_1488),
.B1(n_1512),
.B2(n_1490),
.Y(n_3664)
);

AND2x4_ASAP7_75t_L g3665 ( 
.A(n_3439),
.B(n_112),
.Y(n_3665)
);

OAI21x1_ASAP7_75t_SL g3666 ( 
.A1(n_3441),
.A2(n_115),
.B(n_116),
.Y(n_3666)
);

BUFx3_ASAP7_75t_L g3667 ( 
.A(n_3511),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3454),
.B(n_115),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3540),
.Y(n_3669)
);

AOI22xp5_ASAP7_75t_L g3670 ( 
.A1(n_3562),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_3670)
);

OAI21x1_ASAP7_75t_L g3671 ( 
.A1(n_3404),
.A2(n_1572),
.B(n_1558),
.Y(n_3671)
);

OAI21x1_ASAP7_75t_L g3672 ( 
.A1(n_3569),
.A2(n_1572),
.B(n_118),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3427),
.Y(n_3673)
);

HB1xp67_ASAP7_75t_L g3674 ( 
.A(n_3539),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3459),
.B(n_120),
.Y(n_3675)
);

OAI21x1_ASAP7_75t_L g3676 ( 
.A1(n_3550),
.A2(n_121),
.B(n_122),
.Y(n_3676)
);

OAI21x1_ASAP7_75t_L g3677 ( 
.A1(n_3565),
.A2(n_122),
.B(n_123),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3431),
.Y(n_3678)
);

CKINVDCx11_ASAP7_75t_R g3679 ( 
.A(n_3423),
.Y(n_3679)
);

INVx3_ASAP7_75t_L g3680 ( 
.A(n_3429),
.Y(n_3680)
);

HB1xp67_ASAP7_75t_L g3681 ( 
.A(n_3505),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3526),
.B(n_123),
.Y(n_3682)
);

INVx2_ASAP7_75t_L g3683 ( 
.A(n_3477),
.Y(n_3683)
);

INVx2_ASAP7_75t_L g3684 ( 
.A(n_3500),
.Y(n_3684)
);

INVx8_ASAP7_75t_L g3685 ( 
.A(n_3543),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3460),
.A2(n_124),
.B(n_126),
.Y(n_3686)
);

OAI21x1_ASAP7_75t_L g3687 ( 
.A1(n_3460),
.A2(n_124),
.B(n_126),
.Y(n_3687)
);

OAI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_3450),
.A2(n_127),
.B(n_128),
.Y(n_3688)
);

O2A1O1Ixp33_ASAP7_75t_SL g3689 ( 
.A1(n_3520),
.A2(n_132),
.B(n_128),
.C(n_129),
.Y(n_3689)
);

AOI221xp5_ASAP7_75t_L g3690 ( 
.A1(n_3570),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.C(n_134),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3484),
.B(n_133),
.Y(n_3691)
);

NAND2x1p5_ASAP7_75t_L g3692 ( 
.A(n_3551),
.B(n_2028),
.Y(n_3692)
);

OAI21x1_ASAP7_75t_L g3693 ( 
.A1(n_3483),
.A2(n_134),
.B(n_136),
.Y(n_3693)
);

BUFx6f_ASAP7_75t_L g3694 ( 
.A(n_3405),
.Y(n_3694)
);

INVx5_ASAP7_75t_L g3695 ( 
.A(n_3456),
.Y(n_3695)
);

AO31x2_ASAP7_75t_L g3696 ( 
.A1(n_3489),
.A2(n_139),
.A3(n_136),
.B(n_137),
.Y(n_3696)
);

OAI21x1_ASAP7_75t_L g3697 ( 
.A1(n_3483),
.A2(n_141),
.B(n_143),
.Y(n_3697)
);

INVx3_ASAP7_75t_L g3698 ( 
.A(n_3515),
.Y(n_3698)
);

BUFx2_ASAP7_75t_L g3699 ( 
.A(n_3572),
.Y(n_3699)
);

BUFx8_ASAP7_75t_L g3700 ( 
.A(n_3423),
.Y(n_3700)
);

OAI22xp33_ASAP7_75t_L g3701 ( 
.A1(n_3456),
.A2(n_144),
.B1(n_141),
.B2(n_143),
.Y(n_3701)
);

OA21x2_ASAP7_75t_L g3702 ( 
.A1(n_3502),
.A2(n_147),
.B(n_148),
.Y(n_3702)
);

INVx6_ASAP7_75t_L g3703 ( 
.A(n_3521),
.Y(n_3703)
);

AND2x2_ASAP7_75t_L g3704 ( 
.A(n_3442),
.B(n_147),
.Y(n_3704)
);

AND2x2_ASAP7_75t_L g3705 ( 
.A(n_3553),
.B(n_3435),
.Y(n_3705)
);

A2O1A1Ixp33_ASAP7_75t_L g3706 ( 
.A1(n_3544),
.A2(n_149),
.B(n_151),
.C(n_152),
.Y(n_3706)
);

AOI21x1_ASAP7_75t_L g3707 ( 
.A1(n_3504),
.A2(n_3470),
.B(n_3491),
.Y(n_3707)
);

CKINVDCx11_ASAP7_75t_R g3708 ( 
.A(n_3563),
.Y(n_3708)
);

NOR3xp33_ASAP7_75t_L g3709 ( 
.A(n_3547),
.B(n_149),
.C(n_152),
.Y(n_3709)
);

OAI21x1_ASAP7_75t_L g3710 ( 
.A1(n_3515),
.A2(n_3555),
.B(n_3545),
.Y(n_3710)
);

OAI21x1_ASAP7_75t_L g3711 ( 
.A1(n_3555),
.A2(n_153),
.B(n_154),
.Y(n_3711)
);

INVx2_ASAP7_75t_L g3712 ( 
.A(n_3506),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3614),
.B(n_3541),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3699),
.Y(n_3714)
);

AOI22xp33_ASAP7_75t_L g3715 ( 
.A1(n_3633),
.A2(n_3447),
.B1(n_3518),
.B2(n_3575),
.Y(n_3715)
);

BUFx3_ASAP7_75t_L g3716 ( 
.A(n_3700),
.Y(n_3716)
);

OAI22xp33_ASAP7_75t_L g3717 ( 
.A1(n_3580),
.A2(n_3548),
.B1(n_3554),
.B2(n_3542),
.Y(n_3717)
);

INVx3_ASAP7_75t_L g3718 ( 
.A(n_3578),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_3578),
.Y(n_3719)
);

BUFx2_ASAP7_75t_L g3720 ( 
.A(n_3618),
.Y(n_3720)
);

OA21x2_ASAP7_75t_L g3721 ( 
.A1(n_3710),
.A2(n_3527),
.B(n_3574),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_3680),
.Y(n_3722)
);

HB1xp67_ASAP7_75t_L g3723 ( 
.A(n_3681),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3586),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3680),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3663),
.B(n_3510),
.Y(n_3726)
);

AO21x2_ASAP7_75t_L g3727 ( 
.A1(n_3688),
.A2(n_3573),
.B(n_3473),
.Y(n_3727)
);

AOI22xp33_ASAP7_75t_L g3728 ( 
.A1(n_3709),
.A2(n_3463),
.B1(n_3543),
.B2(n_3566),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3587),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3698),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3593),
.Y(n_3731)
);

BUFx4f_ASAP7_75t_SL g3732 ( 
.A(n_3700),
.Y(n_3732)
);

AO21x1_ASAP7_75t_SL g3733 ( 
.A1(n_3609),
.A2(n_3528),
.B(n_3552),
.Y(n_3733)
);

INVx3_ASAP7_75t_L g3734 ( 
.A(n_3698),
.Y(n_3734)
);

INVx2_ASAP7_75t_L g3735 ( 
.A(n_3629),
.Y(n_3735)
);

NOR2xp33_ASAP7_75t_L g3736 ( 
.A(n_3584),
.B(n_3488),
.Y(n_3736)
);

INVx1_ASAP7_75t_SL g3737 ( 
.A(n_3613),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_L g3738 ( 
.A(n_3602),
.B(n_3558),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3598),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3599),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3616),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3602),
.B(n_3558),
.Y(n_3742)
);

OAI21x1_ASAP7_75t_L g3743 ( 
.A1(n_3577),
.A2(n_3535),
.B(n_3545),
.Y(n_3743)
);

AOI21x1_ASAP7_75t_L g3744 ( 
.A1(n_3707),
.A2(n_3529),
.B(n_3517),
.Y(n_3744)
);

INVx1_ASAP7_75t_SL g3745 ( 
.A(n_3679),
.Y(n_3745)
);

AOI22xp33_ASAP7_75t_L g3746 ( 
.A1(n_3584),
.A2(n_3463),
.B1(n_3566),
.B2(n_3416),
.Y(n_3746)
);

HB1xp67_ASAP7_75t_SL g3747 ( 
.A(n_3652),
.Y(n_3747)
);

BUFx2_ASAP7_75t_SL g3748 ( 
.A(n_3579),
.Y(n_3748)
);

BUFx6f_ASAP7_75t_SL g3749 ( 
.A(n_3579),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3642),
.Y(n_3750)
);

INVx3_ASAP7_75t_L g3751 ( 
.A(n_3583),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_SL g3752 ( 
.A1(n_3688),
.A2(n_3421),
.B1(n_3497),
.B2(n_3495),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3674),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3604),
.Y(n_3754)
);

BUFx2_ASAP7_75t_R g3755 ( 
.A(n_3597),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3650),
.Y(n_3756)
);

AOI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3648),
.A2(n_3425),
.B(n_3457),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3581),
.Y(n_3758)
);

AOI22xp5_ASAP7_75t_L g3759 ( 
.A1(n_3643),
.A2(n_3457),
.B1(n_3472),
.B2(n_3462),
.Y(n_3759)
);

BUFx3_ASAP7_75t_L g3760 ( 
.A(n_3703),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3656),
.Y(n_3761)
);

OAI22xp5_ASAP7_75t_L g3762 ( 
.A1(n_3612),
.A2(n_3457),
.B1(n_3472),
.B2(n_3556),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3581),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3617),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3649),
.Y(n_3765)
);

BUFx3_ASAP7_75t_L g3766 ( 
.A(n_3703),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3622),
.Y(n_3767)
);

AO21x2_ASAP7_75t_L g3768 ( 
.A1(n_3691),
.A2(n_3536),
.B(n_3533),
.Y(n_3768)
);

OAI21x1_ASAP7_75t_L g3769 ( 
.A1(n_3640),
.A2(n_3535),
.B(n_3560),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3660),
.Y(n_3770)
);

NAND2x1p5_ASAP7_75t_L g3771 ( 
.A(n_3695),
.B(n_3560),
.Y(n_3771)
);

INVx1_ASAP7_75t_SL g3772 ( 
.A(n_3708),
.Y(n_3772)
);

INVx4_ASAP7_75t_L g3773 ( 
.A(n_3579),
.Y(n_3773)
);

OAI21x1_ASAP7_75t_L g3774 ( 
.A1(n_3610),
.A2(n_3446),
.B(n_3492),
.Y(n_3774)
);

AOI22xp5_ASAP7_75t_L g3775 ( 
.A1(n_3651),
.A2(n_3472),
.B1(n_3498),
.B2(n_3464),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3673),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3678),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3683),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3611),
.Y(n_3779)
);

OAI21x1_ASAP7_75t_L g3780 ( 
.A1(n_3610),
.A2(n_3557),
.B(n_3516),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3637),
.Y(n_3781)
);

AO21x1_ASAP7_75t_L g3782 ( 
.A1(n_3645),
.A2(n_3516),
.B(n_3571),
.Y(n_3782)
);

BUFx3_ASAP7_75t_L g3783 ( 
.A(n_3588),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3661),
.Y(n_3784)
);

OAI21x1_ASAP7_75t_L g3785 ( 
.A1(n_3595),
.A2(n_3557),
.B(n_3419),
.Y(n_3785)
);

OAI22xp33_ASAP7_75t_L g3786 ( 
.A1(n_3580),
.A2(n_3557),
.B1(n_3519),
.B2(n_3531),
.Y(n_3786)
);

HB1xp67_ASAP7_75t_L g3787 ( 
.A(n_3669),
.Y(n_3787)
);

BUFx5_ASAP7_75t_L g3788 ( 
.A(n_3652),
.Y(n_3788)
);

NAND2x1p5_ASAP7_75t_L g3789 ( 
.A(n_3695),
.B(n_3405),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3684),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3712),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3647),
.Y(n_3792)
);

AOI22xp33_ASAP7_75t_L g3793 ( 
.A1(n_3690),
.A2(n_3523),
.B1(n_3532),
.B2(n_3410),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3592),
.Y(n_3794)
);

INVx11_ASAP7_75t_L g3795 ( 
.A(n_3627),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3615),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3606),
.Y(n_3797)
);

BUFx6f_ASAP7_75t_L g3798 ( 
.A(n_3644),
.Y(n_3798)
);

INVx2_ASAP7_75t_SL g3799 ( 
.A(n_3685),
.Y(n_3799)
);

AOI21x1_ASAP7_75t_L g3800 ( 
.A1(n_3648),
.A2(n_3564),
.B(n_3549),
.Y(n_3800)
);

OAI21x1_ASAP7_75t_L g3801 ( 
.A1(n_3609),
.A2(n_3465),
.B(n_3426),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3615),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3628),
.Y(n_3803)
);

AOI22xp5_ASAP7_75t_L g3804 ( 
.A1(n_3651),
.A2(n_3465),
.B1(n_3474),
.B2(n_3426),
.Y(n_3804)
);

NAND2x1p5_ASAP7_75t_L g3805 ( 
.A(n_3695),
.B(n_3426),
.Y(n_3805)
);

OA21x2_ASAP7_75t_L g3806 ( 
.A1(n_3641),
.A2(n_3474),
.B(n_3465),
.Y(n_3806)
);

AOI22xp5_ASAP7_75t_SL g3807 ( 
.A1(n_3665),
.A2(n_3530),
.B1(n_3513),
.B2(n_3474),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3690),
.A2(n_3670),
.B1(n_3582),
.B2(n_3701),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3628),
.Y(n_3809)
);

AOI22xp33_ASAP7_75t_SL g3810 ( 
.A1(n_3702),
.A2(n_3530),
.B1(n_3513),
.B2(n_155),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3668),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3647),
.Y(n_3812)
);

OAI21x1_ASAP7_75t_L g3813 ( 
.A1(n_3603),
.A2(n_3530),
.B(n_3513),
.Y(n_3813)
);

INVx2_ASAP7_75t_SL g3814 ( 
.A(n_3685),
.Y(n_3814)
);

INVx2_ASAP7_75t_SL g3815 ( 
.A(n_3685),
.Y(n_3815)
);

BUFx12f_ASAP7_75t_L g3816 ( 
.A(n_3653),
.Y(n_3816)
);

AOI22xp5_ASAP7_75t_L g3817 ( 
.A1(n_3670),
.A2(n_3631),
.B1(n_3620),
.B2(n_3582),
.Y(n_3817)
);

BUFx3_ASAP7_75t_L g3818 ( 
.A(n_3667),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3583),
.B(n_153),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3668),
.Y(n_3820)
);

AOI222xp33_ASAP7_75t_L g3821 ( 
.A1(n_3658),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.C1(n_158),
.C2(n_160),
.Y(n_3821)
);

AOI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_3620),
.A2(n_1490),
.B1(n_1512),
.B2(n_1524),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3675),
.Y(n_3823)
);

BUFx2_ASAP7_75t_SL g3824 ( 
.A(n_3594),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3675),
.Y(n_3825)
);

HB1xp67_ASAP7_75t_L g3826 ( 
.A(n_3702),
.Y(n_3826)
);

BUFx3_ASAP7_75t_L g3827 ( 
.A(n_3624),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3623),
.A2(n_3635),
.B1(n_3608),
.B2(n_3711),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3705),
.B(n_156),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_3636),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3691),
.Y(n_3831)
);

HB1xp67_ASAP7_75t_L g3832 ( 
.A(n_3696),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3659),
.Y(n_3833)
);

NAND2x1p5_ASAP7_75t_L g3834 ( 
.A(n_3659),
.B(n_2028),
.Y(n_3834)
);

AO21x1_ASAP7_75t_SL g3835 ( 
.A1(n_3623),
.A2(n_161),
.B(n_162),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3634),
.B(n_161),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3626),
.Y(n_3837)
);

INVx3_ASAP7_75t_L g3838 ( 
.A(n_3634),
.Y(n_3838)
);

HB1xp67_ASAP7_75t_L g3839 ( 
.A(n_3696),
.Y(n_3839)
);

INVx2_ASAP7_75t_SL g3840 ( 
.A(n_3760),
.Y(n_3840)
);

INVx4_ASAP7_75t_SL g3841 ( 
.A(n_3732),
.Y(n_3841)
);

HB1xp67_ASAP7_75t_L g3842 ( 
.A(n_3723),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3767),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3802),
.B(n_3630),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3724),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3723),
.Y(n_3846)
);

AOI22xp33_ASAP7_75t_L g3847 ( 
.A1(n_3808),
.A2(n_3646),
.B1(n_3666),
.B2(n_3607),
.Y(n_3847)
);

HB1xp67_ASAP7_75t_L g3848 ( 
.A(n_3826),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3729),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3731),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3767),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3784),
.Y(n_3852)
);

AND2x4_ASAP7_75t_SL g3853 ( 
.A(n_3773),
.B(n_3665),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3739),
.Y(n_3854)
);

HB1xp67_ASAP7_75t_L g3855 ( 
.A(n_3826),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3784),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3740),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3741),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3800),
.Y(n_3859)
);

BUFx2_ASAP7_75t_L g3860 ( 
.A(n_3720),
.Y(n_3860)
);

INVx3_ASAP7_75t_L g3861 ( 
.A(n_3771),
.Y(n_3861)
);

AOI222xp33_ASAP7_75t_L g3862 ( 
.A1(n_3808),
.A2(n_3706),
.B1(n_3585),
.B2(n_3590),
.C1(n_3682),
.C2(n_3704),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3750),
.Y(n_3863)
);

INVx3_ASAP7_75t_L g3864 ( 
.A(n_3771),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3802),
.Y(n_3865)
);

HB1xp67_ASAP7_75t_L g3866 ( 
.A(n_3832),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3765),
.Y(n_3867)
);

NOR2xp33_ASAP7_75t_SL g3868 ( 
.A(n_3755),
.B(n_3590),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3834),
.Y(n_3869)
);

BUFx2_ASAP7_75t_SL g3870 ( 
.A(n_3749),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3834),
.Y(n_3871)
);

OAI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3817),
.A2(n_3621),
.B(n_3605),
.Y(n_3872)
);

INVx3_ASAP7_75t_L g3873 ( 
.A(n_3789),
.Y(n_3873)
);

OAI21x1_ASAP7_75t_L g3874 ( 
.A1(n_3743),
.A2(n_3591),
.B(n_3601),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3797),
.Y(n_3875)
);

OAI21x1_ASAP7_75t_L g3876 ( 
.A1(n_3769),
.A2(n_3813),
.B(n_3780),
.Y(n_3876)
);

CKINVDCx11_ASAP7_75t_R g3877 ( 
.A(n_3745),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3770),
.Y(n_3878)
);

BUFx6f_ASAP7_75t_L g3879 ( 
.A(n_3716),
.Y(n_3879)
);

HB1xp67_ASAP7_75t_L g3880 ( 
.A(n_3832),
.Y(n_3880)
);

OAI21x1_ASAP7_75t_L g3881 ( 
.A1(n_3785),
.A2(n_3805),
.B(n_3789),
.Y(n_3881)
);

AND2x2_ASAP7_75t_L g3882 ( 
.A(n_3751),
.B(n_3601),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3776),
.Y(n_3883)
);

OR2x6_ASAP7_75t_L g3884 ( 
.A(n_3748),
.B(n_3676),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3797),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3838),
.B(n_3624),
.Y(n_3886)
);

OAI21x1_ASAP7_75t_L g3887 ( 
.A1(n_3805),
.A2(n_3638),
.B(n_3662),
.Y(n_3887)
);

BUFx2_ASAP7_75t_L g3888 ( 
.A(n_3760),
.Y(n_3888)
);

OR2x6_ASAP7_75t_L g3889 ( 
.A(n_3798),
.B(n_3600),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3777),
.Y(n_3890)
);

INVx3_ASAP7_75t_L g3891 ( 
.A(n_3798),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3713),
.Y(n_3892)
);

BUFx3_ASAP7_75t_L g3893 ( 
.A(n_3732),
.Y(n_3893)
);

AND2x4_ASAP7_75t_L g3894 ( 
.A(n_3838),
.B(n_3696),
.Y(n_3894)
);

BUFx3_ASAP7_75t_L g3895 ( 
.A(n_3716),
.Y(n_3895)
);

HB1xp67_ASAP7_75t_L g3896 ( 
.A(n_3839),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3744),
.Y(n_3897)
);

BUFx3_ASAP7_75t_L g3898 ( 
.A(n_3766),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3713),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3794),
.Y(n_3900)
);

BUFx3_ASAP7_75t_L g3901 ( 
.A(n_3766),
.Y(n_3901)
);

AOI22xp33_ASAP7_75t_SL g3902 ( 
.A1(n_3798),
.A2(n_3677),
.B1(n_3625),
.B2(n_3644),
.Y(n_3902)
);

AO21x2_ASAP7_75t_L g3903 ( 
.A1(n_3782),
.A2(n_3596),
.B(n_3689),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3751),
.B(n_3624),
.Y(n_3904)
);

HB1xp67_ASAP7_75t_L g3905 ( 
.A(n_3839),
.Y(n_3905)
);

AND2x2_ASAP7_75t_L g3906 ( 
.A(n_3799),
.B(n_3694),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3753),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3831),
.B(n_3619),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3726),
.Y(n_3909)
);

OR2x2_ASAP7_75t_L g3910 ( 
.A(n_3796),
.B(n_3639),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3726),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3754),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3721),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3721),
.Y(n_3914)
);

INVx1_ASAP7_75t_L g3915 ( 
.A(n_3787),
.Y(n_3915)
);

INVx2_ASAP7_75t_SL g3916 ( 
.A(n_3773),
.Y(n_3916)
);

OR2x6_ASAP7_75t_L g3917 ( 
.A(n_3798),
.B(n_3589),
.Y(n_3917)
);

INVx3_ASAP7_75t_L g3918 ( 
.A(n_3718),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_L g3919 ( 
.A(n_3736),
.B(n_3686),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3721),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3787),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3756),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3761),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3735),
.Y(n_3924)
);

AND2x2_ASAP7_75t_L g3925 ( 
.A(n_3758),
.B(n_3694),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3781),
.Y(n_3926)
);

INVx2_ASAP7_75t_L g3927 ( 
.A(n_3764),
.Y(n_3927)
);

OAI22xp33_ASAP7_75t_L g3928 ( 
.A1(n_3806),
.A2(n_3644),
.B1(n_3576),
.B2(n_3619),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3778),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3790),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3779),
.Y(n_3931)
);

CKINVDCx5p33_ASAP7_75t_R g3932 ( 
.A(n_3755),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3791),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3811),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3820),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3803),
.Y(n_3936)
);

INVx3_ASAP7_75t_L g3937 ( 
.A(n_3718),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3823),
.Y(n_3938)
);

INVx2_ASAP7_75t_L g3939 ( 
.A(n_3809),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3825),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3768),
.B(n_3694),
.Y(n_3941)
);

INVx1_ASAP7_75t_SL g3942 ( 
.A(n_3824),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3738),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3738),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3742),
.Y(n_3945)
);

INVx2_ASAP7_75t_L g3946 ( 
.A(n_3792),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3768),
.B(n_3687),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3742),
.Y(n_3948)
);

OR2x6_ASAP7_75t_L g3949 ( 
.A(n_3806),
.B(n_3671),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3763),
.B(n_3692),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3812),
.Y(n_3951)
);

AOI22xp33_ASAP7_75t_L g3952 ( 
.A1(n_3821),
.A2(n_3664),
.B1(n_3657),
.B2(n_3697),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3833),
.Y(n_3953)
);

HB1xp67_ASAP7_75t_SL g3954 ( 
.A(n_3747),
.Y(n_3954)
);

NAND2xp5_ASAP7_75t_L g3955 ( 
.A(n_3715),
.B(n_3693),
.Y(n_3955)
);

HB1xp67_ASAP7_75t_L g3956 ( 
.A(n_3757),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3837),
.Y(n_3957)
);

OAI21x1_ASAP7_75t_L g3958 ( 
.A1(n_3801),
.A2(n_3692),
.B(n_3639),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3830),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3714),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3827),
.Y(n_3961)
);

HB1xp67_ASAP7_75t_L g3962 ( 
.A(n_3727),
.Y(n_3962)
);

BUFx3_ASAP7_75t_L g3963 ( 
.A(n_3893),
.Y(n_3963)
);

AOI222xp33_ASAP7_75t_L g3964 ( 
.A1(n_3872),
.A2(n_3736),
.B1(n_3715),
.B2(n_3793),
.C1(n_3828),
.C2(n_3728),
.Y(n_3964)
);

BUFx12f_ASAP7_75t_L g3965 ( 
.A(n_3877),
.Y(n_3965)
);

BUFx2_ASAP7_75t_L g3966 ( 
.A(n_3898),
.Y(n_3966)
);

AOI21xp33_ASAP7_75t_L g3967 ( 
.A1(n_3928),
.A2(n_3903),
.B(n_3955),
.Y(n_3967)
);

NOR2xp33_ASAP7_75t_L g3968 ( 
.A(n_3932),
.B(n_3737),
.Y(n_3968)
);

AOI221xp5_ASAP7_75t_L g3969 ( 
.A1(n_3928),
.A2(n_3793),
.B1(n_3828),
.B2(n_3717),
.C(n_3810),
.Y(n_3969)
);

AOI22xp33_ASAP7_75t_L g3970 ( 
.A1(n_3903),
.A2(n_3727),
.B1(n_3762),
.B2(n_3746),
.Y(n_3970)
);

OAI221xp5_ASAP7_75t_L g3971 ( 
.A1(n_3902),
.A2(n_3810),
.B1(n_3759),
.B2(n_3746),
.C(n_3775),
.Y(n_3971)
);

AOI22xp33_ASAP7_75t_L g3972 ( 
.A1(n_3919),
.A2(n_3762),
.B1(n_3835),
.B2(n_3728),
.Y(n_3972)
);

AOI21xp5_ASAP7_75t_L g3973 ( 
.A1(n_3868),
.A2(n_3717),
.B(n_3772),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3888),
.B(n_3807),
.Y(n_3974)
);

AOI22xp33_ASAP7_75t_L g3975 ( 
.A1(n_3919),
.A2(n_3806),
.B1(n_3752),
.B2(n_3788),
.Y(n_3975)
);

CKINVDCx5p33_ASAP7_75t_R g3976 ( 
.A(n_3877),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3848),
.Y(n_3977)
);

OAI22xp33_ASAP7_75t_L g3978 ( 
.A1(n_3917),
.A2(n_3804),
.B1(n_3786),
.B2(n_3814),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3886),
.B(n_3815),
.Y(n_3979)
);

AOI221xp5_ASAP7_75t_L g3980 ( 
.A1(n_3908),
.A2(n_3786),
.B1(n_3752),
.B2(n_3836),
.C(n_3749),
.Y(n_3980)
);

AOI22xp33_ASAP7_75t_SL g3981 ( 
.A1(n_3891),
.A2(n_3788),
.B1(n_3783),
.B2(n_3818),
.Y(n_3981)
);

AND2x2_ASAP7_75t_SL g3982 ( 
.A(n_3847),
.B(n_3819),
.Y(n_3982)
);

OAI22xp5_ASAP7_75t_L g3983 ( 
.A1(n_3954),
.A2(n_3747),
.B1(n_3818),
.B2(n_3822),
.Y(n_3983)
);

AOI222xp33_ASAP7_75t_L g3984 ( 
.A1(n_3891),
.A2(n_3783),
.B1(n_3829),
.B2(n_3816),
.C1(n_3774),
.C2(n_3827),
.Y(n_3984)
);

AOI221xp5_ASAP7_75t_L g3985 ( 
.A1(n_3891),
.A2(n_3725),
.B1(n_3719),
.B2(n_3722),
.C(n_3730),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3898),
.B(n_3901),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3855),
.Y(n_3987)
);

OAI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3862),
.A2(n_3734),
.B(n_3596),
.Y(n_3988)
);

AOI22xp33_ASAP7_75t_L g3989 ( 
.A1(n_3895),
.A2(n_3788),
.B1(n_3733),
.B2(n_3734),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3842),
.Y(n_3990)
);

OR2x2_ASAP7_75t_L g3991 ( 
.A(n_3946),
.B(n_3788),
.Y(n_3991)
);

AOI22xp33_ASAP7_75t_SL g3992 ( 
.A1(n_3962),
.A2(n_3788),
.B1(n_3576),
.B2(n_3632),
.Y(n_3992)
);

OAI211xp5_ASAP7_75t_SL g3993 ( 
.A1(n_3847),
.A2(n_3788),
.B(n_3795),
.C(n_3576),
.Y(n_3993)
);

AOI22xp33_ASAP7_75t_L g3994 ( 
.A1(n_3895),
.A2(n_3879),
.B1(n_3901),
.B2(n_3889),
.Y(n_3994)
);

OAI221xp5_ASAP7_75t_L g3995 ( 
.A1(n_3942),
.A2(n_3654),
.B1(n_164),
.B2(n_165),
.C(n_166),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3840),
.B(n_3655),
.Y(n_3996)
);

AOI22xp33_ASAP7_75t_L g3997 ( 
.A1(n_3879),
.A2(n_3672),
.B1(n_1562),
.B2(n_1557),
.Y(n_3997)
);

OAI22xp5_ASAP7_75t_L g3998 ( 
.A1(n_3952),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_3998)
);

AOI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_3932),
.A2(n_163),
.B(n_167),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3846),
.Y(n_4000)
);

AND2x4_ASAP7_75t_L g4001 ( 
.A(n_3840),
.B(n_168),
.Y(n_4001)
);

AOI22xp5_ASAP7_75t_L g4002 ( 
.A1(n_3870),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_4002)
);

BUFx2_ASAP7_75t_L g4003 ( 
.A(n_3860),
.Y(n_4003)
);

AOI22xp33_ASAP7_75t_L g4004 ( 
.A1(n_3879),
.A2(n_1490),
.B1(n_1524),
.B2(n_1536),
.Y(n_4004)
);

AOI22xp33_ASAP7_75t_SL g4005 ( 
.A1(n_3956),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_4005)
);

CKINVDCx5p33_ASAP7_75t_R g4006 ( 
.A(n_3893),
.Y(n_4006)
);

NOR2xp33_ASAP7_75t_L g4007 ( 
.A(n_3879),
.B(n_3841),
.Y(n_4007)
);

OAI211xp5_ASAP7_75t_SL g4008 ( 
.A1(n_3947),
.A2(n_174),
.B(n_175),
.C(n_176),
.Y(n_4008)
);

OR2x6_ASAP7_75t_L g4009 ( 
.A(n_3916),
.B(n_176),
.Y(n_4009)
);

AO221x2_ASAP7_75t_L g4010 ( 
.A1(n_3897),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.C(n_181),
.Y(n_4010)
);

AOI22xp33_ASAP7_75t_SL g4011 ( 
.A1(n_3853),
.A2(n_3873),
.B1(n_3917),
.B2(n_3864),
.Y(n_4011)
);

AOI221xp5_ASAP7_75t_L g4012 ( 
.A1(n_3897),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.C(n_182),
.Y(n_4012)
);

INVx3_ASAP7_75t_L g4013 ( 
.A(n_3861),
.Y(n_4013)
);

AOI22xp33_ASAP7_75t_SL g4014 ( 
.A1(n_3853),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_4014)
);

NOR2xp33_ASAP7_75t_SL g4015 ( 
.A(n_3916),
.B(n_187),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3961),
.B(n_188),
.Y(n_4016)
);

BUFx6f_ASAP7_75t_L g4017 ( 
.A(n_3873),
.Y(n_4017)
);

INVx3_ASAP7_75t_L g4018 ( 
.A(n_3861),
.Y(n_4018)
);

AOI21xp5_ASAP7_75t_L g4019 ( 
.A1(n_3889),
.A2(n_189),
.B(n_190),
.Y(n_4019)
);

AND2x4_ASAP7_75t_L g4020 ( 
.A(n_3904),
.B(n_189),
.Y(n_4020)
);

INVx2_ASAP7_75t_L g4021 ( 
.A(n_3918),
.Y(n_4021)
);

OAI211xp5_ASAP7_75t_SL g4022 ( 
.A1(n_3941),
.A2(n_190),
.B(n_192),
.C(n_193),
.Y(n_4022)
);

INVx4_ASAP7_75t_L g4023 ( 
.A(n_3841),
.Y(n_4023)
);

OAI222xp33_ASAP7_75t_L g4024 ( 
.A1(n_3917),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.C1(n_196),
.C2(n_197),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3866),
.Y(n_4025)
);

OAI22xp5_ASAP7_75t_L g4026 ( 
.A1(n_3952),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_4026)
);

AOI221xp5_ASAP7_75t_L g4027 ( 
.A1(n_3909),
.A2(n_198),
.B1(n_202),
.B2(n_203),
.C(n_204),
.Y(n_4027)
);

OAI22xp5_ASAP7_75t_L g4028 ( 
.A1(n_3917),
.A2(n_3889),
.B1(n_3884),
.B2(n_3873),
.Y(n_4028)
);

AOI22xp33_ASAP7_75t_SL g4029 ( 
.A1(n_3861),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_L g4030 ( 
.A1(n_3889),
.A2(n_1524),
.B1(n_1536),
.B2(n_1551),
.Y(n_4030)
);

AOI22xp5_ASAP7_75t_L g4031 ( 
.A1(n_3960),
.A2(n_3900),
.B1(n_3953),
.B2(n_3926),
.Y(n_4031)
);

AOI22xp33_ASAP7_75t_L g4032 ( 
.A1(n_3943),
.A2(n_1524),
.B1(n_1536),
.B2(n_1551),
.Y(n_4032)
);

AOI21x1_ASAP7_75t_L g4033 ( 
.A1(n_3880),
.A2(n_205),
.B(n_206),
.Y(n_4033)
);

AOI221xp5_ASAP7_75t_L g4034 ( 
.A1(n_3911),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.C(n_210),
.Y(n_4034)
);

AOI22xp33_ASAP7_75t_L g4035 ( 
.A1(n_3944),
.A2(n_1536),
.B1(n_1551),
.B2(n_1557),
.Y(n_4035)
);

OAI22xp33_ASAP7_75t_L g4036 ( 
.A1(n_3884),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_4036)
);

CKINVDCx5p33_ASAP7_75t_R g4037 ( 
.A(n_3841),
.Y(n_4037)
);

OAI22xp33_ASAP7_75t_L g4038 ( 
.A1(n_3884),
.A2(n_211),
.B1(n_213),
.B2(n_215),
.Y(n_4038)
);

OAI21xp5_ASAP7_75t_SL g4039 ( 
.A1(n_3864),
.A2(n_211),
.B(n_215),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3896),
.Y(n_4040)
);

OAI211xp5_ASAP7_75t_L g4041 ( 
.A1(n_3859),
.A2(n_216),
.B(n_217),
.C(n_218),
.Y(n_4041)
);

AOI22xp33_ASAP7_75t_L g4042 ( 
.A1(n_3945),
.A2(n_3948),
.B1(n_3951),
.B2(n_3946),
.Y(n_4042)
);

OAI221xp5_ASAP7_75t_L g4043 ( 
.A1(n_3864),
.A2(n_216),
.B1(n_219),
.B2(n_220),
.C(n_221),
.Y(n_4043)
);

AOI22xp33_ASAP7_75t_L g4044 ( 
.A1(n_3951),
.A2(n_1551),
.B1(n_1557),
.B2(n_1562),
.Y(n_4044)
);

OAI21xp33_ASAP7_75t_L g4045 ( 
.A1(n_3892),
.A2(n_219),
.B(n_222),
.Y(n_4045)
);

AOI22xp33_ASAP7_75t_L g4046 ( 
.A1(n_3922),
.A2(n_1562),
.B1(n_1557),
.B2(n_223),
.Y(n_4046)
);

OAI22xp5_ASAP7_75t_L g4047 ( 
.A1(n_3884),
.A2(n_223),
.B1(n_227),
.B2(n_2039),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3923),
.A2(n_3931),
.B1(n_3907),
.B2(n_3859),
.Y(n_4048)
);

AOI22xp33_ASAP7_75t_L g4049 ( 
.A1(n_3882),
.A2(n_1562),
.B1(n_227),
.B2(n_2043),
.Y(n_4049)
);

OAI21xp5_ASAP7_75t_L g4050 ( 
.A1(n_3881),
.A2(n_229),
.B(n_230),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3925),
.B(n_235),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3934),
.B(n_239),
.Y(n_4052)
);

AOI221xp5_ASAP7_75t_L g4053 ( 
.A1(n_3905),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.C(n_245),
.Y(n_4053)
);

AOI22xp33_ASAP7_75t_L g4054 ( 
.A1(n_3882),
.A2(n_2043),
.B1(n_2039),
.B2(n_1478),
.Y(n_4054)
);

NAND4xp25_ASAP7_75t_L g4055 ( 
.A(n_3935),
.B(n_248),
.C(n_249),
.D(n_250),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3938),
.B(n_253),
.Y(n_4056)
);

INVxp67_ASAP7_75t_L g4057 ( 
.A(n_3940),
.Y(n_4057)
);

AO31x2_ASAP7_75t_L g4058 ( 
.A1(n_3913),
.A2(n_255),
.A3(n_256),
.B(n_258),
.Y(n_4058)
);

OAI22xp5_ASAP7_75t_L g4059 ( 
.A1(n_3906),
.A2(n_2043),
.B1(n_2039),
.B2(n_266),
.Y(n_4059)
);

AO22x1_ASAP7_75t_L g4060 ( 
.A1(n_3894),
.A2(n_262),
.B1(n_264),
.B2(n_268),
.Y(n_4060)
);

OAI211xp5_ASAP7_75t_L g4061 ( 
.A1(n_3910),
.A2(n_3899),
.B(n_3921),
.C(n_3915),
.Y(n_4061)
);

AND2x2_ASAP7_75t_L g4062 ( 
.A(n_3925),
.B(n_273),
.Y(n_4062)
);

OAI21xp5_ASAP7_75t_L g4063 ( 
.A1(n_3881),
.A2(n_275),
.B(n_276),
.Y(n_4063)
);

AOI221xp5_ASAP7_75t_L g4064 ( 
.A1(n_3894),
.A2(n_277),
.B1(n_281),
.B2(n_287),
.C(n_289),
.Y(n_4064)
);

INVx11_ASAP7_75t_L g4065 ( 
.A(n_3950),
.Y(n_4065)
);

NAND3xp33_ASAP7_75t_L g4066 ( 
.A(n_3894),
.B(n_2039),
.C(n_2043),
.Y(n_4066)
);

AOI21xp33_ASAP7_75t_SL g4067 ( 
.A1(n_3876),
.A2(n_290),
.B(n_291),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_SL g4068 ( 
.A1(n_3844),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_4068)
);

AOI22xp33_ASAP7_75t_SL g4069 ( 
.A1(n_3844),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3950),
.B(n_301),
.Y(n_4070)
);

AOI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_3844),
.A2(n_302),
.B1(n_303),
.B2(n_305),
.Y(n_4071)
);

AND2x2_ASAP7_75t_L g4072 ( 
.A(n_3957),
.B(n_306),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3845),
.Y(n_4073)
);

CKINVDCx5p33_ASAP7_75t_R g4074 ( 
.A(n_3949),
.Y(n_4074)
);

INVx3_ASAP7_75t_L g4075 ( 
.A(n_3918),
.Y(n_4075)
);

BUFx6f_ASAP7_75t_L g4076 ( 
.A(n_3876),
.Y(n_4076)
);

OAI21x1_ASAP7_75t_L g4077 ( 
.A1(n_3958),
.A2(n_307),
.B(n_312),
.Y(n_4077)
);

OAI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_3949),
.A2(n_3937),
.B1(n_3918),
.B2(n_3957),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3924),
.A2(n_317),
.B1(n_320),
.B2(n_321),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3937),
.Y(n_4080)
);

BUFx3_ASAP7_75t_L g4081 ( 
.A(n_3937),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_4003),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_3986),
.B(n_3966),
.Y(n_4083)
);

INVx2_ASAP7_75t_SL g4084 ( 
.A(n_3965),
.Y(n_4084)
);

BUFx2_ASAP7_75t_L g4085 ( 
.A(n_3963),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_4073),
.Y(n_4086)
);

INVx1_ASAP7_75t_SL g4087 ( 
.A(n_3976),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3977),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_4075),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_4075),
.Y(n_4090)
);

BUFx3_ASAP7_75t_L g4091 ( 
.A(n_4037),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_4033),
.Y(n_4092)
);

AND2x2_ASAP7_75t_L g4093 ( 
.A(n_3974),
.B(n_3927),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3987),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3967),
.B(n_3849),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_3969),
.B(n_3850),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_3981),
.B(n_3927),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_4025),
.Y(n_4098)
);

INVx2_ASAP7_75t_L g4099 ( 
.A(n_3991),
.Y(n_4099)
);

BUFx2_ASAP7_75t_L g4100 ( 
.A(n_4023),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_4001),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_4001),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_4011),
.B(n_3929),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4040),
.Y(n_4104)
);

OR2x2_ASAP7_75t_L g4105 ( 
.A(n_3990),
.B(n_3936),
.Y(n_4105)
);

AND2x2_ASAP7_75t_L g4106 ( 
.A(n_4081),
.B(n_3929),
.Y(n_4106)
);

OR2x2_ASAP7_75t_SL g4107 ( 
.A(n_4017),
.B(n_3913),
.Y(n_4107)
);

AND2x2_ASAP7_75t_L g4108 ( 
.A(n_4013),
.B(n_3930),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_4013),
.B(n_3930),
.Y(n_4109)
);

INVx2_ASAP7_75t_L g4110 ( 
.A(n_4009),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_4018),
.B(n_3933),
.Y(n_4111)
);

OR2x2_ASAP7_75t_SL g4112 ( 
.A(n_4017),
.B(n_3914),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3982),
.B(n_3854),
.Y(n_4113)
);

HB1xp67_ASAP7_75t_L g4114 ( 
.A(n_4009),
.Y(n_4114)
);

OR2x2_ASAP7_75t_L g4115 ( 
.A(n_4000),
.B(n_3936),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_4057),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_3964),
.B(n_3857),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_4031),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4016),
.Y(n_4119)
);

OR2x2_ASAP7_75t_L g4120 ( 
.A(n_4042),
.B(n_3939),
.Y(n_4120)
);

INVx3_ASAP7_75t_L g4121 ( 
.A(n_4023),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_4017),
.Y(n_4122)
);

INVx2_ASAP7_75t_L g4123 ( 
.A(n_4076),
.Y(n_4123)
);

HB1xp67_ASAP7_75t_L g4124 ( 
.A(n_4021),
.Y(n_4124)
);

INVx3_ASAP7_75t_L g4125 ( 
.A(n_4076),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4010),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_4076),
.Y(n_4127)
);

AND2x2_ASAP7_75t_L g4128 ( 
.A(n_4018),
.B(n_3933),
.Y(n_4128)
);

HB1xp67_ASAP7_75t_L g4129 ( 
.A(n_4080),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_3994),
.B(n_3939),
.Y(n_4130)
);

BUFx3_ASAP7_75t_L g4131 ( 
.A(n_4010),
.Y(n_4131)
);

INVx2_ASAP7_75t_L g4132 ( 
.A(n_4020),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_3979),
.B(n_3875),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4052),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4048),
.B(n_3858),
.Y(n_4135)
);

BUFx2_ASAP7_75t_L g4136 ( 
.A(n_4006),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_4056),
.Y(n_4137)
);

BUFx3_ASAP7_75t_L g4138 ( 
.A(n_4007),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4020),
.Y(n_4139)
);

AND2x2_ASAP7_75t_L g4140 ( 
.A(n_3989),
.B(n_3875),
.Y(n_4140)
);

INVx2_ASAP7_75t_L g4141 ( 
.A(n_4077),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4072),
.Y(n_4142)
);

HB1xp67_ASAP7_75t_L g4143 ( 
.A(n_4028),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_4074),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_3984),
.B(n_3885),
.Y(n_4145)
);

NOR2x1_ASAP7_75t_L g4146 ( 
.A(n_4024),
.B(n_3914),
.Y(n_4146)
);

AND2x2_ASAP7_75t_L g4147 ( 
.A(n_3975),
.B(n_3885),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_4065),
.Y(n_4148)
);

HB1xp67_ASAP7_75t_L g4149 ( 
.A(n_4047),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_3980),
.B(n_3869),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_3996),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4061),
.B(n_3863),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_4019),
.B(n_3867),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3998),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_4066),
.Y(n_4155)
);

AND2x4_ASAP7_75t_L g4156 ( 
.A(n_3988),
.B(n_3865),
.Y(n_4156)
);

INVx2_ASAP7_75t_L g4157 ( 
.A(n_4070),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_3970),
.B(n_3869),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_3973),
.B(n_3871),
.Y(n_4159)
);

HB1xp67_ASAP7_75t_L g4160 ( 
.A(n_3983),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4026),
.Y(n_4161)
);

OR2x2_ASAP7_75t_L g4162 ( 
.A(n_3978),
.B(n_3865),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_4051),
.Y(n_4163)
);

OR2x2_ASAP7_75t_L g4164 ( 
.A(n_3972),
.B(n_3843),
.Y(n_4164)
);

BUFx2_ASAP7_75t_L g4165 ( 
.A(n_4050),
.Y(n_4165)
);

BUFx3_ASAP7_75t_L g4166 ( 
.A(n_3968),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4036),
.Y(n_4167)
);

HB1xp67_ASAP7_75t_L g4168 ( 
.A(n_3971),
.Y(n_4168)
);

INVxp67_ASAP7_75t_SL g4169 ( 
.A(n_4038),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_3992),
.B(n_3871),
.Y(n_4170)
);

AND2x2_ASAP7_75t_L g4171 ( 
.A(n_3985),
.B(n_3843),
.Y(n_4171)
);

AND2x2_ASAP7_75t_L g4172 ( 
.A(n_4062),
.B(n_3851),
.Y(n_4172)
);

INVx4_ASAP7_75t_L g4173 ( 
.A(n_4005),
.Y(n_4173)
);

AND2x4_ASAP7_75t_L g4174 ( 
.A(n_4063),
.B(n_3851),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_4131),
.B(n_3999),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_4107),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_4107),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_4083),
.B(n_3852),
.Y(n_4178)
);

HB1xp67_ASAP7_75t_L g4179 ( 
.A(n_4114),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4082),
.Y(n_4180)
);

OR2x2_ASAP7_75t_L g4181 ( 
.A(n_4082),
.B(n_3852),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_4131),
.B(n_4126),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_4082),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_4112),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4101),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_4112),
.Y(n_4186)
);

AOI22xp33_ASAP7_75t_L g4187 ( 
.A1(n_4173),
.A2(n_3993),
.B1(n_4008),
.B2(n_4022),
.Y(n_4187)
);

NOR2xp67_ASAP7_75t_L g4188 ( 
.A(n_4084),
.B(n_4039),
.Y(n_4188)
);

AND2x2_ASAP7_75t_L g4189 ( 
.A(n_4083),
.B(n_3856),
.Y(n_4189)
);

OR2x2_ASAP7_75t_L g4190 ( 
.A(n_4167),
.B(n_3878),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_4085),
.Y(n_4191)
);

AND2x2_ASAP7_75t_L g4192 ( 
.A(n_4085),
.B(n_3856),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4101),
.Y(n_4193)
);

AOI22xp33_ASAP7_75t_L g4194 ( 
.A1(n_4173),
.A2(n_4012),
.B1(n_3995),
.B2(n_4034),
.Y(n_4194)
);

NAND2x1p5_ASAP7_75t_L g4195 ( 
.A(n_4131),
.B(n_4002),
.Y(n_4195)
);

AND2x4_ASAP7_75t_L g4196 ( 
.A(n_4121),
.B(n_3883),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_4100),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_4126),
.B(n_4173),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4101),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_4166),
.B(n_3912),
.Y(n_4200)
);

HB1xp67_ASAP7_75t_L g4201 ( 
.A(n_4102),
.Y(n_4201)
);

OAI22xp5_ASAP7_75t_L g4202 ( 
.A1(n_4173),
.A2(n_4029),
.B1(n_4043),
.B2(n_4014),
.Y(n_4202)
);

INVx3_ASAP7_75t_L g4203 ( 
.A(n_4121),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4102),
.Y(n_4204)
);

AND2x2_ASAP7_75t_L g4205 ( 
.A(n_4166),
.B(n_3890),
.Y(n_4205)
);

AND2x4_ASAP7_75t_L g4206 ( 
.A(n_4121),
.B(n_3949),
.Y(n_4206)
);

INVxp67_ASAP7_75t_SL g4207 ( 
.A(n_4166),
.Y(n_4207)
);

INVx2_ASAP7_75t_L g4208 ( 
.A(n_4100),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4102),
.Y(n_4209)
);

AND2x4_ASAP7_75t_L g4210 ( 
.A(n_4121),
.B(n_4084),
.Y(n_4210)
);

HB1xp67_ASAP7_75t_L g4211 ( 
.A(n_4110),
.Y(n_4211)
);

OR2x2_ASAP7_75t_L g4212 ( 
.A(n_4092),
.B(n_3959),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4105),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_4110),
.B(n_4015),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_SL g4215 ( 
.A(n_4146),
.B(n_4078),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4105),
.Y(n_4216)
);

OR2x2_ASAP7_75t_L g4217 ( 
.A(n_4092),
.B(n_3920),
.Y(n_4217)
);

AND2x4_ASAP7_75t_L g4218 ( 
.A(n_4136),
.B(n_3949),
.Y(n_4218)
);

HB1xp67_ASAP7_75t_L g4219 ( 
.A(n_4110),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4115),
.Y(n_4220)
);

OR2x2_ASAP7_75t_L g4221 ( 
.A(n_4167),
.B(n_4045),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4115),
.Y(n_4222)
);

HB1xp67_ASAP7_75t_L g4223 ( 
.A(n_4132),
.Y(n_4223)
);

NOR2x1_ASAP7_75t_L g4224 ( 
.A(n_4136),
.B(n_4041),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4086),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_4169),
.B(n_4027),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_4089),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4132),
.B(n_4049),
.Y(n_4228)
);

INVx2_ASAP7_75t_L g4229 ( 
.A(n_4203),
.Y(n_4229)
);

INVxp67_ASAP7_75t_L g4230 ( 
.A(n_4207),
.Y(n_4230)
);

INVxp67_ASAP7_75t_SL g4231 ( 
.A(n_4215),
.Y(n_4231)
);

INVx2_ASAP7_75t_L g4232 ( 
.A(n_4203),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_4210),
.B(n_4091),
.Y(n_4233)
);

OR2x2_ASAP7_75t_L g4234 ( 
.A(n_4182),
.B(n_4092),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_4191),
.B(n_4132),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_4203),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4210),
.B(n_4091),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4201),
.Y(n_4238)
);

AND2x4_ASAP7_75t_L g4239 ( 
.A(n_4191),
.B(n_4091),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4210),
.Y(n_4240)
);

HB1xp67_ASAP7_75t_L g4241 ( 
.A(n_4176),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4223),
.Y(n_4242)
);

INVx2_ASAP7_75t_L g4243 ( 
.A(n_4176),
.Y(n_4243)
);

INVx2_ASAP7_75t_SL g4244 ( 
.A(n_4197),
.Y(n_4244)
);

INVx2_ASAP7_75t_SL g4245 ( 
.A(n_4197),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_4179),
.B(n_4159),
.Y(n_4246)
);

BUFx2_ASAP7_75t_L g4247 ( 
.A(n_4208),
.Y(n_4247)
);

AND2x4_ASAP7_75t_L g4248 ( 
.A(n_4208),
.B(n_4138),
.Y(n_4248)
);

OR2x2_ASAP7_75t_L g4249 ( 
.A(n_4198),
.B(n_4095),
.Y(n_4249)
);

BUFx3_ASAP7_75t_L g4250 ( 
.A(n_4180),
.Y(n_4250)
);

OR2x2_ASAP7_75t_L g4251 ( 
.A(n_4211),
.B(n_4095),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4219),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4185),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4193),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4199),
.Y(n_4255)
);

AND2x4_ASAP7_75t_L g4256 ( 
.A(n_4177),
.B(n_4138),
.Y(n_4256)
);

OR2x2_ASAP7_75t_L g4257 ( 
.A(n_4221),
.B(n_4152),
.Y(n_4257)
);

BUFx6f_ASAP7_75t_L g4258 ( 
.A(n_4227),
.Y(n_4258)
);

OR2x2_ASAP7_75t_L g4259 ( 
.A(n_4215),
.B(n_4183),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_4177),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_4184),
.Y(n_4261)
);

AND2x2_ASAP7_75t_L g4262 ( 
.A(n_4178),
.B(n_4159),
.Y(n_4262)
);

OR2x2_ASAP7_75t_L g4263 ( 
.A(n_4204),
.B(n_4152),
.Y(n_4263)
);

INVx3_ASAP7_75t_SL g4264 ( 
.A(n_4218),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4209),
.Y(n_4265)
);

BUFx3_ASAP7_75t_L g4266 ( 
.A(n_4218),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_4187),
.B(n_4139),
.Y(n_4267)
);

AND2x2_ASAP7_75t_L g4268 ( 
.A(n_4178),
.B(n_4138),
.Y(n_4268)
);

INVx3_ASAP7_75t_L g4269 ( 
.A(n_4184),
.Y(n_4269)
);

HB1xp67_ASAP7_75t_L g4270 ( 
.A(n_4186),
.Y(n_4270)
);

INVx4_ASAP7_75t_L g4271 ( 
.A(n_4227),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4187),
.B(n_4139),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4181),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4181),
.Y(n_4274)
);

AND2x4_ASAP7_75t_L g4275 ( 
.A(n_4186),
.B(n_4122),
.Y(n_4275)
);

AND2x2_ASAP7_75t_L g4276 ( 
.A(n_4189),
.B(n_4093),
.Y(n_4276)
);

INVx3_ASAP7_75t_L g4277 ( 
.A(n_4206),
.Y(n_4277)
);

OR2x2_ASAP7_75t_L g4278 ( 
.A(n_4190),
.B(n_4096),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_4189),
.B(n_4093),
.Y(n_4279)
);

INVx3_ASAP7_75t_L g4280 ( 
.A(n_4206),
.Y(n_4280)
);

HB1xp67_ASAP7_75t_L g4281 ( 
.A(n_4240),
.Y(n_4281)
);

INVx2_ASAP7_75t_L g4282 ( 
.A(n_4258),
.Y(n_4282)
);

INVx2_ASAP7_75t_L g4283 ( 
.A(n_4258),
.Y(n_4283)
);

OA211x2_ASAP7_75t_L g4284 ( 
.A1(n_4230),
.A2(n_4194),
.B(n_4175),
.C(n_4214),
.Y(n_4284)
);

OR2x2_ASAP7_75t_L g4285 ( 
.A(n_4259),
.B(n_4096),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4258),
.Y(n_4286)
);

AND2x2_ASAP7_75t_SL g4287 ( 
.A(n_4259),
.B(n_4194),
.Y(n_4287)
);

OR2x2_ASAP7_75t_L g4288 ( 
.A(n_4231),
.B(n_4226),
.Y(n_4288)
);

INVx2_ASAP7_75t_L g4289 ( 
.A(n_4258),
.Y(n_4289)
);

OR2x2_ASAP7_75t_L g4290 ( 
.A(n_4244),
.B(n_4213),
.Y(n_4290)
);

BUFx2_ASAP7_75t_SL g4291 ( 
.A(n_4248),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_4244),
.B(n_4216),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4269),
.Y(n_4293)
);

AND2x2_ASAP7_75t_L g4294 ( 
.A(n_4233),
.B(n_4148),
.Y(n_4294)
);

INVx2_ASAP7_75t_L g4295 ( 
.A(n_4269),
.Y(n_4295)
);

BUFx2_ASAP7_75t_L g4296 ( 
.A(n_4248),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4246),
.B(n_4239),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4247),
.Y(n_4298)
);

NOR2x1_ASAP7_75t_L g4299 ( 
.A(n_4248),
.B(n_4224),
.Y(n_4299)
);

OR2x2_ASAP7_75t_L g4300 ( 
.A(n_4257),
.B(n_4164),
.Y(n_4300)
);

NAND2x1p5_ASAP7_75t_L g4301 ( 
.A(n_4233),
.B(n_4087),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_4269),
.Y(n_4302)
);

INVxp67_ASAP7_75t_L g4303 ( 
.A(n_4246),
.Y(n_4303)
);

OR2x2_ASAP7_75t_L g4304 ( 
.A(n_4257),
.B(n_4164),
.Y(n_4304)
);

OR2x2_ASAP7_75t_L g4305 ( 
.A(n_4245),
.B(n_4220),
.Y(n_4305)
);

HB1xp67_ASAP7_75t_L g4306 ( 
.A(n_4240),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4245),
.Y(n_4307)
);

AND2x2_ASAP7_75t_L g4308 ( 
.A(n_4237),
.B(n_4148),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4237),
.B(n_4148),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_4239),
.B(n_4202),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_4239),
.B(n_4188),
.Y(n_4311)
);

AND2x2_ASAP7_75t_L g4312 ( 
.A(n_4268),
.B(n_4087),
.Y(n_4312)
);

AND2x2_ASAP7_75t_L g4313 ( 
.A(n_4268),
.B(n_4192),
.Y(n_4313)
);

INVxp67_ASAP7_75t_L g4314 ( 
.A(n_4262),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4256),
.B(n_4168),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4262),
.B(n_4192),
.Y(n_4316)
);

OAI22xp5_ASAP7_75t_L g4317 ( 
.A1(n_4278),
.A2(n_4195),
.B1(n_4146),
.B2(n_4165),
.Y(n_4317)
);

HB1xp67_ASAP7_75t_L g4318 ( 
.A(n_4256),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4276),
.B(n_4279),
.Y(n_4319)
);

AND2x2_ASAP7_75t_L g4320 ( 
.A(n_4312),
.B(n_4319),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4312),
.B(n_4276),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_4313),
.B(n_4256),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_L g4323 ( 
.A(n_4313),
.B(n_4279),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4316),
.B(n_4264),
.Y(n_4324)
);

AND2x2_ASAP7_75t_L g4325 ( 
.A(n_4316),
.B(n_4319),
.Y(n_4325)
);

OR2x6_ASAP7_75t_L g4326 ( 
.A(n_4291),
.B(n_4243),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4318),
.Y(n_4327)
);

AOI22xp33_ASAP7_75t_L g4328 ( 
.A1(n_4287),
.A2(n_4160),
.B1(n_4118),
.B2(n_4150),
.Y(n_4328)
);

BUFx2_ASAP7_75t_L g4329 ( 
.A(n_4301),
.Y(n_4329)
);

HB1xp67_ASAP7_75t_L g4330 ( 
.A(n_4299),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4296),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_4294),
.B(n_4144),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4293),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_4294),
.B(n_4252),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_L g4335 ( 
.A(n_4308),
.B(n_4275),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_4308),
.B(n_4275),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4293),
.Y(n_4337)
);

NOR2x1_ASAP7_75t_SL g4338 ( 
.A(n_4290),
.B(n_4266),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4295),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4295),
.Y(n_4340)
);

INVx6_ASAP7_75t_L g4341 ( 
.A(n_4290),
.Y(n_4341)
);

AND2x2_ASAP7_75t_L g4342 ( 
.A(n_4309),
.B(n_4144),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4309),
.B(n_4275),
.Y(n_4343)
);

AND2x2_ASAP7_75t_L g4344 ( 
.A(n_4301),
.B(n_4264),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4303),
.B(n_4241),
.Y(n_4345)
);

NOR3xp33_ASAP7_75t_L g4346 ( 
.A(n_4329),
.B(n_4317),
.C(n_4311),
.Y(n_4346)
);

AND2x2_ASAP7_75t_L g4347 ( 
.A(n_4320),
.B(n_4321),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_4341),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_4321),
.B(n_4314),
.Y(n_4349)
);

AND2x2_ASAP7_75t_L g4350 ( 
.A(n_4325),
.B(n_4298),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4325),
.B(n_4144),
.Y(n_4351)
);

NAND3xp33_ASAP7_75t_SL g4352 ( 
.A(n_4328),
.B(n_4288),
.C(n_4330),
.Y(n_4352)
);

OR2x2_ASAP7_75t_L g4353 ( 
.A(n_4335),
.B(n_4297),
.Y(n_4353)
);

OR2x2_ASAP7_75t_L g4354 ( 
.A(n_4336),
.B(n_4343),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4332),
.B(n_4266),
.Y(n_4355)
);

AND2x2_ASAP7_75t_L g4356 ( 
.A(n_4342),
.B(n_4270),
.Y(n_4356)
);

OR2x2_ASAP7_75t_L g4357 ( 
.A(n_4323),
.B(n_4300),
.Y(n_4357)
);

AND2x2_ASAP7_75t_L g4358 ( 
.A(n_4324),
.B(n_4344),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_4341),
.B(n_4287),
.Y(n_4359)
);

NAND2xp5_ASAP7_75t_SL g4360 ( 
.A(n_4344),
.B(n_4156),
.Y(n_4360)
);

AND2x2_ASAP7_75t_L g4361 ( 
.A(n_4324),
.B(n_4281),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4341),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_4328),
.B(n_4302),
.Y(n_4363)
);

OAI211xp5_ASAP7_75t_L g4364 ( 
.A1(n_4330),
.A2(n_4285),
.B(n_4288),
.C(n_4310),
.Y(n_4364)
);

AND2x4_ASAP7_75t_L g4365 ( 
.A(n_4338),
.B(n_4326),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4365),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_4347),
.B(n_4307),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4361),
.Y(n_4368)
);

NOR3xp33_ASAP7_75t_L g4369 ( 
.A(n_4359),
.B(n_4352),
.C(n_4364),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_4365),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_4355),
.B(n_4331),
.Y(n_4371)
);

AOI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_4358),
.A2(n_4284),
.B1(n_4150),
.B2(n_4118),
.Y(n_4372)
);

AOI221xp5_ASAP7_75t_L g4373 ( 
.A1(n_4352),
.A2(n_4272),
.B1(n_4267),
.B2(n_4117),
.C(n_4285),
.Y(n_4373)
);

A2O1A1Ixp33_ASAP7_75t_L g4374 ( 
.A1(n_4359),
.A2(n_4251),
.B(n_4278),
.C(n_4149),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4356),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4348),
.Y(n_4376)
);

OR2x2_ASAP7_75t_L g4377 ( 
.A(n_4362),
.B(n_4304),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4351),
.Y(n_4378)
);

INVx3_ASAP7_75t_L g4379 ( 
.A(n_4350),
.Y(n_4379)
);

HB1xp67_ASAP7_75t_L g4380 ( 
.A(n_4349),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4357),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4353),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4379),
.Y(n_4383)
);

OR2x2_ASAP7_75t_L g4384 ( 
.A(n_4379),
.B(n_4326),
.Y(n_4384)
);

OR2x2_ASAP7_75t_L g4385 ( 
.A(n_4366),
.B(n_4326),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_4380),
.B(n_4345),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4377),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4370),
.B(n_4243),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_L g4389 ( 
.A(n_4369),
.B(n_4302),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_4367),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4378),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_4368),
.B(n_4260),
.Y(n_4392)
);

OR2x2_ASAP7_75t_L g4393 ( 
.A(n_4371),
.B(n_4322),
.Y(n_4393)
);

AND2x2_ASAP7_75t_L g4394 ( 
.A(n_4375),
.B(n_4345),
.Y(n_4394)
);

AND2x2_ASAP7_75t_L g4395 ( 
.A(n_4394),
.B(n_4327),
.Y(n_4395)
);

AND2x4_ASAP7_75t_L g4396 ( 
.A(n_4386),
.B(n_4306),
.Y(n_4396)
);

INVx1_ASAP7_75t_SL g4397 ( 
.A(n_4384),
.Y(n_4397)
);

INVx1_ASAP7_75t_SL g4398 ( 
.A(n_4385),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4388),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_4387),
.B(n_4260),
.Y(n_4400)
);

AOI22xp33_ASAP7_75t_L g4401 ( 
.A1(n_4390),
.A2(n_4373),
.B1(n_4143),
.B2(n_4346),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4383),
.B(n_4261),
.Y(n_4402)
);

NOR2xp33_ASAP7_75t_L g4403 ( 
.A(n_4396),
.B(n_4360),
.Y(n_4403)
);

NAND3xp33_ASAP7_75t_SL g4404 ( 
.A(n_4401),
.B(n_4364),
.C(n_4363),
.Y(n_4404)
);

OAI221xp5_ASAP7_75t_SL g4405 ( 
.A1(n_4397),
.A2(n_4372),
.B1(n_4249),
.B2(n_4251),
.C(n_4374),
.Y(n_4405)
);

OAI221xp5_ASAP7_75t_L g4406 ( 
.A1(n_4400),
.A2(n_4363),
.B1(n_4315),
.B2(n_4389),
.C(n_4235),
.Y(n_4406)
);

AOI22xp5_ASAP7_75t_L g4407 ( 
.A1(n_4398),
.A2(n_4381),
.B1(n_4376),
.B2(n_4382),
.Y(n_4407)
);

NOR2xp33_ASAP7_75t_L g4408 ( 
.A(n_4396),
.B(n_4334),
.Y(n_4408)
);

O2A1O1Ixp5_ASAP7_75t_L g4409 ( 
.A1(n_4395),
.A2(n_4271),
.B(n_4283),
.C(n_4289),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4402),
.Y(n_4410)
);

OAI21xp5_ASAP7_75t_SL g4411 ( 
.A1(n_4399),
.A2(n_4242),
.B(n_4238),
.Y(n_4411)
);

AOI21xp33_ASAP7_75t_SL g4412 ( 
.A1(n_4396),
.A2(n_4389),
.B(n_4305),
.Y(n_4412)
);

AOI22xp5_ASAP7_75t_L g4413 ( 
.A1(n_4397),
.A2(n_4261),
.B1(n_4277),
.B2(n_4280),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_4396),
.B(n_4250),
.Y(n_4414)
);

AND2x2_ASAP7_75t_L g4415 ( 
.A(n_4395),
.B(n_4391),
.Y(n_4415)
);

AOI22xp33_ASAP7_75t_L g4416 ( 
.A1(n_4404),
.A2(n_4218),
.B1(n_4280),
.B2(n_4277),
.Y(n_4416)
);

INVx2_ASAP7_75t_SL g4417 ( 
.A(n_4414),
.Y(n_4417)
);

OAI21xp33_ASAP7_75t_L g4418 ( 
.A1(n_4413),
.A2(n_4392),
.B(n_4354),
.Y(n_4418)
);

INVxp67_ASAP7_75t_L g4419 ( 
.A(n_4403),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4409),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_4412),
.B(n_4333),
.Y(n_4421)
);

BUFx2_ASAP7_75t_L g4422 ( 
.A(n_4415),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_4410),
.Y(n_4423)
);

O2A1O1Ixp33_ASAP7_75t_SL g4424 ( 
.A1(n_4408),
.A2(n_4286),
.B(n_4283),
.C(n_4282),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_4407),
.B(n_4337),
.Y(n_4425)
);

AOI22xp33_ASAP7_75t_L g4426 ( 
.A1(n_4406),
.A2(n_4280),
.B1(n_4277),
.B2(n_4250),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4411),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_4405),
.B(n_4339),
.Y(n_4428)
);

INVxp67_ASAP7_75t_SL g4429 ( 
.A(n_4413),
.Y(n_4429)
);

NAND2xp5_ASAP7_75t_L g4430 ( 
.A(n_4413),
.B(n_4340),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_4413),
.Y(n_4431)
);

OAI22xp33_ASAP7_75t_SL g4432 ( 
.A1(n_4405),
.A2(n_4305),
.B1(n_4292),
.B2(n_4234),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_4409),
.Y(n_4433)
);

OAI22xp5_ASAP7_75t_L g4434 ( 
.A1(n_4413),
.A2(n_4249),
.B1(n_4234),
.B2(n_4292),
.Y(n_4434)
);

AND2x2_ASAP7_75t_SL g4435 ( 
.A(n_4403),
.B(n_4393),
.Y(n_4435)
);

NOR2xp33_ASAP7_75t_L g4436 ( 
.A(n_4413),
.B(n_4282),
.Y(n_4436)
);

OAI22xp5_ASAP7_75t_L g4437 ( 
.A1(n_4413),
.A2(n_4263),
.B1(n_4228),
.B2(n_4116),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4416),
.B(n_4289),
.Y(n_4438)
);

INVx1_ASAP7_75t_L g4439 ( 
.A(n_4434),
.Y(n_4439)
);

INVx1_ASAP7_75t_SL g4440 ( 
.A(n_4422),
.Y(n_4440)
);

NOR2xp33_ASAP7_75t_L g4441 ( 
.A(n_4432),
.B(n_4263),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4424),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_4426),
.B(n_4273),
.Y(n_4443)
);

AND2x2_ASAP7_75t_L g4444 ( 
.A(n_4435),
.B(n_4205),
.Y(n_4444)
);

AOI221xp5_ASAP7_75t_L g4445 ( 
.A1(n_4437),
.A2(n_4253),
.B1(n_4254),
.B2(n_4265),
.C(n_4255),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_4436),
.B(n_4274),
.Y(n_4446)
);

NOR2xp33_ASAP7_75t_L g4447 ( 
.A(n_4418),
.B(n_4271),
.Y(n_4447)
);

INVxp67_ASAP7_75t_L g4448 ( 
.A(n_4421),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4429),
.B(n_4205),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_4418),
.B(n_4195),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_4423),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4431),
.B(n_4116),
.Y(n_4452)
);

OR2x2_ASAP7_75t_L g4453 ( 
.A(n_4425),
.B(n_4222),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4430),
.Y(n_4454)
);

AND2x2_ASAP7_75t_L g4455 ( 
.A(n_4419),
.B(n_4200),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_4417),
.B(n_4200),
.Y(n_4456)
);

AOI22xp5_ASAP7_75t_L g4457 ( 
.A1(n_4420),
.A2(n_4271),
.B1(n_4236),
.B2(n_4232),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_4433),
.B(n_4119),
.Y(n_4458)
);

OR2x2_ASAP7_75t_L g4459 ( 
.A(n_4428),
.B(n_4088),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4427),
.B(n_4119),
.Y(n_4460)
);

NOR2xp33_ASAP7_75t_L g4461 ( 
.A(n_4432),
.B(n_4229),
.Y(n_4461)
);

AOI22xp33_ASAP7_75t_L g4462 ( 
.A1(n_4422),
.A2(n_4125),
.B1(n_4232),
.B2(n_4229),
.Y(n_4462)
);

BUFx4f_ASAP7_75t_SL g4463 ( 
.A(n_4422),
.Y(n_4463)
);

INVx4_ASAP7_75t_L g4464 ( 
.A(n_4463),
.Y(n_4464)
);

OR2x2_ASAP7_75t_L g4465 ( 
.A(n_4450),
.B(n_4088),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4444),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_4449),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4456),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_L g4469 ( 
.A(n_4462),
.B(n_4236),
.Y(n_4469)
);

NOR2xp33_ASAP7_75t_L g4470 ( 
.A(n_4438),
.B(n_4225),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4457),
.Y(n_4471)
);

INVx2_ASAP7_75t_L g4472 ( 
.A(n_4455),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4457),
.Y(n_4473)
);

XNOR2xp5_ASAP7_75t_L g4474 ( 
.A(n_4440),
.B(n_4154),
.Y(n_4474)
);

OR2x2_ASAP7_75t_L g4475 ( 
.A(n_4446),
.B(n_4094),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4461),
.Y(n_4476)
);

AOI22xp5_ASAP7_75t_L g4477 ( 
.A1(n_4441),
.A2(n_4122),
.B1(n_4127),
.B2(n_4123),
.Y(n_4477)
);

OR2x2_ASAP7_75t_L g4478 ( 
.A(n_4443),
.B(n_4094),
.Y(n_4478)
);

INVxp67_ASAP7_75t_SL g4479 ( 
.A(n_4447),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4442),
.B(n_4098),
.Y(n_4480)
);

XNOR2x2_ASAP7_75t_SL g4481 ( 
.A(n_4453),
.B(n_4212),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_4445),
.B(n_4098),
.Y(n_4482)
);

XNOR2xp5_ASAP7_75t_L g4483 ( 
.A(n_4439),
.B(n_4154),
.Y(n_4483)
);

INVxp67_ASAP7_75t_L g4484 ( 
.A(n_4452),
.Y(n_4484)
);

OR2x2_ASAP7_75t_L g4485 ( 
.A(n_4459),
.B(n_4104),
.Y(n_4485)
);

INVx1_ASAP7_75t_SL g4486 ( 
.A(n_4458),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4451),
.Y(n_4487)
);

NOR3xp33_ASAP7_75t_L g4488 ( 
.A(n_4464),
.B(n_4448),
.C(n_4454),
.Y(n_4488)
);

OAI211xp5_ASAP7_75t_SL g4489 ( 
.A1(n_4476),
.A2(n_4460),
.B(n_4217),
.C(n_4123),
.Y(n_4489)
);

NOR3xp33_ASAP7_75t_L g4490 ( 
.A(n_4464),
.B(n_4125),
.C(n_4123),
.Y(n_4490)
);

AO22x2_ASAP7_75t_L g4491 ( 
.A1(n_4467),
.A2(n_4127),
.B1(n_4125),
.B2(n_4122),
.Y(n_4491)
);

NOR2x1_ASAP7_75t_L g4492 ( 
.A(n_4480),
.B(n_4125),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_4481),
.Y(n_4493)
);

NAND2xp33_ASAP7_75t_SL g4494 ( 
.A(n_4474),
.B(n_4483),
.Y(n_4494)
);

AOI21xp5_ASAP7_75t_L g4495 ( 
.A1(n_4482),
.A2(n_4127),
.B(n_4212),
.Y(n_4495)
);

INVx1_ASAP7_75t_L g4496 ( 
.A(n_4477),
.Y(n_4496)
);

OAI21xp33_ASAP7_75t_L g4497 ( 
.A1(n_4468),
.A2(n_4206),
.B(n_4217),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_4466),
.B(n_4104),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4472),
.B(n_4103),
.Y(n_4499)
);

OR2x2_ASAP7_75t_L g4500 ( 
.A(n_4469),
.B(n_4465),
.Y(n_4500)
);

OAI211xp5_ASAP7_75t_SL g4501 ( 
.A1(n_4487),
.A2(n_4161),
.B(n_4113),
.C(n_4135),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4471),
.B(n_4196),
.Y(n_4502)
);

NOR4xp25_ASAP7_75t_L g4503 ( 
.A(n_4473),
.B(n_4089),
.C(n_4090),
.D(n_4086),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4479),
.B(n_4103),
.Y(n_4504)
);

OAI21xp33_ASAP7_75t_L g4505 ( 
.A1(n_4499),
.A2(n_4470),
.B(n_4486),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4504),
.Y(n_4506)
);

INVx2_ASAP7_75t_L g4507 ( 
.A(n_4491),
.Y(n_4507)
);

OAI21xp5_ASAP7_75t_L g4508 ( 
.A1(n_4497),
.A2(n_4484),
.B(n_4478),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4502),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4491),
.Y(n_4510)
);

AOI221xp5_ASAP7_75t_L g4511 ( 
.A1(n_4503),
.A2(n_4475),
.B1(n_4485),
.B2(n_4196),
.C(n_4156),
.Y(n_4511)
);

INVx2_ASAP7_75t_SL g4512 ( 
.A(n_4492),
.Y(n_4512)
);

OAI32xp33_ASAP7_75t_L g4513 ( 
.A1(n_4490),
.A2(n_4089),
.A3(n_4090),
.B1(n_4099),
.B2(n_4124),
.Y(n_4513)
);

NOR2xp33_ASAP7_75t_R g4514 ( 
.A(n_4494),
.B(n_4134),
.Y(n_4514)
);

OAI22xp5_ASAP7_75t_L g4515 ( 
.A1(n_4493),
.A2(n_4196),
.B1(n_4162),
.B2(n_4090),
.Y(n_4515)
);

A2O1A1Ixp33_ASAP7_75t_L g4516 ( 
.A1(n_4495),
.A2(n_4156),
.B(n_4145),
.C(n_4158),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4496),
.B(n_4161),
.Y(n_4517)
);

OAI211xp5_ASAP7_75t_L g4518 ( 
.A1(n_4498),
.A2(n_4145),
.B(n_4129),
.C(n_4099),
.Y(n_4518)
);

OAI311xp33_ASAP7_75t_L g4519 ( 
.A1(n_4500),
.A2(n_4135),
.A3(n_4162),
.B1(n_4120),
.C1(n_4153),
.Y(n_4519)
);

OAI221xp5_ASAP7_75t_SL g4520 ( 
.A1(n_4511),
.A2(n_4488),
.B1(n_4489),
.B2(n_4501),
.C(n_4099),
.Y(n_4520)
);

NAND4xp25_ASAP7_75t_L g4521 ( 
.A(n_4517),
.B(n_4158),
.C(n_4156),
.D(n_4130),
.Y(n_4521)
);

O2A1O1Ixp33_ASAP7_75t_L g4522 ( 
.A1(n_4512),
.A2(n_4120),
.B(n_4165),
.C(n_4151),
.Y(n_4522)
);

OAI221xp5_ASAP7_75t_L g4523 ( 
.A1(n_4515),
.A2(n_4151),
.B1(n_4130),
.B2(n_4155),
.C(n_4153),
.Y(n_4523)
);

AOI22xp5_ASAP7_75t_L g4524 ( 
.A1(n_4506),
.A2(n_4170),
.B1(n_4097),
.B2(n_4147),
.Y(n_4524)
);

AOI211xp5_ASAP7_75t_L g4525 ( 
.A1(n_4505),
.A2(n_4508),
.B(n_4509),
.C(n_4513),
.Y(n_4525)
);

AOI211xp5_ASAP7_75t_L g4526 ( 
.A1(n_4519),
.A2(n_4097),
.B(n_4170),
.C(n_4147),
.Y(n_4526)
);

NAND4xp25_ASAP7_75t_L g4527 ( 
.A(n_4516),
.B(n_4140),
.C(n_4151),
.D(n_4171),
.Y(n_4527)
);

AOI221xp5_ASAP7_75t_L g4528 ( 
.A1(n_4514),
.A2(n_4140),
.B1(n_4171),
.B2(n_4155),
.C(n_4137),
.Y(n_4528)
);

O2A1O1Ixp33_ASAP7_75t_L g4529 ( 
.A1(n_4510),
.A2(n_4141),
.B(n_4155),
.C(n_4134),
.Y(n_4529)
);

A2O1A1Ixp33_ASAP7_75t_L g4530 ( 
.A1(n_4507),
.A2(n_4518),
.B(n_4137),
.C(n_4106),
.Y(n_4530)
);

NAND3xp33_ASAP7_75t_L g4531 ( 
.A(n_4506),
.B(n_4106),
.C(n_4108),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4515),
.Y(n_4532)
);

AOI221xp5_ASAP7_75t_L g4533 ( 
.A1(n_4515),
.A2(n_4128),
.B1(n_4108),
.B2(n_4109),
.C(n_4111),
.Y(n_4533)
);

AOI21xp33_ASAP7_75t_L g4534 ( 
.A1(n_4506),
.A2(n_4142),
.B(n_4141),
.Y(n_4534)
);

AOI211xp5_ASAP7_75t_SL g4535 ( 
.A1(n_4505),
.A2(n_4141),
.B(n_4109),
.C(n_4128),
.Y(n_4535)
);

NOR3xp33_ASAP7_75t_L g4536 ( 
.A(n_4505),
.B(n_4142),
.C(n_4163),
.Y(n_4536)
);

AOI322xp5_ASAP7_75t_L g4537 ( 
.A1(n_4506),
.A2(n_4111),
.A3(n_4174),
.B1(n_4163),
.B2(n_4157),
.C1(n_4133),
.C2(n_4172),
.Y(n_4537)
);

NOR3x2_ASAP7_75t_L g4538 ( 
.A(n_4525),
.B(n_4174),
.C(n_4163),
.Y(n_4538)
);

OAI211xp5_ASAP7_75t_SL g4539 ( 
.A1(n_4532),
.A2(n_4157),
.B(n_4064),
.C(n_4053),
.Y(n_4539)
);

OR2x2_ASAP7_75t_L g4540 ( 
.A(n_4521),
.B(n_4157),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4531),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_4535),
.B(n_4174),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4529),
.Y(n_4543)
);

NOR2x1_ASAP7_75t_L g4544 ( 
.A(n_4530),
.B(n_4174),
.Y(n_4544)
);

NAND4xp75_ASAP7_75t_L g4545 ( 
.A(n_4534),
.B(n_4133),
.C(n_4172),
.D(n_3920),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4536),
.B(n_3874),
.Y(n_4546)
);

NOR2x1_ASAP7_75t_L g4547 ( 
.A(n_4522),
.B(n_4055),
.Y(n_4547)
);

NOR2x1_ASAP7_75t_L g4548 ( 
.A(n_4527),
.B(n_4059),
.Y(n_4548)
);

NAND3xp33_ASAP7_75t_SL g4549 ( 
.A(n_4526),
.B(n_4067),
.C(n_4068),
.Y(n_4549)
);

NOR3xp33_ASAP7_75t_L g4550 ( 
.A(n_4520),
.B(n_4060),
.C(n_4069),
.Y(n_4550)
);

NAND3xp33_ASAP7_75t_SL g4551 ( 
.A(n_4524),
.B(n_4030),
.C(n_4046),
.Y(n_4551)
);

INVx1_ASAP7_75t_SL g4552 ( 
.A(n_4523),
.Y(n_4552)
);

NOR3x1_ASAP7_75t_L g4553 ( 
.A(n_4528),
.B(n_3874),
.C(n_3958),
.Y(n_4553)
);

XNOR2x1_ASAP7_75t_L g4554 ( 
.A(n_4537),
.B(n_322),
.Y(n_4554)
);

AOI21x1_ASAP7_75t_L g4555 ( 
.A1(n_4543),
.A2(n_4533),
.B(n_326),
.Y(n_4555)
);

NAND4xp25_ASAP7_75t_SL g4556 ( 
.A(n_4544),
.B(n_4054),
.C(n_4071),
.D(n_4004),
.Y(n_4556)
);

NOR2x1_ASAP7_75t_L g4557 ( 
.A(n_4541),
.B(n_325),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4538),
.Y(n_4558)
);

AOI211xp5_ASAP7_75t_L g4559 ( 
.A1(n_4552),
.A2(n_327),
.B(n_330),
.C(n_331),
.Y(n_4559)
);

NAND4xp25_ASAP7_75t_L g4560 ( 
.A(n_4540),
.B(n_4079),
.C(n_4035),
.D(n_4032),
.Y(n_4560)
);

OAI211xp5_ASAP7_75t_SL g4561 ( 
.A1(n_4542),
.A2(n_333),
.B(n_336),
.C(n_339),
.Y(n_4561)
);

A2O1A1Ixp33_ASAP7_75t_L g4562 ( 
.A1(n_4548),
.A2(n_4044),
.B(n_3997),
.C(n_3887),
.Y(n_4562)
);

NOR4xp25_ASAP7_75t_L g4563 ( 
.A(n_4546),
.B(n_343),
.C(n_344),
.D(n_345),
.Y(n_4563)
);

NAND4xp25_ASAP7_75t_L g4564 ( 
.A(n_4547),
.B(n_347),
.C(n_350),
.D(n_351),
.Y(n_4564)
);

OAI221xp5_ASAP7_75t_L g4565 ( 
.A1(n_4554),
.A2(n_4058),
.B1(n_354),
.B2(n_358),
.C(n_359),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_4557),
.B(n_4550),
.Y(n_4566)
);

NAND2xp33_ASAP7_75t_L g4567 ( 
.A(n_4558),
.B(n_4545),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4563),
.B(n_4549),
.Y(n_4568)
);

NOR2xp33_ASAP7_75t_L g4569 ( 
.A(n_4555),
.B(n_4551),
.Y(n_4569)
);

AOI22xp5_ASAP7_75t_L g4570 ( 
.A1(n_4565),
.A2(n_4539),
.B1(n_4553),
.B2(n_3887),
.Y(n_4570)
);

NOR2xp67_ASAP7_75t_L g4571 ( 
.A(n_4564),
.B(n_353),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_L g4572 ( 
.A(n_4571),
.B(n_4570),
.Y(n_4572)
);

OR2x2_ASAP7_75t_L g4573 ( 
.A(n_4568),
.B(n_4556),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4566),
.Y(n_4574)
);

NOR2xp33_ASAP7_75t_L g4575 ( 
.A(n_4574),
.B(n_4567),
.Y(n_4575)
);

NOR2xp67_ASAP7_75t_L g4576 ( 
.A(n_4573),
.B(n_4569),
.Y(n_4576)
);

AOI22xp5_ASAP7_75t_L g4577 ( 
.A1(n_4575),
.A2(n_4561),
.B1(n_4572),
.B2(n_4559),
.Y(n_4577)
);

XNOR2x2_ASAP7_75t_L g4578 ( 
.A(n_4577),
.B(n_4576),
.Y(n_4578)
);

AOI22xp5_ASAP7_75t_L g4579 ( 
.A1(n_4578),
.A2(n_4560),
.B1(n_4562),
.B2(n_366),
.Y(n_4579)
);

OR2x2_ASAP7_75t_L g4580 ( 
.A(n_4579),
.B(n_361),
.Y(n_4580)
);

NOR3xp33_ASAP7_75t_L g4581 ( 
.A(n_4580),
.B(n_363),
.C(n_369),
.Y(n_4581)
);

AND2x2_ASAP7_75t_SL g4582 ( 
.A(n_4581),
.B(n_372),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4582),
.Y(n_4583)
);

NAND3xp33_ASAP7_75t_L g4584 ( 
.A(n_4583),
.B(n_1554),
.C(n_383),
.Y(n_4584)
);

XOR2xp5_ASAP7_75t_L g4585 ( 
.A(n_4584),
.B(n_379),
.Y(n_4585)
);

OAI21xp5_ASAP7_75t_L g4586 ( 
.A1(n_4585),
.A2(n_1554),
.B(n_384),
.Y(n_4586)
);

INVx3_ASAP7_75t_L g4587 ( 
.A(n_4586),
.Y(n_4587)
);

OAI22xp5_ASAP7_75t_L g4588 ( 
.A1(n_4587),
.A2(n_1554),
.B1(n_395),
.B2(n_396),
.Y(n_4588)
);

OAI221xp5_ASAP7_75t_R g4589 ( 
.A1(n_4588),
.A2(n_389),
.B1(n_399),
.B2(n_402),
.C(n_403),
.Y(n_4589)
);

AOI22xp5_ASAP7_75t_L g4590 ( 
.A1(n_4589),
.A2(n_404),
.B1(n_405),
.B2(n_406),
.Y(n_4590)
);

AOI211xp5_ASAP7_75t_L g4591 ( 
.A1(n_4590),
.A2(n_408),
.B(n_409),
.C(n_413),
.Y(n_4591)
);


endmodule