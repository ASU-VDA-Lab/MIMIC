module real_aes_6333_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_717;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g259 ( .A1(n_0), .A2(n_260), .B(n_261), .C(n_264), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_1), .B(n_201), .Y(n_265) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_3), .B(n_171), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_4), .A2(n_141), .B(n_144), .C(n_451), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_5), .A2(n_161), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_6), .A2(n_161), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_7), .B(n_201), .Y(n_497) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_8), .A2(n_128), .B(n_181), .Y(n_180) );
AND2x6_ASAP7_75t_L g141 ( .A(n_9), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_10), .A2(n_141), .B(n_144), .C(n_147), .Y(n_143) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_11), .A2(n_44), .B1(n_115), .B2(n_116), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_11), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_12), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_12), .B(n_40), .Y(n_439) );
INVx1_ASAP7_75t_L g467 ( .A(n_13), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_14), .B(n_151), .Y(n_453) );
INVx1_ASAP7_75t_L g133 ( .A(n_15), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_16), .B(n_171), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_17), .A2(n_149), .B(n_475), .C(n_477), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_18), .B(n_201), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_19), .B(n_225), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_20), .A2(n_144), .B(n_188), .C(n_221), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_21), .A2(n_153), .B(n_263), .C(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_22), .B(n_151), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_23), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_24), .B(n_151), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_25), .Y(n_525) );
INVx1_ASAP7_75t_L g517 ( .A(n_26), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_27), .A2(n_144), .B(n_184), .C(n_188), .Y(n_183) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_28), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_29), .Y(n_449) );
INVx1_ASAP7_75t_L g508 ( .A(n_30), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_31), .A2(n_161), .B(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g139 ( .A(n_32), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_33), .A2(n_163), .B(n_174), .C(n_209), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_34), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_35), .A2(n_263), .B(n_494), .C(n_496), .Y(n_493) );
INVxp67_ASAP7_75t_L g509 ( .A(n_36), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_37), .B(n_186), .Y(n_185) );
CKINVDCx14_ASAP7_75t_R g492 ( .A(n_38), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_39), .A2(n_144), .B(n_188), .C(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g111 ( .A(n_40), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_41), .A2(n_264), .B(n_465), .C(n_466), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_42), .B(n_219), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_43), .Y(n_156) );
INVx1_ASAP7_75t_L g116 ( .A(n_44), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_45), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_46), .B(n_161), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_47), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_48), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_49), .A2(n_163), .B(n_165), .C(n_174), .Y(n_162) );
INVx1_ASAP7_75t_L g262 ( .A(n_50), .Y(n_262) );
INVx1_ASAP7_75t_L g166 ( .A(n_51), .Y(n_166) );
INVx1_ASAP7_75t_L g482 ( .A(n_52), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_53), .B(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_54), .A2(n_58), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_54), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_55), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_56), .Y(n_228) );
CKINVDCx14_ASAP7_75t_R g463 ( .A(n_57), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_58), .Y(n_731) );
INVx1_ASAP7_75t_L g142 ( .A(n_59), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_60), .B(n_161), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_61), .B(n_201), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_62), .A2(n_195), .B(n_197), .C(n_199), .Y(n_194) );
INVx1_ASAP7_75t_L g132 ( .A(n_63), .Y(n_132) );
INVx1_ASAP7_75t_SL g495 ( .A(n_64), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_65), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_66), .B(n_171), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_67), .B(n_201), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_68), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g528 ( .A(n_69), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_70), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_71), .B(n_168), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_72), .A2(n_144), .B(n_174), .C(n_235), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_73), .Y(n_193) );
INVx1_ASAP7_75t_L g108 ( .A(n_74), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_75), .A2(n_161), .B(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_76), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_77), .A2(n_161), .B(n_472), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_78), .A2(n_219), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g473 ( .A(n_79), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_80), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_81), .B(n_167), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_82), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_83), .A2(n_161), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g476 ( .A(n_84), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_85), .A2(n_102), .B1(n_112), .B2(n_742), .Y(n_101) );
INVx2_ASAP7_75t_L g130 ( .A(n_86), .Y(n_130) );
INVx1_ASAP7_75t_L g452 ( .A(n_87), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_88), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_89), .B(n_151), .Y(n_150) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_90), .B(n_105), .C(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g437 ( .A(n_90), .B(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g709 ( .A(n_90), .Y(n_709) );
OR2x2_ASAP7_75t_L g735 ( .A(n_90), .B(n_722), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_91), .A2(n_144), .B(n_174), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_92), .B(n_161), .Y(n_207) );
INVx1_ASAP7_75t_L g210 ( .A(n_93), .Y(n_210) );
INVxp67_ASAP7_75t_L g198 ( .A(n_94), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_95), .B(n_128), .Y(n_468) );
INVx2_ASAP7_75t_L g485 ( .A(n_96), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_97), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
INVx1_ASAP7_75t_L g236 ( .A(n_99), .Y(n_236) );
AND2x2_ASAP7_75t_L g177 ( .A(n_100), .B(n_176), .Y(n_177) );
INVx5_ASAP7_75t_SL g742 ( .A(n_102), .Y(n_742) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_109), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g438 ( .A(n_105), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AO221x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_723), .B1(n_726), .B2(n_736), .C(n_738), .Y(n_112) );
OAI222xp33_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_117), .B1(n_710), .B2(n_711), .C1(n_717), .C2(n_718), .Y(n_113) );
INVx1_ASAP7_75t_L g710 ( .A(n_114), .Y(n_710) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_435), .B1(n_440), .B2(n_706), .Y(n_118) );
INVx2_ASAP7_75t_L g714 ( .A(n_119), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_119), .A2(n_714), .B1(n_729), .B2(n_730), .Y(n_728) );
OR3x1_ASAP7_75t_L g119 ( .A(n_120), .B(n_333), .C(n_398), .Y(n_119) );
NAND4xp25_ASAP7_75t_SL g120 ( .A(n_121), .B(n_274), .C(n_300), .D(n_323), .Y(n_120) );
AOI221xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_202), .B1(n_243), .B2(n_250), .C(n_266), .Y(n_121) );
CKINVDCx14_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_123), .A2(n_267), .B1(n_291), .B2(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_178), .Y(n_123) );
INVx1_ASAP7_75t_SL g327 ( .A(n_124), .Y(n_327) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_158), .Y(n_124) );
OR2x2_ASAP7_75t_L g248 ( .A(n_125), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g269 ( .A(n_125), .B(n_179), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_125), .B(n_189), .Y(n_282) );
AND2x2_ASAP7_75t_L g299 ( .A(n_125), .B(n_158), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_125), .B(n_246), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_125), .B(n_298), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_125), .B(n_178), .Y(n_420) );
AOI211xp5_ASAP7_75t_SL g431 ( .A1(n_125), .A2(n_337), .B(n_432), .C(n_433), .Y(n_431) );
INVx5_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_126), .B(n_179), .Y(n_303) );
AND2x2_ASAP7_75t_L g306 ( .A(n_126), .B(n_180), .Y(n_306) );
OR2x2_ASAP7_75t_L g351 ( .A(n_126), .B(n_179), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_126), .B(n_189), .Y(n_360) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_134), .B(n_155), .Y(n_126) );
INVx3_ASAP7_75t_L g201 ( .A(n_127), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_127), .B(n_213), .Y(n_212) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_127), .A2(n_233), .B(n_241), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_127), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_127), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_127), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_127), .A2(n_524), .B(n_530), .Y(n_523) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_128), .A2(n_182), .B(n_183), .Y(n_181) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_128), .Y(n_190) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g157 ( .A(n_129), .Y(n_157) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_130), .B(n_131), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_136), .B(n_143), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_136), .A2(n_449), .B(n_450), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_136), .A2(n_176), .B(n_514), .C(n_515), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_136), .A2(n_525), .B(n_526), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
AND2x4_ASAP7_75t_L g161 ( .A(n_137), .B(n_141), .Y(n_161) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx1_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
INVx1_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx3_ASAP7_75t_L g149 ( .A(n_140), .Y(n_149) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
INVx1_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
INVx4_ASAP7_75t_SL g175 ( .A(n_141), .Y(n_175) );
BUFx3_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
INVx5_ASAP7_75t_L g164 ( .A(n_144), .Y(n_164) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx3_ASAP7_75t_L g173 ( .A(n_145), .Y(n_173) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_145), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_150), .B(n_152), .Y(n_147) );
INVx5_ASAP7_75t_L g171 ( .A(n_149), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_149), .B(n_467), .Y(n_466) );
INVx4_ASAP7_75t_L g263 ( .A(n_151), .Y(n_263) );
INVx2_ASAP7_75t_L g465 ( .A(n_151), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_152), .A2(n_185), .B(n_187), .Y(n_184) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx2_ASAP7_75t_L g502 ( .A(n_157), .Y(n_502) );
INVx5_ASAP7_75t_SL g249 ( .A(n_158), .Y(n_249) );
AND2x2_ASAP7_75t_L g268 ( .A(n_158), .B(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_158), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g354 ( .A(n_158), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g386 ( .A(n_158), .B(n_189), .Y(n_386) );
OR2x2_ASAP7_75t_L g392 ( .A(n_158), .B(n_282), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_158), .B(n_342), .Y(n_401) );
OR2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_177), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_176), .Y(n_159) );
BUFx2_ASAP7_75t_L g219 ( .A(n_161), .Y(n_219) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_164), .A2(n_175), .B(n_193), .C(n_194), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_164), .A2(n_175), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g462 ( .A1(n_164), .A2(n_175), .B(n_463), .C(n_464), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_SL g472 ( .A1(n_164), .A2(n_175), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_164), .A2(n_175), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_164), .A2(n_175), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_164), .A2(n_175), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_170), .C(n_172), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g209 ( .A1(n_167), .A2(n_172), .B(n_210), .C(n_211), .Y(n_209) );
O2A1O1Ixp5_ASAP7_75t_L g451 ( .A1(n_167), .A2(n_452), .B(n_453), .C(n_454), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_167), .A2(n_454), .B(n_528), .C(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx4_ASAP7_75t_L g196 ( .A(n_169), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_171), .B(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g260 ( .A(n_171), .Y(n_260) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_171), .A2(n_196), .B1(n_508), .B2(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_171), .A2(n_224), .B(n_517), .C(n_518), .Y(n_516) );
HB1xp67_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g264 ( .A(n_173), .Y(n_264) );
INVx1_ASAP7_75t_L g477 ( .A(n_173), .Y(n_477) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_176), .A2(n_207), .B(n_208), .Y(n_206) );
INVx2_ASAP7_75t_L g226 ( .A(n_176), .Y(n_226) );
INVx1_ASAP7_75t_L g229 ( .A(n_176), .Y(n_229) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_176), .A2(n_461), .B(n_468), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_189), .Y(n_178) );
AND2x2_ASAP7_75t_L g283 ( .A(n_179), .B(n_249), .Y(n_283) );
INVx1_ASAP7_75t_SL g296 ( .A(n_179), .Y(n_296) );
OR2x2_ASAP7_75t_L g331 ( .A(n_179), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g337 ( .A(n_179), .B(n_189), .Y(n_337) );
AND2x2_ASAP7_75t_L g395 ( .A(n_179), .B(n_246), .Y(n_395) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_180), .B(n_249), .Y(n_322) );
INVx3_ASAP7_75t_L g246 ( .A(n_189), .Y(n_246) );
OR2x2_ASAP7_75t_L g288 ( .A(n_189), .B(n_249), .Y(n_288) );
AND2x2_ASAP7_75t_L g298 ( .A(n_189), .B(n_296), .Y(n_298) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_189), .Y(n_346) );
AND2x2_ASAP7_75t_L g355 ( .A(n_189), .B(n_269), .Y(n_355) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_200), .Y(n_189) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_190), .A2(n_471), .B(n_478), .Y(n_470) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_190), .A2(n_480), .B(n_486), .Y(n_479) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_190), .A2(n_490), .B(n_497), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_195), .A2(n_236), .B(n_237), .C(n_238), .Y(n_235) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_196), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_196), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g224 ( .A(n_199), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_199), .B(n_507), .Y(n_506) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_201), .A2(n_256), .B(n_265), .Y(n_255) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_202), .A2(n_372), .B1(n_374), .B2(n_376), .C(n_379), .Y(n_371) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
AND2x2_ASAP7_75t_L g345 ( .A(n_204), .B(n_326), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_204), .B(n_404), .Y(n_408) );
OR2x2_ASAP7_75t_L g429 ( .A(n_204), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_204), .B(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx5_ASAP7_75t_L g276 ( .A(n_205), .Y(n_276) );
AND2x2_ASAP7_75t_L g353 ( .A(n_205), .B(n_216), .Y(n_353) );
AND2x2_ASAP7_75t_L g414 ( .A(n_205), .B(n_293), .Y(n_414) );
AND2x2_ASAP7_75t_L g427 ( .A(n_205), .B(n_246), .Y(n_427) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_212), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_230), .Y(n_214) );
AND2x4_ASAP7_75t_L g253 ( .A(n_215), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g272 ( .A(n_215), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g279 ( .A(n_215), .Y(n_279) );
AND2x2_ASAP7_75t_L g348 ( .A(n_215), .B(n_326), .Y(n_348) );
AND2x2_ASAP7_75t_L g358 ( .A(n_215), .B(n_276), .Y(n_358) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_215), .Y(n_366) );
AND2x2_ASAP7_75t_L g378 ( .A(n_215), .B(n_255), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_215), .B(n_310), .Y(n_382) );
AND2x2_ASAP7_75t_L g419 ( .A(n_215), .B(n_414), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_215), .B(n_293), .Y(n_430) );
OR2x2_ASAP7_75t_L g432 ( .A(n_215), .B(n_368), .Y(n_432) );
INVx5_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g318 ( .A(n_216), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g328 ( .A(n_216), .B(n_273), .Y(n_328) );
AND2x2_ASAP7_75t_L g340 ( .A(n_216), .B(n_255), .Y(n_340) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_216), .Y(n_370) );
AND2x4_ASAP7_75t_L g404 ( .A(n_216), .B(n_254), .Y(n_404) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_227), .Y(n_216) );
AOI21xp5_ASAP7_75t_SL g217 ( .A1(n_218), .A2(n_220), .B(n_225), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_226), .B(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
AO21x2_ASAP7_75t_L g447 ( .A1(n_229), .A2(n_448), .B(n_455), .Y(n_447) );
BUFx2_ASAP7_75t_L g252 ( .A(n_230), .Y(n_252) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g293 ( .A(n_231), .Y(n_293) );
AND2x2_ASAP7_75t_L g326 ( .A(n_231), .B(n_255), .Y(n_326) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g273 ( .A(n_232), .B(n_255), .Y(n_273) );
BUFx2_ASAP7_75t_L g319 ( .A(n_232), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx3_ASAP7_75t_L g496 ( .A(n_239), .Y(n_496) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_245), .B(n_327), .Y(n_406) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_246), .B(n_269), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_246), .B(n_249), .Y(n_308) );
AND2x2_ASAP7_75t_L g363 ( .A(n_246), .B(n_299), .Y(n_363) );
AOI221xp5_ASAP7_75t_SL g300 ( .A1(n_247), .A2(n_301), .B1(n_309), .B2(n_311), .C(n_315), .Y(n_300) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g295 ( .A(n_248), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g336 ( .A(n_248), .B(n_337), .Y(n_336) );
OAI321xp33_ASAP7_75t_L g343 ( .A1(n_248), .A2(n_302), .A3(n_344), .B1(n_346), .B2(n_347), .C(n_349), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_249), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_252), .B(n_404), .Y(n_422) );
AND2x2_ASAP7_75t_L g309 ( .A(n_253), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_253), .B(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_254), .Y(n_285) );
AND2x2_ASAP7_75t_L g292 ( .A(n_254), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_254), .B(n_367), .Y(n_397) );
INVx1_ASAP7_75t_L g434 ( .A(n_254), .Y(n_434) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_263), .B(n_495), .Y(n_494) );
INVx2_ASAP7_75t_L g454 ( .A(n_264), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .B(n_271), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g426 ( .A1(n_268), .A2(n_378), .B(n_427), .C(n_428), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_269), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_269), .B(n_307), .Y(n_373) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g316 ( .A(n_273), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_273), .B(n_276), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_273), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_273), .B(n_358), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_277), .B1(n_289), .B2(n_294), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g290 ( .A(n_276), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g313 ( .A(n_276), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g325 ( .A(n_276), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_276), .B(n_319), .Y(n_361) );
OR2x2_ASAP7_75t_L g368 ( .A(n_276), .B(n_293), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_276), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g418 ( .A(n_276), .B(n_404), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .B1(n_284), .B2(n_286), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g324 ( .A(n_279), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_282), .A2(n_297), .B1(n_365), .B2(n_369), .Y(n_364) );
INVx1_ASAP7_75t_L g412 ( .A(n_283), .Y(n_412) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_287), .A2(n_324), .B1(n_327), .B2(n_328), .C(n_329), .Y(n_323) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g302 ( .A(n_288), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_292), .B(n_358), .Y(n_390) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_293), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_293), .Y(n_314) );
NAND2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g332 ( .A(n_299), .Y(n_332) );
AND2x2_ASAP7_75t_L g341 ( .A(n_299), .B(n_342), .Y(n_341) );
NAND2xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x2_ASAP7_75t_L g385 ( .A(n_306), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_309), .A2(n_335), .B1(n_338), .B2(n_341), .C(n_343), .Y(n_334) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_313), .B(n_370), .Y(n_369) );
AOI21xp33_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_317), .B(n_320), .Y(n_315) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_320), .Y(n_417) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
OR2x2_ASAP7_75t_L g359 ( .A(n_322), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g380 ( .A(n_325), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_325), .B(n_385), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_328), .B(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND4xp25_ASAP7_75t_L g333 ( .A(n_334), .B(n_352), .C(n_371), .D(n_384), .Y(n_333) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g342 ( .A(n_337), .Y(n_342) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g375 ( .A(n_346), .B(n_351), .Y(n_375) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI211xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B(n_356), .C(n_364), .Y(n_352) );
AOI211xp5_ASAP7_75t_L g423 ( .A1(n_354), .A2(n_396), .B(n_424), .C(n_431), .Y(n_423) );
INVx1_ASAP7_75t_SL g383 ( .A(n_355), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B1(n_361), .B2(n_362), .Y(n_356) );
INVx1_ASAP7_75t_L g387 ( .A(n_361), .Y(n_387) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_367), .B(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_367), .B(n_378), .Y(n_411) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g388 ( .A(n_378), .Y(n_388) );
AOI21xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B(n_383), .Y(n_379) );
INVxp33_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI322xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .A3(n_388), .B1(n_389), .B2(n_391), .C1(n_393), .C2(n_396), .Y(n_384) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND3xp33_ASAP7_75t_SL g398 ( .A(n_399), .B(n_416), .C(n_423), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B1(n_405), .B2(n_407), .C(n_409), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g415 ( .A(n_404), .Y(n_415) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_412), .B2(n_413), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_419), .B2(n_420), .C(n_421), .Y(n_416) );
NAND2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g713 ( .A(n_436), .Y(n_713) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g708 ( .A(n_438), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g722 ( .A(n_438), .Y(n_722) );
INVx2_ASAP7_75t_L g715 ( .A(n_440), .Y(n_715) );
OR2x2_ASAP7_75t_SL g440 ( .A(n_441), .B(n_661), .Y(n_440) );
NAND5xp2_ASAP7_75t_L g441 ( .A(n_442), .B(n_573), .C(n_611), .D(n_632), .E(n_649), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_545), .C(n_566), .Y(n_442) );
OAI221xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_487), .B1(n_511), .B2(n_532), .C(n_536), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_457), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_446), .B(n_534), .Y(n_553) );
OR2x2_ASAP7_75t_L g580 ( .A(n_446), .B(n_470), .Y(n_580) );
AND2x2_ASAP7_75t_L g594 ( .A(n_446), .B(n_470), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_446), .B(n_460), .Y(n_608) );
AND2x2_ASAP7_75t_L g646 ( .A(n_446), .B(n_610), .Y(n_646) );
AND2x2_ASAP7_75t_L g675 ( .A(n_446), .B(n_585), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_446), .B(n_557), .Y(n_692) );
INVx4_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g572 ( .A(n_447), .B(n_469), .Y(n_572) );
BUFx3_ASAP7_75t_L g597 ( .A(n_447), .Y(n_597) );
AND2x2_ASAP7_75t_L g626 ( .A(n_447), .B(n_470), .Y(n_626) );
AND3x2_ASAP7_75t_L g639 ( .A(n_447), .B(n_640), .C(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g562 ( .A(n_457), .Y(n_562) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_469), .Y(n_457) );
AOI32xp33_ASAP7_75t_L g617 ( .A1(n_458), .A2(n_569), .A3(n_618), .B1(n_621), .B2(n_622), .Y(n_617) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g544 ( .A(n_459), .B(n_469), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_459), .B(n_572), .Y(n_615) );
AND2x2_ASAP7_75t_L g622 ( .A(n_459), .B(n_594), .Y(n_622) );
OR2x2_ASAP7_75t_L g628 ( .A(n_459), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_459), .B(n_583), .Y(n_653) );
OR2x2_ASAP7_75t_L g671 ( .A(n_459), .B(n_499), .Y(n_671) );
BUFx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g535 ( .A(n_460), .B(n_479), .Y(n_535) );
INVx2_ASAP7_75t_L g557 ( .A(n_460), .Y(n_557) );
OR2x2_ASAP7_75t_L g579 ( .A(n_460), .B(n_479), .Y(n_579) );
AND2x2_ASAP7_75t_L g584 ( .A(n_460), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_460), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g640 ( .A(n_460), .B(n_534), .Y(n_640) );
INVx1_ASAP7_75t_SL g691 ( .A(n_469), .Y(n_691) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
INVx1_ASAP7_75t_SL g534 ( .A(n_470), .Y(n_534) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_470), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_470), .B(n_620), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_470), .B(n_557), .C(n_675), .Y(n_686) );
INVx2_ASAP7_75t_L g585 ( .A(n_479), .Y(n_585) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_479), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_488), .B(n_498), .Y(n_487) );
INVx1_ASAP7_75t_L g621 ( .A(n_488), .Y(n_621) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g539 ( .A(n_489), .B(n_522), .Y(n_539) );
INVx2_ASAP7_75t_L g556 ( .A(n_489), .Y(n_556) );
AND2x2_ASAP7_75t_L g561 ( .A(n_489), .B(n_523), .Y(n_561) );
AND2x2_ASAP7_75t_L g576 ( .A(n_489), .B(n_512), .Y(n_576) );
AND2x2_ASAP7_75t_L g588 ( .A(n_489), .B(n_560), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_498), .B(n_604), .Y(n_603) );
NAND2x1p5_ASAP7_75t_L g660 ( .A(n_498), .B(n_561), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_498), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_498), .B(n_555), .Y(n_683) );
BUFx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g521 ( .A(n_499), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_499), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g565 ( .A(n_499), .B(n_512), .Y(n_565) );
AND2x2_ASAP7_75t_L g591 ( .A(n_499), .B(n_522), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_499), .B(n_631), .Y(n_630) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_503), .B(n_510), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_501), .A2(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g550 ( .A(n_503), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_510), .Y(n_551) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_512), .B(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g555 ( .A(n_512), .B(n_556), .Y(n_555) );
INVx3_ASAP7_75t_SL g560 ( .A(n_512), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_512), .B(n_547), .Y(n_613) );
OR2x2_ASAP7_75t_L g623 ( .A(n_512), .B(n_549), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_512), .B(n_591), .Y(n_651) );
OR2x2_ASAP7_75t_L g681 ( .A(n_512), .B(n_522), .Y(n_681) );
AND2x2_ASAP7_75t_L g685 ( .A(n_512), .B(n_523), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_512), .B(n_561), .Y(n_698) );
AND2x2_ASAP7_75t_L g705 ( .A(n_512), .B(n_587), .Y(n_705) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_519), .Y(n_512) );
INVx1_ASAP7_75t_SL g648 ( .A(n_521), .Y(n_648) );
AND2x2_ASAP7_75t_L g587 ( .A(n_522), .B(n_549), .Y(n_587) );
AND2x2_ASAP7_75t_L g601 ( .A(n_522), .B(n_556), .Y(n_601) );
AND2x2_ASAP7_75t_L g604 ( .A(n_522), .B(n_560), .Y(n_604) );
INVx1_ASAP7_75t_L g631 ( .A(n_522), .Y(n_631) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
BUFx2_ASAP7_75t_L g543 ( .A(n_523), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_533), .A2(n_579), .B(n_703), .C(n_704), .Y(n_702) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g609 ( .A(n_534), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_535), .B(n_552), .Y(n_567) );
AND2x2_ASAP7_75t_L g593 ( .A(n_535), .B(n_594), .Y(n_593) );
OAI21xp5_ASAP7_75t_SL g536 ( .A1(n_537), .A2(n_540), .B(n_544), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_538), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g564 ( .A(n_539), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_539), .B(n_560), .Y(n_605) );
AND2x2_ASAP7_75t_L g696 ( .A(n_539), .B(n_547), .Y(n_696) );
INVxp67_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g569 ( .A(n_543), .B(n_556), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_543), .B(n_554), .Y(n_570) );
OAI322xp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_553), .A3(n_554), .B1(n_557), .B2(n_558), .C1(n_562), .C2(n_563), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_552), .Y(n_546) );
AND2x2_ASAP7_75t_L g657 ( .A(n_547), .B(n_569), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_547), .B(n_621), .Y(n_703) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g600 ( .A(n_549), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g666 ( .A(n_553), .B(n_579), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_554), .B(n_648), .Y(n_647) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_555), .B(n_587), .Y(n_644) );
AND2x2_ASAP7_75t_L g590 ( .A(n_556), .B(n_560), .Y(n_590) );
AND2x2_ASAP7_75t_L g598 ( .A(n_557), .B(n_599), .Y(n_598) );
A2O1A1Ixp33_ASAP7_75t_L g695 ( .A1(n_557), .A2(n_636), .B(n_696), .C(n_697), .Y(n_695) );
AOI21xp33_ASAP7_75t_L g668 ( .A1(n_558), .A2(n_571), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_560), .B(n_587), .Y(n_627) );
AND2x2_ASAP7_75t_L g633 ( .A(n_560), .B(n_601), .Y(n_633) );
AND2x2_ASAP7_75t_L g667 ( .A(n_560), .B(n_569), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_561), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_SL g677 ( .A(n_561), .Y(n_677) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_565), .A2(n_593), .B1(n_595), .B2(n_600), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g566 ( .A1(n_567), .A2(n_568), .B1(n_570), .B2(n_571), .Y(n_566) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_567), .A2(n_603), .B1(n_605), .B2(n_606), .Y(n_602) );
INVxp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_572), .A2(n_674), .B1(n_676), .B2(n_678), .C(n_682), .Y(n_673) );
AOI211xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_577), .B(n_581), .C(n_602), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OR2x2_ASAP7_75t_L g643 ( .A(n_579), .B(n_596), .Y(n_643) );
INVx1_ASAP7_75t_L g694 ( .A(n_579), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g581 ( .A1(n_580), .A2(n_582), .B1(n_586), .B2(n_589), .C(n_592), .Y(n_581) );
INVx2_ASAP7_75t_SL g636 ( .A(n_580), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g701 ( .A(n_583), .Y(n_701) );
AND2x2_ASAP7_75t_L g625 ( .A(n_584), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g610 ( .A(n_585), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g672 ( .A(n_588), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_596), .B(n_698), .Y(n_697) );
CKINVDCx16_ASAP7_75t_R g596 ( .A(n_597), .Y(n_596) );
INVxp67_ASAP7_75t_L g641 ( .A(n_599), .Y(n_641) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_600), .A2(n_612), .B(n_614), .C(n_616), .Y(n_611) );
INVx1_ASAP7_75t_L g689 ( .A(n_603), .Y(n_689) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_607), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx2_ASAP7_75t_L g620 ( .A(n_610), .Y(n_620) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI222xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_623), .B1(n_624), .B2(n_627), .C1(n_628), .C2(n_630), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g656 ( .A(n_620), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_623), .B(n_677), .Y(n_676) );
NAND2xp33_ASAP7_75t_SL g654 ( .A(n_624), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g629 ( .A(n_626), .Y(n_629) );
AND2x2_ASAP7_75t_L g693 ( .A(n_626), .B(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g659 ( .A(n_629), .B(n_656), .Y(n_659) );
INVx1_ASAP7_75t_L g688 ( .A(n_630), .Y(n_688) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_637), .C(n_642), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_636), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
AOI322xp5_ASAP7_75t_L g687 ( .A1(n_639), .A2(n_667), .A3(n_672), .B1(n_688), .B2(n_689), .C1(n_690), .C2(n_693), .Y(n_687) );
AND2x2_ASAP7_75t_L g674 ( .A(n_640), .B(n_675), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B1(n_645), .B2(n_647), .Y(n_642) );
INVxp33_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B1(n_654), .B2(n_657), .C(n_658), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND5xp2_ASAP7_75t_L g661 ( .A(n_662), .B(n_673), .C(n_687), .D(n_695), .E(n_699), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_667), .B(n_668), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVxp33_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_675), .A2(n_700), .B(n_701), .C(n_702), .Y(n_699) );
AOI31xp33_ASAP7_75t_L g682 ( .A1(n_677), .A2(n_683), .A3(n_684), .B(n_686), .Y(n_682) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g700 ( .A(n_698), .Y(n_700) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g716 ( .A(n_707), .Y(n_716) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR2x2_ASAP7_75t_L g721 ( .A(n_709), .B(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
OAI22x1_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_712) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
BUFx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g737 ( .A(n_725), .Y(n_737) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_728), .B(n_733), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g741 ( .A(n_735), .Y(n_741) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
endmodule