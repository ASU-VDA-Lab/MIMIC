module fake_jpeg_14629_n_43 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_43);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_43;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx11_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_12),
.A2(n_1),
.B1(n_7),
.B2(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_4),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_30),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.C(n_25),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_19),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_8),
.B1(n_15),
.B2(n_13),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_23),
.B1(n_24),
.B2(n_2),
.Y(n_31)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_0),
.Y(n_36)
);

OAI22x1_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_19),
.B1(n_20),
.B2(n_10),
.Y(n_33)
);

A2O1A1O1Ixp25_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_37),
.B(n_38),
.C(n_32),
.D(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_37),
.B(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_5),
.B(n_11),
.Y(n_42)
);

AOI221xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_1),
.B1(n_3),
.B2(n_18),
.C(n_23),
.Y(n_43)
);


endmodule