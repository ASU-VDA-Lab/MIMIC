module fake_jpeg_30412_n_360 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_360);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_60),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_49),
.B(n_34),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_22),
.B(n_10),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_10),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_65),
.Y(n_72)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_15),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_67),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_75),
.B(n_89),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_79),
.B(n_82),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_32),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_27),
.B1(n_36),
.B2(n_40),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_83),
.A2(n_107),
.B1(n_41),
.B2(n_39),
.Y(n_131)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_28),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_37),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_37),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_93),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_44),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_95),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_96),
.A2(n_103),
.B1(n_67),
.B2(n_36),
.Y(n_126)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_42),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_111),
.B(n_72),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_26),
.B1(n_33),
.B2(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_29),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_61),
.A2(n_27),
.B1(n_36),
.B2(n_39),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_48),
.B(n_38),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_59),
.B(n_38),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

AO22x2_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_41),
.B1(n_39),
.B2(n_36),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_118),
.A2(n_147),
.A3(n_153),
.B1(n_122),
.B2(n_130),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_78),
.B(n_2),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_86),
.C(n_76),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_103),
.B1(n_86),
.B2(n_109),
.Y(n_157)
);

NOR2x1_ASAP7_75t_R g184 ( 
.A(n_127),
.B(n_34),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_70),
.B1(n_76),
.B2(n_115),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_20),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_68),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_107),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_144),
.B(n_2),
.Y(n_187)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_84),
.A2(n_26),
.B1(n_33),
.B2(n_23),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_146),
.B1(n_150),
.B2(n_113),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_35),
.B1(n_34),
.B2(n_13),
.Y(n_144)
);

BUFx6f_ASAP7_75t_SL g145 ( 
.A(n_112),
.Y(n_145)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_67),
.B1(n_41),
.B2(n_39),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_83),
.A2(n_34),
.B1(n_41),
.B2(n_25),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_88),
.A2(n_35),
.B1(n_34),
.B2(n_25),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_163),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_155),
.B(n_159),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_169),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_120),
.A2(n_87),
.B1(n_91),
.B2(n_69),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_183),
.B1(n_185),
.B2(n_118),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_105),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_160),
.Y(n_215)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_73),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_162),
.B(n_80),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_130),
.B1(n_147),
.B2(n_124),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_105),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_180),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_115),
.B1(n_77),
.B2(n_97),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_141),
.B(n_134),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_184),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_70),
.B1(n_77),
.B2(n_91),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_118),
.B1(n_100),
.B2(n_119),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_118),
.B1(n_133),
.B2(n_125),
.Y(n_201)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_117),
.C(n_134),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_178),
.C(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_105),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_179),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_112),
.C(n_71),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_34),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_71),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_92),
.C(n_80),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_131),
.A2(n_147),
.B1(n_118),
.B2(n_152),
.Y(n_183)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_187),
.A2(n_8),
.B(n_9),
.Y(n_222)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_100),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_136),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_191),
.A2(n_218),
.B1(n_220),
.B2(n_174),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_124),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_194),
.B(n_195),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_190),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_198),
.B(n_210),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_199),
.B(n_206),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_200),
.A2(n_201),
.B1(n_207),
.B2(n_225),
.Y(n_243)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_177),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_169),
.A2(n_133),
.B1(n_125),
.B2(n_92),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_3),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_176),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_211),
.B(n_213),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_175),
.B(n_12),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_219),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_25),
.B1(n_11),
.B2(n_6),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_172),
.B(n_3),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_11),
.B1(n_6),
.B2(n_8),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_176),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_221),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_222),
.A2(n_165),
.B(n_182),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_170),
.B(n_156),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_226),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_149),
.B1(n_8),
.B2(n_9),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_5),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_178),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_251),
.C(n_223),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_228),
.A2(n_225),
.B1(n_203),
.B2(n_199),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_157),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_244),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_223),
.B(n_208),
.Y(n_256)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_238),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_170),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_165),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_239),
.B(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_197),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_242),
.Y(n_274)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_201),
.A2(n_158),
.B1(n_156),
.B2(n_171),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_191),
.B1(n_243),
.B2(n_218),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_188),
.C(n_186),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_198),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_255),
.B(n_258),
.C(n_262),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_261),
.B(n_220),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_223),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_208),
.B(n_207),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_206),
.C(n_219),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_192),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_265),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_206),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_253),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_211),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_247),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_267),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_228),
.B1(n_209),
.B2(n_222),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_206),
.C(n_192),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_275),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_243),
.B1(n_249),
.B2(n_203),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_194),
.Y(n_275)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_210),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_278),
.C(n_236),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_214),
.C(n_213),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_263),
.Y(n_299)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_282),
.Y(n_300)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_275),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_258),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_259),
.B1(n_271),
.B2(n_250),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_292),
.B1(n_212),
.B2(n_254),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_230),
.B(n_248),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_290),
.A2(n_297),
.B(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_266),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_295),
.B(n_221),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_231),
.B1(n_235),
.B2(n_234),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_296),
.A2(n_257),
.B1(n_274),
.B2(n_264),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_231),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_299),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_308),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_310),
.B1(n_311),
.B2(n_297),
.Y(n_314)
);

OA21x2_ASAP7_75t_SL g305 ( 
.A1(n_284),
.A2(n_278),
.B(n_255),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_307),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_262),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_281),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_292),
.A2(n_274),
.B1(n_233),
.B2(n_240),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_290),
.A2(n_241),
.B(n_242),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_282),
.B(n_279),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_314),
.A2(n_320),
.B1(n_325),
.B2(n_326),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_237),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_301),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_317),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_283),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_318),
.A2(n_313),
.B1(n_304),
.B2(n_301),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_291),
.C(n_286),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_323),
.C(n_299),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_300),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_291),
.C(n_296),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_280),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_195),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_327),
.B(n_334),
.C(n_336),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_331),
.B(n_315),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_332),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_322),
.A2(n_309),
.B(n_313),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_SL g332 ( 
.A1(n_318),
.A2(n_288),
.A3(n_302),
.B1(n_310),
.B2(n_312),
.C1(n_297),
.C2(n_306),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_294),
.C(n_281),
.Y(n_334)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_244),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_321),
.C(n_316),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_316),
.C(n_314),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_338),
.B(n_340),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_328),
.Y(n_346)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_333),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_343),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_181),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_334),
.A2(n_161),
.B(n_9),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_344),
.B(n_345),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_335),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_14),
.Y(n_353)
);

FAx1_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_329),
.CI(n_336),
.CON(n_347),
.SN(n_347)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_347),
.A2(n_14),
.B1(n_15),
.B2(n_5),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_181),
.C(n_11),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_350),
.B(n_343),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_352),
.B(n_353),
.C(n_354),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_353),
.A2(n_351),
.B(n_347),
.Y(n_355)
);

OAI21x1_ASAP7_75t_SL g357 ( 
.A1(n_355),
.A2(n_348),
.B(n_349),
.Y(n_357)
);

AOI21x1_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_348),
.B(n_356),
.Y(n_358)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_358),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_14),
.Y(n_360)
);


endmodule