module fake_netlist_1_9628_n_608 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_608);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_608;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_67;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_70;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_68;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g67 ( .A(n_6), .Y(n_67) );
CKINVDCx5p33_ASAP7_75t_R g68 ( .A(n_29), .Y(n_68) );
INVxp33_ASAP7_75t_L g69 ( .A(n_17), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_43), .Y(n_70) );
CKINVDCx20_ASAP7_75t_R g71 ( .A(n_66), .Y(n_71) );
INVxp67_ASAP7_75t_SL g72 ( .A(n_37), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_51), .Y(n_73) );
INVx1_ASAP7_75t_SL g74 ( .A(n_65), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_8), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_62), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_64), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_12), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_41), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_53), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_60), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_61), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_45), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_63), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_57), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_34), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_32), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_54), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_55), .Y(n_89) );
NOR2xp67_ASAP7_75t_L g90 ( .A(n_0), .B(n_31), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_35), .Y(n_91) );
INVxp67_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_27), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_28), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_22), .Y(n_95) );
BUFx10_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_44), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_10), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_52), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_12), .Y(n_100) );
HB1xp67_ASAP7_75t_L g101 ( .A(n_56), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_33), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_42), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_30), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_19), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
BUFx2_ASAP7_75t_SL g107 ( .A(n_16), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_49), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_58), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_48), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_16), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_96), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_70), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_70), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_78), .B(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_73), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_71), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_77), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_93), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_111), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_111), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_96), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_93), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_96), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_96), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_67), .B(n_1), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_103), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_84), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_101), .B(n_1), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_107), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_92), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_94), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_107), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_68), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_76), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_103), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_81), .B(n_2), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_82), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_82), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_69), .B(n_2), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_110), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_67), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_83), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_74), .Y(n_150) );
OAI22xp5_ASAP7_75t_SL g151 ( .A1(n_98), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_83), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_147), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_147), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_112), .B(n_91), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_147), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_118), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_130), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_130), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_130), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_112), .B(n_86), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_130), .Y(n_166) );
NAND3x1_ASAP7_75t_L g167 ( .A(n_115), .B(n_75), .C(n_100), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_130), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_130), .Y(n_169) );
NOR2xp33_ASAP7_75t_R g170 ( .A(n_123), .B(n_110), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_112), .B(n_109), .Y(n_171) );
AO22x2_ASAP7_75t_L g172 ( .A1(n_128), .A2(n_109), .B1(n_108), .B2(n_85), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_112), .B(n_108), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
BUFx2_ASAP7_75t_L g175 ( .A(n_125), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_125), .B(n_97), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
NOR3xp33_ASAP7_75t_L g178 ( .A(n_151), .B(n_106), .C(n_105), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_133), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
NAND2x1p5_ASAP7_75t_L g182 ( .A(n_128), .B(n_99), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_133), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_125), .B(n_106), .Y(n_184) );
INVx8_ASAP7_75t_L g185 ( .A(n_125), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_148), .B(n_105), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_133), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_128), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_128), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_124), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_124), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_124), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_148), .B(n_75), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_129), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_129), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_129), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_142), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_113), .B(n_104), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_142), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_113), .B(n_104), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_114), .B(n_100), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_114), .A2(n_89), .B1(n_99), .B2(n_97), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_142), .Y(n_204) );
INVx4_ASAP7_75t_L g205 ( .A(n_185), .Y(n_205) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_194), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_157), .B(n_134), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_165), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_172), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_194), .B(n_140), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_157), .B(n_134), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_185), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_170), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_175), .B(n_141), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_194), .B(n_150), .Y(n_217) );
BUFx4f_ASAP7_75t_L g218 ( .A(n_182), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_175), .B(n_132), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_182), .A2(n_139), .B1(n_122), .B2(n_121), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_194), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_193), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_172), .A2(n_149), .B1(n_119), .B2(n_117), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_184), .B(n_149), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_181), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_184), .B(n_119), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_160), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_181), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_184), .B(n_131), .Y(n_229) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_171), .A2(n_117), .B(n_116), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_184), .B(n_137), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_193), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_172), .Y(n_233) );
BUFx2_ASAP7_75t_L g234 ( .A(n_172), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_182), .Y(n_235) );
NOR3xp33_ASAP7_75t_SL g236 ( .A(n_199), .B(n_136), .C(n_146), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_202), .B(n_116), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_167), .A2(n_178), .B1(n_202), .B2(n_189), .Y(n_238) );
NAND3xp33_ASAP7_75t_SL g239 ( .A(n_203), .B(n_126), .C(n_143), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_193), .Y(n_240) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_167), .A2(n_144), .B1(n_138), .B2(n_137), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_202), .B(n_144), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
AOI211xp5_ASAP7_75t_L g244 ( .A1(n_187), .A2(n_138), .B(n_135), .C(n_127), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_186), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_193), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_193), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_185), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_187), .B(n_135), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_189), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_185), .Y(n_251) );
NOR2xp33_ASAP7_75t_R g252 ( .A(n_185), .B(n_127), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_193), .Y(n_253) );
NOR3xp33_ASAP7_75t_SL g254 ( .A(n_201), .B(n_72), .C(n_80), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_202), .B(n_145), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_164), .B(n_145), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_173), .Y(n_257) );
BUFx10_ASAP7_75t_L g258 ( .A(n_186), .Y(n_258) );
NAND3xp33_ASAP7_75t_L g259 ( .A(n_189), .B(n_120), .C(n_102), .Y(n_259) );
NOR3xp33_ASAP7_75t_SL g260 ( .A(n_176), .B(n_85), .C(n_87), .Y(n_260) );
INVxp67_ASAP7_75t_SL g261 ( .A(n_190), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_243), .Y(n_262) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_218), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_249), .B(n_190), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_208), .A2(n_190), .B1(n_200), .B2(n_195), .Y(n_265) );
NOR2xp33_ASAP7_75t_R g266 ( .A(n_227), .B(n_190), .Y(n_266) );
BUFx12f_ASAP7_75t_L g267 ( .A(n_227), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_258), .Y(n_268) );
OAI22xp5_ASAP7_75t_SL g269 ( .A1(n_257), .A2(n_87), .B1(n_88), .B2(n_89), .Y(n_269) );
AO21x1_ASAP7_75t_L g270 ( .A1(n_244), .A2(n_168), .B(n_161), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_258), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_208), .A2(n_200), .B1(n_191), .B2(n_195), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_257), .B(n_191), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_258), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_249), .B(n_204), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_218), .Y(n_276) );
AOI22xp33_ASAP7_75t_SL g277 ( .A1(n_210), .A2(n_204), .B1(n_198), .B2(n_192), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_218), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_214), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_205), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_248), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_205), .B(n_204), .Y(n_282) );
NAND2xp33_ASAP7_75t_L g283 ( .A(n_252), .B(n_197), .Y(n_283) );
INVxp67_ASAP7_75t_L g284 ( .A(n_207), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_SL g285 ( .A1(n_235), .A2(n_154), .B(n_153), .C(n_158), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_214), .Y(n_286) );
INVx2_ASAP7_75t_SL g287 ( .A(n_235), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_220), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_237), .A2(n_159), .B(n_158), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_205), .B(n_198), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_249), .B(n_198), .Y(n_291) );
AO22x1_ASAP7_75t_L g292 ( .A1(n_210), .A2(n_88), .B1(n_95), .B2(n_102), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_213), .B(n_196), .Y(n_293) );
NOR2x1_ASAP7_75t_L g294 ( .A(n_233), .B(n_196), .Y(n_294) );
NAND2x2_ASAP7_75t_L g295 ( .A(n_212), .B(n_4), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_209), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_213), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_222), .A2(n_192), .B(n_196), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_213), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_249), .B(n_192), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_243), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_211), .B(n_217), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_233), .A2(n_197), .B1(n_120), .B2(n_95), .Y(n_303) );
INVx3_ASAP7_75t_SL g304 ( .A(n_248), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_243), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_234), .A2(n_197), .B1(n_90), .B2(n_153), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_234), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
AOI222xp33_ASAP7_75t_L g309 ( .A1(n_284), .A2(n_239), .B1(n_221), .B2(n_206), .C1(n_229), .C2(n_223), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_267), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_267), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_296), .B(n_244), .Y(n_312) );
BUFx4f_ASAP7_75t_SL g313 ( .A(n_304), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_298), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_273), .B(n_219), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_269), .A2(n_229), .B1(n_238), .B2(n_250), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
INVx6_ASAP7_75t_L g319 ( .A(n_280), .Y(n_319) );
BUFx10_ASAP7_75t_L g320 ( .A(n_268), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_264), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g322 ( .A1(n_272), .A2(n_256), .B(n_241), .C(n_238), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_288), .B(n_216), .Y(n_323) );
NOR2xp67_ASAP7_75t_SL g324 ( .A(n_280), .B(n_251), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_280), .Y(n_325) );
NOR2xp33_ASAP7_75t_R g326 ( .A(n_279), .B(n_251), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_298), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_280), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_282), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_280), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_264), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_272), .A2(n_241), .B(n_230), .C(n_260), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_275), .B(n_229), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_269), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_307), .A2(n_229), .B1(n_242), .B2(n_254), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_275), .B(n_209), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_302), .A2(n_236), .B1(n_231), .B2(n_224), .C(n_226), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_315), .B(n_291), .Y(n_338) );
NAND2x1p5_ASAP7_75t_L g339 ( .A(n_324), .B(n_280), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_332), .A2(n_215), .B(n_225), .C(n_228), .Y(n_340) );
OAI21x1_ASAP7_75t_SL g341 ( .A1(n_312), .A2(n_270), .B(n_299), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_318), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_329), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_318), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_336), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_315), .B(n_291), .Y(n_346) );
INVx4_ASAP7_75t_SL g347 ( .A(n_319), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_334), .B(n_300), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_323), .A2(n_295), .B1(n_270), .B2(n_266), .Y(n_349) );
OAI21x1_ASAP7_75t_L g350 ( .A1(n_314), .A2(n_294), .B(n_289), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_322), .A2(n_317), .B1(n_312), .B2(n_277), .Y(n_351) );
INVx4_ASAP7_75t_SL g352 ( .A(n_319), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_336), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_329), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_314), .A2(n_294), .B(n_306), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_333), .B(n_300), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_337), .A2(n_279), .B1(n_286), .B2(n_292), .C(n_255), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
O2A1O1Ixp33_ASAP7_75t_L g359 ( .A1(n_337), .A2(n_263), .B(n_278), .C(n_276), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_314), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_321), .B(n_292), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_327), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_335), .A2(n_295), .B1(n_265), .B2(n_268), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_351), .A2(n_338), .B1(n_353), .B2(n_345), .C(n_331), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_357), .A2(n_331), .B1(n_321), .B2(n_333), .C(n_335), .Y(n_365) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_349), .B(n_309), .C(n_306), .D(n_259), .Y(n_366) );
OAI33xp33_ASAP7_75t_L g367 ( .A1(n_363), .A2(n_259), .A3(n_286), .B1(n_159), .B2(n_154), .B3(n_155), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_346), .Y(n_368) );
AO21x2_ASAP7_75t_L g369 ( .A1(n_341), .A2(n_327), .B(n_285), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_342), .B(n_325), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_360), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_339), .Y(n_372) );
OAI321xp33_ASAP7_75t_L g373 ( .A1(n_361), .A2(n_316), .A3(n_308), .B1(n_303), .B2(n_327), .C(n_225), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_344), .B(n_325), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_360), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_354), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_362), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_355), .A2(n_330), .B(n_328), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_362), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_346), .B(n_308), .Y(n_380) );
AOI33xp33_ASAP7_75t_L g381 ( .A1(n_359), .A2(n_155), .A3(n_177), .B1(n_179), .B2(n_161), .B3(n_162), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_348), .A2(n_309), .B1(n_316), .B2(n_276), .C(n_330), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_326), .B(n_328), .C(n_330), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_340), .A2(n_330), .B1(n_328), .B2(n_325), .C(n_274), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_343), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_358), .B(n_325), .Y(n_386) );
OAI31xp33_ASAP7_75t_SL g387 ( .A1(n_355), .A2(n_282), .A3(n_290), .B(n_293), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_356), .B(n_311), .Y(n_388) );
OAI22xp33_ASAP7_75t_L g389 ( .A1(n_361), .A2(n_313), .B1(n_304), .B2(n_328), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_343), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_356), .A2(n_319), .B1(n_299), .B2(n_324), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_350), .Y(n_392) );
NAND3xp33_ASAP7_75t_L g393 ( .A(n_340), .B(n_169), .C(n_163), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_347), .B(n_215), .Y(n_395) );
NAND3xp33_ASAP7_75t_L g396 ( .A(n_387), .B(n_197), .C(n_169), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_385), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_379), .B(n_347), .Y(n_398) );
AOI211x1_ASAP7_75t_L g399 ( .A1(n_382), .A2(n_5), .B(n_6), .C(n_7), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_379), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_365), .A2(n_339), .B1(n_304), .B2(n_319), .C(n_287), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_372), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_364), .A2(n_310), .B1(n_197), .B2(n_245), .C(n_228), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_378), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_371), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_378), .B(n_352), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_375), .B(n_347), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_375), .B(n_352), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_385), .B(n_350), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_377), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_372), .Y(n_413) );
INVx4_ASAP7_75t_L g414 ( .A(n_372), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_377), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_380), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_368), .B(n_352), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_377), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_368), .B(n_352), .Y(n_419) );
BUFx2_ASAP7_75t_L g420 ( .A(n_378), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_390), .B(n_197), .Y(n_421) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_387), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_376), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_390), .B(n_245), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_392), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_364), .B(n_163), .C(n_169), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_380), .B(n_7), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_376), .B(n_365), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_382), .A2(n_319), .B1(n_287), .B2(n_299), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_370), .B(n_374), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_386), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_370), .B(n_8), .Y(n_432) );
OAI31xp33_ASAP7_75t_L g433 ( .A1(n_383), .A2(n_290), .A3(n_282), .B(n_293), .Y(n_433) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_381), .B(n_163), .C(n_169), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_386), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_374), .B(n_9), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_392), .B(n_395), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_366), .B(n_163), .C(n_169), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_394), .B(n_9), .Y(n_439) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_388), .A2(n_283), .B1(n_282), .B2(n_290), .C1(n_293), .C2(n_262), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_369), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_437), .B(n_369), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_405), .B(n_383), .C(n_366), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_437), .B(n_369), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_423), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_423), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_416), .B(n_389), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_430), .B(n_369), .Y(n_448) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_414), .B(n_395), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_430), .B(n_391), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_397), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_402), .B(n_393), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_402), .B(n_393), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_402), .B(n_11), .Y(n_454) );
NAND2xp33_ASAP7_75t_R g455 ( .A(n_408), .B(n_11), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_403), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_403), .B(n_13), .Y(n_457) );
AOI21xp33_ASAP7_75t_SL g458 ( .A1(n_396), .A2(n_13), .B(n_14), .Y(n_458) );
NOR2xp67_ASAP7_75t_SL g459 ( .A(n_396), .B(n_373), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_403), .B(n_14), .Y(n_460) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_414), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_415), .B(n_15), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_415), .B(n_15), .Y(n_463) );
NAND4xp25_ASAP7_75t_SL g464 ( .A(n_440), .B(n_384), .C(n_367), .D(n_19), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_400), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_415), .B(n_17), .Y(n_466) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_422), .A2(n_384), .B1(n_274), .B2(n_168), .C(n_177), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_431), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_439), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_428), .B(n_18), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_414), .Y(n_471) );
NOR2xp33_ASAP7_75t_R g472 ( .A(n_413), .B(n_18), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_411), .B(n_20), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_407), .B(n_21), .Y(n_474) );
INVxp33_ASAP7_75t_L g475 ( .A(n_398), .Y(n_475) );
AOI32xp33_ASAP7_75t_L g476 ( .A1(n_436), .A2(n_373), .A3(n_21), .B1(n_290), .B2(n_293), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_435), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_426), .A2(n_367), .B(n_297), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_411), .B(n_166), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_412), .B(n_418), .Y(n_480) );
NOR2xp67_ASAP7_75t_SL g481 ( .A(n_426), .B(n_438), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_433), .A2(n_297), .B(n_281), .C(n_301), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_412), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_429), .A2(n_166), .B1(n_183), .B2(n_180), .C(n_179), .Y(n_484) );
NAND2xp33_ASAP7_75t_L g485 ( .A(n_413), .B(n_297), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_418), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_427), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_414), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_425), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_427), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_432), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_398), .Y(n_493) );
AOI21xp33_ASAP7_75t_L g494 ( .A1(n_455), .A2(n_432), .B(n_404), .Y(n_494) );
OAI32xp33_ASAP7_75t_L g495 ( .A1(n_461), .A2(n_438), .A3(n_419), .B1(n_417), .B2(n_410), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_443), .A2(n_436), .B1(n_409), .B2(n_410), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_488), .B(n_399), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_451), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_481), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_491), .B(n_399), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_449), .A2(n_408), .B(n_409), .C(n_434), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_464), .A2(n_401), .B1(n_434), .B2(n_408), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_449), .A2(n_408), .B(n_420), .C(n_406), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_492), .A2(n_425), .B1(n_424), .B2(n_420), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_468), .B(n_424), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_465), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_471), .A2(n_421), .B1(n_406), .B2(n_441), .Y(n_507) );
OAI32xp33_ASAP7_75t_L g508 ( .A1(n_475), .A2(n_406), .A3(n_441), .B1(n_421), .B2(n_168), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_471), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_445), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_459), .B(n_406), .C(n_441), .Y(n_511) );
OAI32xp33_ASAP7_75t_L g512 ( .A1(n_475), .A2(n_183), .A3(n_180), .B1(n_179), .B2(n_177), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_477), .B(n_162), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_489), .A2(n_320), .B1(n_305), .B2(n_301), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_490), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_446), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_493), .B(n_23), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_469), .B(n_162), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_483), .Y(n_519) );
AOI32xp33_ASAP7_75t_L g520 ( .A1(n_489), .A2(n_281), .A3(n_166), .B1(n_161), .B2(n_183), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_486), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_473), .B(n_180), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_487), .A2(n_163), .B1(n_169), .B2(n_174), .C(n_188), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_472), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_458), .A2(n_305), .B(n_262), .C(n_320), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_473), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_480), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_481), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_470), .A2(n_163), .B1(n_174), .B2(n_188), .C(n_156), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_476), .A2(n_174), .B1(n_188), .B2(n_156), .C(n_250), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g531 ( .A(n_459), .B(n_174), .C(n_188), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_485), .A2(n_246), .B(n_232), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_448), .B(n_24), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_450), .A2(n_174), .B1(n_188), .B2(n_320), .Y(n_534) );
NOR2x1_ASAP7_75t_L g535 ( .A(n_485), .B(n_188), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_474), .B(n_174), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_467), .A2(n_320), .B1(n_156), .B2(n_253), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_527), .B(n_448), .Y(n_538) );
AND3x2_ASAP7_75t_L g539 ( .A(n_499), .B(n_457), .C(n_454), .Y(n_539) );
AOI222xp33_ASAP7_75t_L g540 ( .A1(n_524), .A2(n_442), .B1(n_444), .B2(n_447), .C1(n_457), .C2(n_460), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g541 ( .A1(n_526), .A2(n_442), .B1(n_444), .B2(n_460), .C1(n_462), .C2(n_463), .Y(n_541) );
AOI211xp5_ASAP7_75t_L g542 ( .A1(n_494), .A2(n_462), .B(n_466), .C(n_478), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_506), .Y(n_543) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_509), .B(n_466), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_498), .B(n_490), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_515), .B(n_453), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_510), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_497), .B(n_479), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_496), .A2(n_502), .B1(n_500), .B2(n_528), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_516), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_505), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_504), .B(n_453), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_515), .B(n_452), .Y(n_553) );
CKINVDCx16_ASAP7_75t_R g554 ( .A(n_533), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_499), .A2(n_452), .B1(n_456), .B2(n_482), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_507), .B(n_456), .Y(n_556) );
OA22x2_ASAP7_75t_L g557 ( .A1(n_528), .A2(n_25), .B1(n_26), .B2(n_36), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_503), .B(n_38), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_519), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_517), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_535), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_511), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_530), .A2(n_484), .B1(n_156), .B2(n_250), .Y(n_563) );
NAND3xp33_ASAP7_75t_SL g564 ( .A(n_525), .B(n_39), .C(n_40), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_504), .B(n_46), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_521), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_501), .B(n_156), .Y(n_567) );
NAND3xp33_ASAP7_75t_SL g568 ( .A(n_542), .B(n_537), .C(n_520), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_564), .A2(n_495), .B(n_508), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_562), .A2(n_518), .B(n_513), .C(n_522), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_544), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_540), .B(n_536), .Y(n_572) );
XNOR2xp5_ASAP7_75t_L g573 ( .A(n_560), .B(n_551), .Y(n_573) );
NAND2xp33_ASAP7_75t_SL g574 ( .A(n_554), .B(n_537), .Y(n_574) );
OAI211xp5_ASAP7_75t_L g575 ( .A1(n_549), .A2(n_514), .B(n_534), .C(n_531), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_545), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_548), .A2(n_529), .B1(n_523), .B2(n_532), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_557), .A2(n_512), .B(n_246), .Y(n_578) );
OAI221xp5_ASAP7_75t_L g579 ( .A1(n_562), .A2(n_261), .B1(n_247), .B2(n_240), .C(n_232), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_548), .A2(n_541), .B1(n_552), .B2(n_555), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_546), .B(n_47), .Y(n_581) );
BUFx3_ASAP7_75t_L g582 ( .A(n_561), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_543), .Y(n_583) );
AOI322xp5_ASAP7_75t_L g584 ( .A1(n_574), .A2(n_538), .A3(n_553), .B1(n_545), .B2(n_547), .C1(n_559), .C2(n_550), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_582), .B(n_556), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_571), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_580), .B(n_566), .Y(n_587) );
AOI21xp33_ASAP7_75t_SL g588 ( .A1(n_573), .A2(n_557), .B(n_558), .Y(n_588) );
NAND2xp33_ASAP7_75t_R g589 ( .A(n_569), .B(n_539), .Y(n_589) );
XNOR2xp5_ASAP7_75t_L g590 ( .A(n_572), .B(n_539), .Y(n_590) );
OA22x2_ASAP7_75t_L g591 ( .A1(n_576), .A2(n_565), .B1(n_563), .B2(n_567), .Y(n_591) );
AOI211xp5_ASAP7_75t_L g592 ( .A1(n_568), .A2(n_253), .B(n_247), .C(n_240), .Y(n_592) );
AOI21xp33_ASAP7_75t_L g593 ( .A1(n_570), .A2(n_50), .B(n_59), .Y(n_593) );
NAND5xp2_ASAP7_75t_L g594 ( .A(n_569), .B(n_575), .C(n_577), .D(n_578), .E(n_581), .Y(n_594) );
NAND3xp33_ASAP7_75t_SL g595 ( .A(n_575), .B(n_253), .C(n_579), .Y(n_595) );
AOI211xp5_ASAP7_75t_SL g596 ( .A1(n_583), .A2(n_494), .B(n_568), .C(n_575), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g597 ( .A1(n_574), .A2(n_582), .B(n_571), .C(n_569), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_590), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_586), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_589), .Y(n_600) );
OR3x2_ASAP7_75t_L g601 ( .A(n_594), .B(n_596), .C(n_588), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_600), .A2(n_597), .B1(n_595), .B2(n_591), .C(n_584), .Y(n_602) );
NOR3xp33_ASAP7_75t_L g603 ( .A(n_598), .B(n_592), .C(n_593), .Y(n_603) );
INVx3_ASAP7_75t_L g604 ( .A(n_602), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_603), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_605), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_606), .A2(n_604), .B1(n_601), .B2(n_599), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_607), .A2(n_604), .B1(n_601), .B2(n_587), .C(n_585), .Y(n_608) );
endmodule