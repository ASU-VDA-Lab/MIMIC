module fake_jpeg_19106_n_236 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_28),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_52),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_59),
.Y(n_78)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_44),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_17),
.B1(n_27),
.B2(n_16),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_33),
.B1(n_19),
.B2(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_31),
.Y(n_64)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_45),
.B1(n_41),
.B2(n_42),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_36),
.A2(n_31),
.B1(n_26),
.B2(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_71),
.B1(n_25),
.B2(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_42),
.B1(n_41),
.B2(n_26),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_30),
.CON(n_72),
.SN(n_72)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_30),
.B(n_23),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_38),
.A2(n_33),
.B1(n_19),
.B2(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_47),
.Y(n_81)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_99),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_89),
.B(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_92),
.B(n_95),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_44),
.B(n_38),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_46),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_44),
.B(n_21),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_44),
.B(n_21),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_10),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_10),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_101),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_11),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_105),
.B(n_1),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_107),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_108),
.B(n_110),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_75),
.B(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_15),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_11),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_23),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_91),
.B1(n_68),
.B2(n_58),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_77),
.B1(n_54),
.B2(n_69),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_124),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_21),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_83),
.C(n_88),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_22),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_46),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_22),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_102),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_151),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_88),
.B1(n_105),
.B2(n_79),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_154),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_103),
.B1(n_79),
.B2(n_77),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_117),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_102),
.B1(n_54),
.B2(n_56),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_155),
.B1(n_125),
.B2(n_117),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_146),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_86),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_86),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_150),
.B(n_152),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_94),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_12),
.C(n_14),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_87),
.B1(n_76),
.B2(n_84),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_84),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_156),
.B(n_132),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_145),
.B1(n_142),
.B2(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_121),
.C(n_131),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_133),
.C(n_134),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_110),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_171),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_169),
.B1(n_149),
.B2(n_145),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_114),
.B(n_122),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_115),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_114),
.B(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_109),
.B1(n_127),
.B2(n_126),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_143),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_181),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_158),
.B1(n_170),
.B2(n_166),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_2),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_189),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_109),
.C(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_169),
.A2(n_153),
.B1(n_135),
.B2(n_132),
.C(n_22),
.Y(n_190)
);

OA21x2_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_174),
.B(n_158),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_167),
.C(n_171),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_157),
.C(n_172),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_196),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_198),
.C(n_184),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_183),
.B(n_153),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_173),
.C(n_154),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_188),
.A2(n_160),
.B1(n_126),
.B2(n_118),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_204),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_160),
.B(n_3),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_2),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_192),
.C(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_212),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_197),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_211),
.B(n_213),
.Y(n_217)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_186),
.C(n_180),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_214),
.B(n_3),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_216),
.C(n_221),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_200),
.B(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_218),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_207),
.B(n_203),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_201),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_177),
.B(n_185),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_205),
.B(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_208),
.C(n_180),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_220),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_226),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_224),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_14),
.B(n_5),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_230),
.A2(n_6),
.B(n_7),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_231),
.B(n_232),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_4),
.C(n_5),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_233),
.A2(n_227),
.B(n_7),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_234),
.Y(n_236)
);


endmodule