module fake_jpeg_1281_n_443 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_443);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_443;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_11),
.B(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_47),
.Y(n_133)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_48),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_8),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_63),
.Y(n_104)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_57),
.Y(n_117)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_8),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_73),
.Y(n_89)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_81),
.Y(n_92)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_84),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_18),
.B(n_8),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_87),
.B(n_20),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_57),
.B1(n_73),
.B2(n_51),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_88),
.A2(n_108),
.B1(n_125),
.B2(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_90),
.B(n_111),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_17),
.B1(n_39),
.B2(n_37),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_91),
.A2(n_29),
.B1(n_43),
.B2(n_40),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_45),
.A2(n_20),
.B1(n_16),
.B2(n_39),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_95),
.A2(n_123),
.B1(n_43),
.B2(n_32),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_44),
.A2(n_20),
.B1(n_27),
.B2(n_39),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_33),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_50),
.A2(n_16),
.B1(n_27),
.B2(n_21),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_17),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_136),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_46),
.A2(n_33),
.B1(n_29),
.B2(n_37),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_49),
.A2(n_17),
.B1(n_21),
.B2(n_37),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_77),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_33),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_140),
.B(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_78),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_141),
.B(n_170),
.Y(n_195)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_134),
.Y(n_144)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_144),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_145),
.A2(n_174),
.B1(n_156),
.B2(n_148),
.Y(n_192)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_65),
.B1(n_54),
.B2(n_71),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_155),
.B1(n_166),
.B2(n_175),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_43),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_100),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_89),
.A2(n_36),
.B(n_35),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_157),
.B(n_140),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_21),
.B1(n_27),
.B2(n_29),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_173),
.B1(n_32),
.B2(n_34),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_69),
.B1(n_55),
.B2(n_74),
.Y(n_155)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_103),
.A2(n_35),
.B1(n_30),
.B2(n_32),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_158),
.Y(n_216)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_164),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_119),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_167),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_172),
.Y(n_203)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_180),
.C(n_98),
.Y(n_202)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_113),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_0),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_97),
.C(n_98),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_115),
.A2(n_35),
.B1(n_30),
.B2(n_40),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_118),
.A2(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_84),
.B1(n_82),
.B2(n_36),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_177),
.Y(n_207)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_101),
.Y(n_206)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_144),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_129),
.B(n_34),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_139),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_183),
.B(n_208),
.C(n_210),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_135),
.B(n_126),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_148),
.B(n_175),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_192),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_145),
.C(n_179),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_159),
.A2(n_133),
.B1(n_132),
.B2(n_116),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_201),
.B1(n_178),
.B2(n_152),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_200),
.B(n_3),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_132),
.B1(n_121),
.B2(n_130),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_144),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_109),
.B(n_114),
.C(n_121),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_157),
.Y(n_224)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_105),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_143),
.B(n_105),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_101),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_130),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_220),
.A2(n_234),
.B(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_149),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_224),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_210),
.C(n_193),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_184),
.A2(n_190),
.B1(n_191),
.B2(n_188),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_226),
.A2(n_230),
.B1(n_241),
.B2(n_247),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_145),
.B1(n_146),
.B2(n_165),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_228),
.A2(n_239),
.B1(n_240),
.B2(n_251),
.Y(n_280)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_184),
.A2(n_145),
.B1(n_106),
.B2(n_142),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_232),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_190),
.A2(n_158),
.B1(n_160),
.B2(n_162),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_196),
.A2(n_170),
.B1(n_172),
.B2(n_168),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_188),
.B(n_163),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_242),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_138),
.B1(n_176),
.B2(n_161),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_106),
.B1(n_177),
.B2(n_169),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_196),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_217),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_206),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_243),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_8),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_244),
.B(n_245),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_195),
.B(n_191),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_189),
.A2(n_0),
.B(n_1),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_246),
.A2(n_220),
.B(n_224),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_211),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_249),
.A2(n_250),
.B1(n_214),
.B2(n_194),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_204),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_254),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_231),
.A2(n_232),
.B1(n_218),
.B2(n_243),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_256),
.A2(n_257),
.B1(n_262),
.B2(n_267),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_181),
.B1(n_186),
.B2(n_183),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_236),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_260),
.A2(n_261),
.B(n_270),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_181),
.B(n_199),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_228),
.A2(n_215),
.B1(n_205),
.B2(n_200),
.Y(n_262)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_230),
.A2(n_199),
.B(n_209),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_223),
.B(n_205),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_266),
.B(n_273),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_237),
.A2(n_207),
.B1(n_209),
.B2(n_182),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_214),
.B(n_187),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_234),
.B1(n_235),
.B2(n_239),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_223),
.A2(n_182),
.B1(n_194),
.B2(n_185),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_272),
.A2(n_229),
.B1(n_247),
.B2(n_241),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_236),
.B(n_185),
.CI(n_216),
.CON(n_273),
.SN(n_273)
);

NAND4xp25_ASAP7_75t_SL g276 ( 
.A(n_251),
.B(n_216),
.C(n_5),
.D(n_6),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_281),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_4),
.C(n_7),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_246),
.C(n_238),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_222),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_227),
.B(n_4),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_283),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_293),
.C(n_295),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_285),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_298),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_255),
.B1(n_261),
.B2(n_263),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_225),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_264),
.B1(n_265),
.B2(n_275),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_294),
.A2(n_253),
.B1(n_268),
.B2(n_254),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_225),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_260),
.A2(n_219),
.B(n_246),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_296),
.A2(n_255),
.B(n_275),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_256),
.B(n_238),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_299),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_264),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_238),
.C(n_252),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_301),
.C(n_281),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_252),
.B(n_226),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_259),
.A2(n_242),
.B1(n_250),
.B2(n_244),
.Y(n_302)
);

OAI22x1_ASAP7_75t_SL g329 ( 
.A1(n_302),
.A2(n_306),
.B1(n_234),
.B2(n_273),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_278),
.A2(n_250),
.B1(n_221),
.B2(n_240),
.Y(n_303)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_304),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_267),
.A2(n_250),
.B1(n_248),
.B2(n_227),
.Y(n_306)
);

NOR2x1_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_235),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_310),
.Y(n_335)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_254),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_301),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_320),
.B1(n_329),
.B2(n_334),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_287),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_315),
.B(n_318),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_287),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_319),
.A2(n_306),
.B(n_307),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_280),
.B1(n_263),
.B2(n_265),
.Y(n_320)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_302),
.Y(n_358)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_328),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_284),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_336),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_269),
.C(n_279),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_296),
.C(n_299),
.Y(n_354)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_288),
.A2(n_280),
.B1(n_263),
.B2(n_262),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_300),
.B(n_253),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_338),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_291),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_340),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_312),
.B(n_289),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_343),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_337),
.Y(n_344)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_319),
.A2(n_308),
.B(n_292),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_347),
.A2(n_353),
.B1(n_356),
.B2(n_328),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_335),
.A2(n_288),
.B(n_292),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_291),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_352),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_297),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_312),
.B(n_282),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_358),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_316),
.B(n_286),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_355),
.A2(n_324),
.B1(n_316),
.B2(n_335),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_317),
.A2(n_310),
.B1(n_286),
.B2(n_309),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_359),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_274),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_360),
.B(n_326),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_368),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_365),
.A2(n_357),
.B1(n_339),
.B2(n_356),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_360),
.B(n_326),
.C(n_327),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_370),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_361),
.A2(n_317),
.B1(n_322),
.B2(n_323),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_367),
.B(n_369),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_351),
.B(n_336),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_361),
.A2(n_322),
.B1(n_323),
.B2(n_330),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_332),
.C(n_329),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_338),
.C(n_314),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_374),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_348),
.A2(n_343),
.B1(n_320),
.B2(n_350),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_321),
.C(n_334),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_355),
.C(n_357),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_358),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_385),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_378),
.A2(n_341),
.B(n_359),
.Y(n_382)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_378),
.A2(n_346),
.B(n_348),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_384),
.A2(n_396),
.B(n_362),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_352),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_353),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_387),
.B(n_391),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_347),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_393),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_390),
.A2(n_333),
.B1(n_377),
.B2(n_274),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_345),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_339),
.C(n_321),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_229),
.C(n_276),
.Y(n_404)
);

AOI21x1_ASAP7_75t_L g396 ( 
.A1(n_371),
.A2(n_345),
.B(n_349),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_397),
.A2(n_399),
.B(n_402),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_390),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_404),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_386),
.A2(n_364),
.B(n_365),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_392),
.A2(n_373),
.B1(n_349),
.B2(n_370),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_400),
.A2(n_405),
.B1(n_383),
.B2(n_12),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_401),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_384),
.A2(n_368),
.B(n_277),
.Y(n_402)
);

INVx11_ASAP7_75t_L g405 ( 
.A(n_395),
.Y(n_405)
);

XOR2x2_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_229),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_383),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_392),
.A2(n_9),
.B(n_10),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_408),
.A2(n_11),
.B(n_12),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_407),
.B(n_394),
.C(n_389),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_413),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_381),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_388),
.C(n_385),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_415),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_402),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_397),
.C(n_399),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_418),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_11),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_420),
.B(n_421),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_12),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_403),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_416),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_401),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_427),
.A2(n_413),
.B(n_411),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_430),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_419),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_433),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_423),
.B(n_422),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_434),
.A2(n_405),
.B(n_408),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_422),
.Y(n_435)
);

AO21x2_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_424),
.B(n_425),
.Y(n_436)
);

NAND4xp25_ASAP7_75t_SL g439 ( 
.A(n_436),
.B(n_438),
.C(n_432),
.D(n_429),
.Y(n_439)
);

OAI321xp33_ASAP7_75t_L g440 ( 
.A1(n_439),
.A2(n_437),
.A3(n_404),
.B1(n_15),
.B2(n_14),
.C(n_13),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_440),
.A2(n_13),
.B(n_14),
.Y(n_441)
);

BUFx24_ASAP7_75t_SL g442 ( 
.A(n_441),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_442),
.A2(n_13),
.B(n_15),
.Y(n_443)
);


endmodule