module fake_jpeg_1980_n_474 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_474);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_474;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_73),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_55),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_60),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_16),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_61),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_14),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_79),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_63),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_68),
.Y(n_135)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_18),
.B(n_14),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_31),
.B(n_0),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

HAxp5_ASAP7_75t_SL g81 ( 
.A(n_25),
.B(n_13),
.CON(n_81),
.SN(n_81)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_85),
.Y(n_109)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_34),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_91),
.B(n_107),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_47),
.A2(n_64),
.B1(n_63),
.B2(n_83),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_93),
.A2(n_137),
.B1(n_21),
.B2(n_25),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_49),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_54),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_110),
.B(n_115),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_50),
.B(n_65),
.C(n_59),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_114),
.B(n_13),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_34),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_20),
.B1(n_44),
.B2(n_40),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_117),
.A2(n_128),
.B1(n_147),
.B2(n_4),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_58),
.B(n_41),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_119),
.B(n_123),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_45),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_122),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_45),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_66),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_41),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_124),
.B(n_125),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_67),
.B(n_19),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_44),
.B1(n_40),
.B2(n_33),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_78),
.B(n_19),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_130),
.B(n_132),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_35),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_74),
.A2(n_20),
.B1(n_40),
.B2(n_33),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_76),
.A2(n_22),
.B1(n_23),
.B2(n_35),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_144),
.A2(n_145),
.B1(n_8),
.B2(n_9),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_80),
.A2(n_22),
.B1(n_23),
.B2(n_33),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_88),
.A2(n_44),
.B1(n_20),
.B2(n_28),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_149),
.A2(n_156),
.B1(n_162),
.B2(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_150),
.Y(n_204)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_153),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_98),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_103),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_169),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_158),
.Y(n_234)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_159),
.B(n_163),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_27),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_176),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_167),
.A2(n_168),
.B1(n_190),
.B2(n_202),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_109),
.A2(n_25),
.B1(n_21),
.B2(n_38),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_136),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_170),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_109),
.A2(n_25),
.B(n_21),
.C(n_38),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_171),
.B(n_203),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_105),
.B(n_1),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_117),
.A2(n_1),
.B(n_2),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_177),
.B(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_95),
.B(n_3),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_180),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_179),
.A2(n_198),
.B1(n_13),
.B2(n_10),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_96),
.B(n_4),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_187),
.Y(n_237)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_108),
.Y(n_213)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_90),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_191),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_93),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_90),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_127),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_97),
.B(n_6),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_196),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_194),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_94),
.B(n_8),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_8),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_133),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_200),
.Y(n_220)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_135),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_205),
.B(n_233),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_213),
.B(n_199),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_99),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_223),
.B(n_231),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_164),
.A2(n_147),
.B1(n_129),
.B2(n_146),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_224),
.A2(n_185),
.B1(n_183),
.B2(n_201),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_167),
.A2(n_140),
.B1(n_141),
.B2(n_133),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_225),
.A2(n_235),
.B1(n_241),
.B2(n_153),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_226),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_152),
.B(n_101),
.C(n_143),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_251),
.C(n_166),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_143),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_152),
.B(n_134),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_190),
.A2(n_140),
.B1(n_141),
.B2(n_135),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_134),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_244),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_172),
.B(n_160),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_239),
.B(n_249),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_174),
.A2(n_202),
.B1(n_177),
.B2(n_180),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_247),
.B1(n_168),
.B2(n_188),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_171),
.A2(n_108),
.B1(n_131),
.B2(n_118),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_193),
.B(n_131),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_165),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_252),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_161),
.A2(n_128),
.B1(n_146),
.B2(n_129),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_176),
.B(n_9),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_150),
.B(n_10),
.C(n_11),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_158),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_255),
.Y(n_309)
);

BUFx12_ASAP7_75t_L g257 ( 
.A(n_252),
.Y(n_257)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_151),
.B(n_188),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_258),
.A2(n_251),
.B(n_216),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_259),
.A2(n_271),
.B(n_285),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_SL g260 ( 
.A1(n_238),
.A2(n_181),
.B(n_203),
.C(n_151),
.Y(n_260)
);

OA21x2_ASAP7_75t_L g301 ( 
.A1(n_260),
.A2(n_219),
.B(n_246),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g319 ( 
.A(n_261),
.B(n_258),
.C(n_264),
.Y(n_319)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_262),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_263),
.A2(n_270),
.B1(n_282),
.B2(n_294),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_264),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_206),
.A2(n_155),
.B1(n_170),
.B2(n_175),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_265),
.A2(n_273),
.B1(n_277),
.B2(n_287),
.Y(n_303)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_214),
.A2(n_200),
.B(n_186),
.Y(n_271)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_272),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_206),
.A2(n_198),
.B1(n_148),
.B2(n_154),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_214),
.A2(n_194),
.B1(n_173),
.B2(n_12),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_278),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_205),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_280),
.B(n_286),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_11),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_281),
.A2(n_291),
.B(n_284),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_212),
.A2(n_11),
.B1(n_12),
.B2(n_223),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_215),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_211),
.B(n_11),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_284),
.B(n_289),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_241),
.A2(n_12),
.B(n_233),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_210),
.B(n_229),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_212),
.A2(n_224),
.B1(n_228),
.B2(n_231),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_227),
.Y(n_288)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_239),
.B(n_250),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_243),
.A2(n_225),
.B1(n_237),
.B2(n_250),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_222),
.A2(n_208),
.B(n_213),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_237),
.A2(n_222),
.B1(n_232),
.B2(n_216),
.Y(n_292)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_208),
.B(n_211),
.C(n_249),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_295),
.C(n_254),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_235),
.A2(n_232),
.B1(n_246),
.B2(n_242),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_217),
.B(n_230),
.C(n_218),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_215),
.B(n_234),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_253),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_299),
.A2(n_301),
.B(n_308),
.Y(n_342)
);

CKINVDCx10_ASAP7_75t_R g302 ( 
.A(n_257),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_219),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_310),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_271),
.B(n_218),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g310 ( 
.A(n_259),
.B(n_230),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_285),
.A2(n_234),
.B(n_221),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_335),
.B(n_260),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_207),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_324),
.C(n_326),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_287),
.A2(n_207),
.B1(n_273),
.B2(n_270),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_317),
.A2(n_260),
.B1(n_257),
.B2(n_288),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_319),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_329),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_254),
.B(n_261),
.C(n_264),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_267),
.C(n_274),
.Y(n_326)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_268),
.C(n_256),
.Y(n_329)
);

NOR3xp33_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_260),
.C(n_269),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g332 ( 
.A(n_275),
.B(n_260),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_281),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_255),
.B(n_276),
.C(n_278),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_265),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_297),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_334),
.B(n_262),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_281),
.A2(n_269),
.B(n_277),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_283),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_348),
.C(n_352),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_302),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_345),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_315),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_346),
.A2(n_358),
.B1(n_363),
.B2(n_368),
.Y(n_380)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_322),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_347),
.B(n_357),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_282),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_300),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_351),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_298),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_272),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_353),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_301),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_342),
.Y(n_388)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_316),
.C(n_321),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_303),
.A2(n_294),
.B1(n_263),
.B2(n_272),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_309),
.Y(n_359)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_331),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_313),
.B(n_266),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_362),
.B(n_364),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_257),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_365),
.Y(n_389)
);

AO21x1_ASAP7_75t_L g366 ( 
.A1(n_306),
.A2(n_332),
.B(n_323),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_366),
.Y(n_379)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_303),
.A2(n_323),
.B1(n_317),
.B2(n_312),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_364),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_344),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_324),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_376),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_375),
.C(n_386),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_326),
.C(n_299),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_330),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_307),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_392),
.Y(n_408)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_381),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_361),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_388),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_331),
.C(n_306),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_308),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_328),
.Y(n_393)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_368),
.A2(n_312),
.B1(n_335),
.B2(n_311),
.Y(n_394)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_394),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_379),
.A2(n_308),
.B1(n_360),
.B2(n_354),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_396),
.A2(n_415),
.B1(n_388),
.B2(n_393),
.Y(n_428)
);

XNOR2x1_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_353),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_395),
.Y(n_424)
);

XOR2x1_ASAP7_75t_SL g399 ( 
.A(n_395),
.B(n_342),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_410),
.C(n_386),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_401),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_351),
.C(n_344),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_374),
.C(n_369),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_366),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_301),
.Y(n_435)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_387),
.Y(n_409)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_409),
.Y(n_422)
);

XOR2x2_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_346),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_340),
.Y(n_411)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_411),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_387),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_412),
.A2(n_414),
.B1(n_416),
.B2(n_382),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_367),
.Y(n_413)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_413),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_343),
.B1(n_308),
.B2(n_363),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_418),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_378),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_420),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_404),
.A2(n_379),
.B(n_384),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_423),
.A2(n_404),
.B(n_396),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_430),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_426),
.C(n_429),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_405),
.C(n_403),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_397),
.A2(n_377),
.B1(n_343),
.B2(n_369),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_427),
.A2(n_402),
.B1(n_414),
.B2(n_413),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_428),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_406),
.C(n_408),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_366),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_410),
.B(n_338),
.C(n_341),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_431),
.B(n_434),
.C(n_435),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_398),
.B(n_310),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_438),
.B(n_441),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_439),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_407),
.C(n_417),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_SL g443 ( 
.A1(n_424),
.A2(n_399),
.B(n_415),
.C(n_431),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_443),
.A2(n_435),
.B1(n_433),
.B2(n_430),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_417),
.C(n_345),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_445),
.B(n_446),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_422),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_432),
.A2(n_365),
.B(n_362),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_448),
.A2(n_371),
.B(n_372),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_437),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_450),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_429),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_421),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_452),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_455),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_325),
.Y(n_457)
);

AOI322xp5_ASAP7_75t_L g460 ( 
.A1(n_457),
.A2(n_318),
.A3(n_372),
.B1(n_371),
.B2(n_355),
.C1(n_359),
.C2(n_348),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_449),
.A2(n_443),
.B1(n_434),
.B2(n_420),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_452),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_460),
.A2(n_461),
.B(n_453),
.Y(n_464)
);

AOI322xp5_ASAP7_75t_L g461 ( 
.A1(n_456),
.A2(n_391),
.A3(n_389),
.B1(n_443),
.B2(n_442),
.C1(n_447),
.C2(n_318),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_466),
.C(n_467),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_463),
.A2(n_462),
.B(n_455),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_465),
.A2(n_458),
.B(n_443),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_450),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_468),
.B(n_447),
.Y(n_470)
);

NOR3xp33_ASAP7_75t_L g472 ( 
.A(n_470),
.B(n_471),
.C(n_442),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_469),
.B(n_389),
.Y(n_471)
);

O2A1O1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_472),
.A2(n_419),
.B(n_391),
.C(n_305),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_473),
.B(n_358),
.Y(n_474)
);


endmodule