module real_jpeg_30745_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_605;
wire n_216;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_0),
.Y(n_245)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_0),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_0),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_1),
.A2(n_337),
.B(n_340),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_1),
.B(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_1),
.Y(n_395)
);

OAI32xp33_ASAP7_75t_L g498 ( 
.A1(n_1),
.A2(n_148),
.A3(n_499),
.B1(n_503),
.B2(n_506),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_1),
.A2(n_395),
.B1(n_540),
.B2(n_541),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_1),
.B(n_120),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_1),
.A2(n_234),
.B1(n_614),
.B2(n_628),
.Y(n_627)
);

INVxp33_ASAP7_75t_L g663 ( 
.A(n_2),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_3),
.A2(n_54),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_3),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g277 ( 
.A1(n_3),
.A2(n_184),
.B1(n_278),
.B2(n_280),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_3),
.A2(n_184),
.B1(n_355),
.B2(n_358),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_3),
.A2(n_184),
.B1(n_377),
.B2(n_381),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_5),
.A2(n_54),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_5),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_5),
.A2(n_344),
.B1(n_367),
.B2(n_370),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_5),
.A2(n_344),
.B1(n_571),
.B2(n_573),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_5),
.A2(n_344),
.B1(n_615),
.B2(n_617),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_6),
.A2(n_57),
.B1(n_223),
.B2(n_226),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_6),
.A2(n_57),
.B1(n_215),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_6),
.A2(n_57),
.B1(n_239),
.B2(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_7),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_112),
.B1(n_132),
.B2(n_137),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_7),
.A2(n_112),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_8),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_8),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_8),
.A2(n_271),
.B1(n_350),
.B2(n_353),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_8),
.A2(n_271),
.B1(n_443),
.B2(n_444),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_8),
.A2(n_271),
.B1(n_515),
.B2(n_518),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_9),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_9),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_9),
.A2(n_263),
.B1(n_327),
.B2(n_331),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_9),
.A2(n_263),
.B1(n_353),
.B2(n_496),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_9),
.A2(n_238),
.B1(n_263),
.B2(n_583),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_10),
.A2(n_63),
.B1(n_67),
.B2(n_73),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_10),
.A2(n_73),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_10),
.A2(n_73),
.B1(n_253),
.B2(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_10),
.A2(n_73),
.B1(n_248),
.B2(n_419),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_11),
.A2(n_156),
.B1(n_160),
.B2(n_164),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_11),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_11),
.A2(n_164),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_11),
.A2(n_164),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_11),
.A2(n_164),
.B1(n_238),
.B2(n_243),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_13),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_13),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_14),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_14),
.Y(n_384)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_14),
.Y(n_587)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_21),
.B(n_662),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_16),
.B(n_663),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_17),
.A2(n_318),
.B1(n_322),
.B2(n_323),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_17),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_17),
.A2(n_54),
.B1(n_322),
.B2(n_435),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_17),
.A2(n_215),
.B1(n_322),
.B2(n_546),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g601 ( 
.A1(n_17),
.A2(n_322),
.B1(n_602),
.B2(n_605),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_18),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_18),
.Y(n_111)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_19),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_19),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_19),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_201),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_R g22 ( 
.A(n_23),
.B(n_199),
.Y(n_22)
);

NOR2x1_ASAP7_75t_R g23 ( 
.A(n_24),
.B(n_178),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_24),
.B(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_165),
.B2(n_166),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_74),
.C(n_117),
.Y(n_26)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_27),
.B(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_28),
.A2(n_61),
.B1(n_62),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_28),
.A2(n_61),
.B1(n_260),
.B2(n_267),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_28),
.A2(n_61),
.B1(n_336),
.B2(n_343),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_28),
.A2(n_61),
.B1(n_260),
.B2(n_434),
.Y(n_454)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_29),
.A2(n_52),
.B1(n_183),
.B2(n_188),
.Y(n_182)
);

AO22x1_ASAP7_75t_L g285 ( 
.A1(n_29),
.A2(n_183),
.B1(n_188),
.B2(n_268),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_29),
.A2(n_188),
.B1(n_433),
.B2(n_439),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_41),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_33),
.Y(n_262)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_33),
.Y(n_438)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_36),
.Y(n_402)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_37),
.Y(n_339)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_38),
.Y(n_342)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_40),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_41)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_42),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_43),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_43),
.Y(n_282)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_48),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_56),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_60),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_60),
.Y(n_266)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_61),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_61),
.B(n_395),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_65),
.Y(n_347)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_66),
.Y(n_406)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_71),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_72),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_74),
.A2(n_191),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_75),
.B(n_118),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_75),
.B(n_181),
.C(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_75),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_89),
.B(n_107),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_76),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_76),
.A2(n_218),
.B1(n_252),
.B2(n_254),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_76),
.A2(n_211),
.B1(n_218),
.B2(n_254),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_76),
.A2(n_218),
.B1(n_349),
.B2(n_354),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_76),
.A2(n_218),
.B1(n_252),
.B2(n_354),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_76),
.A2(n_218),
.B1(n_545),
.B2(n_569),
.Y(n_594)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp33_ASAP7_75t_SL g106 ( 
.A(n_78),
.Y(n_106)
);

AO21x2_ASAP7_75t_L g218 ( 
.A1(n_78),
.A2(n_91),
.B(n_100),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_78)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_79),
.Y(n_236)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_81),
.Y(n_380)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_81),
.Y(n_393)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_83),
.Y(n_562)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_86),
.Y(n_243)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_106),
.Y(n_89)
);

AO21x1_ASAP7_75t_L g554 ( 
.A1(n_90),
.A2(n_555),
.B(n_557),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_94),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_95),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_95),
.Y(n_352)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp67_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_105),
.Y(n_511)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_110),
.Y(n_360)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_110),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_111),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_111),
.Y(n_357)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx4f_ASAP7_75t_L g572 ( 
.A(n_114),
.Y(n_572)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_116),
.Y(n_579)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_131),
.B1(n_141),
.B2(n_155),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_119),
.A2(n_141),
.B1(n_155),
.B2(n_192),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_119),
.A2(n_141),
.B1(n_317),
.B2(n_366),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_119),
.A2(n_141),
.B1(n_326),
.B2(n_442),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_119),
.A2(n_141),
.B1(n_366),
.B2(n_539),
.Y(n_538)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

AOI22x1_ASAP7_75t_L g221 ( 
.A1(n_120),
.A2(n_168),
.B1(n_193),
.B2(n_222),
.Y(n_221)
);

AOI22x1_ASAP7_75t_L g276 ( 
.A1(n_120),
.A2(n_168),
.B1(n_222),
.B2(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_120),
.A2(n_168),
.B1(n_316),
.B2(n_325),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_120),
.A2(n_168),
.B1(n_277),
.B2(n_456),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_120),
.A2(n_168),
.B1(n_277),
.B2(n_456),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_142),
.B(n_148),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.Y(n_121)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_127),
.Y(n_505)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_136),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_136),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_136),
.Y(n_373)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_149),
.Y(n_443)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_150),
.Y(n_399)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_151),
.Y(n_369)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_151),
.Y(n_412)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_160),
.Y(n_540)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_189),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_179),
.B(n_181),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_182),
.Y(n_300)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_189),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_191),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_198),
.Y(n_279)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_658),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_310),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_304),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_292),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_205),
.B(n_292),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_230),
.C(n_283),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_207),
.A2(n_208),
.B1(n_284),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_221),
.B(n_229),
.Y(n_208)
);

NAND2x1p5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_221),
.Y(n_229)
);

AOI22x1_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_212),
.Y(n_353)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

BUFx6f_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_217),
.A2(n_220),
.B1(n_495),
.B2(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_217),
.Y(n_574)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_218),
.A2(n_349),
.B1(n_493),
.B2(n_494),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_220),
.Y(n_493)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_225),
.Y(n_324)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_228),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_229),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_229),
.B(n_293),
.C(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_230),
.B(n_477),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_258),
.C(n_275),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_231),
.A2(n_232),
.B1(n_471),
.B2(n_473),
.Y(n_470)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_251),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_233),
.B(n_251),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_237),
.B1(n_244),
.B2(n_246),
.Y(n_233)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_234),
.A2(n_237),
.B1(n_418),
.B2(n_427),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_234),
.A2(n_582),
.B1(n_588),
.B2(n_591),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_234),
.A2(n_601),
.B1(n_614),
.B2(n_621),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_241),
.Y(n_616)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_242),
.Y(n_517)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_242),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_242),
.Y(n_604)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_245),
.Y(n_416)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_246),
.Y(n_290)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_259),
.A2(n_275),
.B1(n_276),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_259),
.Y(n_472)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_284),
.Y(n_478)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_285),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_286),
.A2(n_296),
.B(n_468),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.Y(n_286)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B(n_290),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_288),
.A2(n_376),
.B1(n_385),
.B2(n_389),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_288),
.A2(n_389),
.B1(n_415),
.B2(n_417),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_288),
.A2(n_376),
.B1(n_514),
.B2(n_522),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_288),
.A2(n_600),
.B1(n_606),
.B2(n_607),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_296),
.B(n_297),
.Y(n_293)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_295),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AOI21x1_ASAP7_75t_SL g659 ( 
.A1(n_305),
.A2(n_660),
.B(n_661),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_SL g661 ( 
.A(n_306),
.B(n_308),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_487),
.B(n_649),
.Y(n_310)
);

NAND4xp25_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_448),
.C(n_474),
.D(n_479),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_422),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_313),
.B(n_422),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_363),
.C(n_396),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_314),
.B(n_646),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_334),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_315),
.B(n_361),
.C(n_362),
.Y(n_428)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_330),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_330),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_348),
.B1(n_361),
.B2(n_362),
.Y(n_334)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_340),
.Y(n_413)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_343),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_357),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_364),
.B(n_396),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_374),
.C(n_394),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_365),
.B(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_373),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_374),
.A2(n_375),
.B1(n_394),
.B2(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_380),
.Y(n_556)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx2_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_384),
.Y(n_560)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_384),
.Y(n_620)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_387),
.Y(n_632)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_388),
.Y(n_624)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_394),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_395),
.B(n_507),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_395),
.B(n_564),
.Y(n_563)
);

OA21x2_ASAP7_75t_SL g575 ( 
.A1(n_395),
.A2(n_563),
.B(n_576),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_SL g625 ( 
.A(n_395),
.B(n_493),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_395),
.B(n_631),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_414),
.B1(n_420),
.B2(n_421),
.Y(n_396)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

OAI32xp33_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_400),
.A3(n_403),
.B1(n_407),
.B2(n_413),
.Y(n_397)
);

OAI32xp33_ASAP7_75t_L g447 ( 
.A1(n_398),
.A2(n_400),
.A3(n_403),
.B1(n_407),
.B2(n_413),
.Y(n_447)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_SL g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_414),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_415),
.Y(n_427)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_419),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_421),
.B(n_447),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_429),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_428),
.Y(n_423)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_424),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_426),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_428),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_429),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_446),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_432),
.B1(n_440),
.B2(n_441),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_432),
.Y(n_459)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_458),
.C(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_442),
.Y(n_456)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_462),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_449),
.A2(n_462),
.B1(n_480),
.B2(n_651),
.Y(n_652)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_449),
.Y(n_655)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_457),
.C(n_460),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_461),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_453),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_452),
.B(n_465),
.C(n_466),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_454),
.Y(n_465)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_457),
.Y(n_485)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_462),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_469),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_467),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_467),
.C(n_470),
.Y(n_475)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_471),
.Y(n_473)
);

A2O1A1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_474),
.A2(n_650),
.B(n_652),
.C(n_653),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_475),
.B(n_476),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_484),
.Y(n_479)
);

OAI21xp33_ASAP7_75t_L g650 ( 
.A1(n_480),
.A2(n_484),
.B(n_651),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.C(n_483),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

AOI21x1_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_644),
.B(n_648),
.Y(n_487)
);

OAI21x1_ASAP7_75t_SL g488 ( 
.A1(n_489),
.A2(n_550),
.B(n_643),
.Y(n_488)
);

AOI211xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_528),
.B(n_533),
.C(n_534),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_L g643 ( 
.A1(n_490),
.A2(n_528),
.B(n_533),
.C(n_534),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_530),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_497),
.B1(n_526),
.B2(n_527),
.Y(n_491)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_492),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_492),
.B(n_526),
.C(n_529),
.Y(n_647)
);

OAI22x1_ASAP7_75t_L g568 ( 
.A1(n_493),
.A2(n_569),
.B1(n_574),
.B2(n_575),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_497),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_512),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_498),
.A2(n_512),
.B1(n_513),
.B2(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_498),
.Y(n_536)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_510),
.Y(n_567)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_511),
.Y(n_549)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_514),
.Y(n_591)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_520),
.Y(n_633)
);

BUFx12f_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_525),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_525),
.Y(n_609)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_537),
.C(n_543),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_535),
.B(n_640),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_537),
.A2(n_538),
.B1(n_543),
.B2(n_641),
.Y(n_640)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_543),
.Y(n_641)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_549),
.Y(n_548)
);

AOI21x1_ASAP7_75t_L g550 ( 
.A1(n_551),
.A2(n_637),
.B(n_642),
.Y(n_550)
);

OAI21x1_ASAP7_75t_SL g551 ( 
.A1(n_552),
.A2(n_597),
.B(n_636),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_553),
.B(n_580),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_553),
.B(n_580),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_568),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_SL g610 ( 
.A(n_554),
.B(n_568),
.Y(n_610)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_558),
.A2(n_561),
.B(n_563),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_581),
.B(n_592),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_581),
.B(n_594),
.C(n_595),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_582),
.Y(n_606)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_593),
.A2(n_594),
.B1(n_595),
.B2(n_596),
.Y(n_592)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_593),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_594),
.Y(n_596)
);

AOI21x1_ASAP7_75t_L g597 ( 
.A1(n_598),
.A2(n_611),
.B(n_635),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_610),
.Y(n_598)
);

NOR2xp67_ASAP7_75t_L g635 ( 
.A(n_599),
.B(n_610),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

INVx3_ASAP7_75t_SL g607 ( 
.A(n_608),
.Y(n_607)
);

INVx8_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_612),
.A2(n_626),
.B(n_634),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_625),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_613),
.B(n_625),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_622),
.Y(n_628)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_624),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_627),
.B(n_629),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_630),
.B(n_633),
.Y(n_629)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_638),
.B(n_639),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_SL g642 ( 
.A(n_638),
.B(n_639),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_645),
.B(n_647),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_645),
.B(n_647),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_654),
.B(n_657),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_655),
.B(n_656),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);


endmodule