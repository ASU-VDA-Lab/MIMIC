module fake_jpeg_22953_n_220 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_0),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_53),
.B1(n_68),
.B2(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_55),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_22),
.B1(n_24),
.B2(n_20),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_26),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_56),
.B(n_62),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_25),
.Y(n_72)
);

BUFx12f_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_3),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_32),
.B1(n_21),
.B2(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_54),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_33),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_75),
.B(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_15),
.Y(n_76)
);

OR2x4_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_37),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_46),
.B(n_51),
.Y(n_119)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_25),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_1),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_42),
.C(n_44),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_69),
.Y(n_110)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_91),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_44),
.B(n_42),
.C(n_25),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_51),
.B(n_61),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_97),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_95),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_11),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_114),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_123),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_91),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_117),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_57),
.B1(n_48),
.B2(n_58),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_118),
.B1(n_89),
.B2(n_93),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_54),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_124),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_97),
.B(n_101),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_77),
.A2(n_6),
.B(n_7),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_122),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_8),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_8),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_10),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_10),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_13),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_135),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_82),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_148),
.B(n_117),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_112),
.B1(n_102),
.B2(n_105),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_80),
.A3(n_95),
.B1(n_92),
.B2(n_78),
.Y(n_134)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_124),
.A3(n_125),
.B1(n_110),
.B2(n_114),
.C1(n_118),
.C2(n_122),
.Y(n_151)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_105),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_121),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_73),
.A3(n_74),
.B1(n_86),
.B2(n_88),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_104),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_162),
.B(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_156),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_159),
.B(n_142),
.Y(n_169)
);

NAND2x1p5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_120),
.Y(n_155)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_147),
.B(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_142),
.B1(n_145),
.B2(n_138),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_106),
.B(n_73),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_107),
.C(n_113),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_163),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_133),
.B1(n_146),
.B2(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_137),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_169),
.A2(n_171),
.B(n_174),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_143),
.B(n_132),
.C(n_141),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_173),
.B1(n_157),
.B2(n_166),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_147),
.B(n_135),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_175),
.A2(n_176),
.B(n_156),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_127),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_181),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_121),
.B(n_136),
.Y(n_179)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_180),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_159),
.B(n_161),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_182),
.A2(n_187),
.B1(n_192),
.B2(n_173),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_160),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_186),
.C(n_170),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_164),
.B(n_158),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_153),
.B1(n_167),
.B2(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_193),
.B(n_179),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_177),
.C(n_170),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_196),
.C(n_199),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_181),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_182),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_158),
.C(n_175),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_201),
.B(n_185),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_207),
.B1(n_171),
.B2(n_195),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_209),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_191),
.C(n_197),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_205),
.B(n_152),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_211),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_214),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_210),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_182),
.Y(n_218)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_209),
.B(n_205),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_218),
.C(n_178),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_175),
.Y(n_220)
);


endmodule