module fake_jpeg_12719_n_454 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_454);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_454;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_6),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_52),
.B(n_61),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_53),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_55),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_57),
.Y(n_117)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_6),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_63),
.Y(n_104)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_65),
.Y(n_119)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_9),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_12),
.Y(n_106)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_72),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_29),
.A2(n_9),
.B1(n_13),
.B2(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_114)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_5),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_91),
.Y(n_110)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_89),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_95),
.Y(n_109)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_35),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_35),
.B1(n_26),
.B2(n_38),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_97),
.A2(n_114),
.B1(n_30),
.B2(n_42),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_106),
.B(n_115),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_34),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_50),
.A2(n_35),
.B1(n_42),
.B2(n_39),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_21),
.B1(n_42),
.B2(n_39),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_20),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_121),
.B(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_20),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_36),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_36),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_136),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_55),
.B(n_19),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_79),
.B(n_19),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_15),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_151),
.Y(n_230)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_155),
.A2(n_169),
.B1(n_171),
.B2(n_173),
.Y(n_206)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_157),
.A2(n_102),
.B1(n_133),
.B2(n_145),
.Y(n_211)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_110),
.A2(n_56),
.B1(n_53),
.B2(n_54),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_172),
.B1(n_119),
.B2(n_104),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_96),
.B(n_90),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_164),
.B(n_176),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_125),
.A2(n_88),
.B1(n_30),
.B2(n_28),
.Y(n_166)
);

OAI22x1_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_102),
.B1(n_117),
.B2(n_127),
.Y(n_209)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_118),
.A2(n_73),
.B1(n_84),
.B2(n_83),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_108),
.A2(n_82),
.B1(n_63),
.B2(n_65),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_110),
.A2(n_78),
.B1(n_59),
.B2(n_89),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_122),
.A2(n_35),
.B1(n_24),
.B2(n_30),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_132),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_177),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_98),
.B(n_0),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_178),
.A2(n_187),
.B1(n_191),
.B2(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_100),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_182),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_111),
.A2(n_15),
.B1(n_28),
.B2(n_27),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_22),
.B1(n_21),
.B2(n_27),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_109),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_128),
.B(n_0),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_194),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_185),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_186),
.B(n_22),
.Y(n_197)
);

BUFx6f_ASAP7_75t_SL g187 ( 
.A(n_141),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_113),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_129),
.B(n_15),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_195),
.Y(n_202)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_140),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_116),
.A2(n_23),
.B1(n_28),
.B2(n_27),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_192),
.A2(n_104),
.B1(n_119),
.B2(n_23),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_99),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_101),
.B(n_0),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_117),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_197),
.B(n_175),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_198),
.A2(n_211),
.B1(n_219),
.B2(n_221),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_203),
.B1(n_195),
.B2(n_24),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_209),
.A2(n_218),
.B(n_225),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_186),
.B(n_101),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_165),
.B(n_137),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_144),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_176),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_153),
.A2(n_126),
.B(n_120),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_157),
.A2(n_148),
.B1(n_112),
.B2(n_145),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_163),
.A2(n_105),
.B1(n_120),
.B2(n_148),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_174),
.A2(n_126),
.B1(n_107),
.B2(n_105),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_124),
.B1(n_127),
.B2(n_21),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_204),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_172),
.B1(n_169),
.B2(n_190),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_232),
.B1(n_240),
.B2(n_249),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_147),
.B1(n_135),
.B2(n_165),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_164),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_241),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_235),
.A2(n_215),
.B1(n_178),
.B2(n_159),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_207),
.A2(n_194),
.B(n_183),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_236),
.A2(n_239),
.B(n_243),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_237),
.Y(n_287)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_194),
.B(n_183),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_196),
.B1(n_212),
.B2(n_201),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_153),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_248),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_207),
.A2(n_153),
.B(n_164),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_244),
.A2(n_255),
.B(n_222),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_251),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_158),
.C(n_179),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_229),
.C(n_189),
.Y(n_268)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_158),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_196),
.A2(n_180),
.B1(n_182),
.B2(n_124),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_180),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_256),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_207),
.A2(n_181),
.B(n_168),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_208),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_210),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_152),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_208),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_263),
.B(n_283),
.Y(n_313)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_242),
.A3(n_248),
.B1(n_250),
.B2(n_240),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_201),
.B1(n_225),
.B2(n_200),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_265),
.A2(n_274),
.B1(n_289),
.B2(n_258),
.Y(n_299)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_270),
.C(n_276),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_209),
.C(n_224),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_258),
.A2(n_198),
.B1(n_203),
.B2(n_221),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_273),
.A2(n_231),
.B1(n_232),
.B2(n_249),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_231),
.A2(n_209),
.B1(n_171),
.B2(n_173),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_224),
.C(n_222),
.Y(n_276)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_259),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_277),
.Y(n_306)
);

A2O1A1O1Ixp25_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_255),
.B(n_239),
.C(n_234),
.D(n_235),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_241),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_236),
.B(n_170),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_234),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_256),
.Y(n_292)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_288),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_292),
.B(n_296),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_244),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_297),
.C(n_303),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_275),
.A2(n_243),
.B(n_259),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_299),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_267),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_244),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_302),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_300),
.A2(n_308),
.B1(n_254),
.B2(n_215),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_301),
.B(n_280),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_277),
.A2(n_243),
.B(n_255),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_236),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_304),
.B(n_305),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_279),
.Y(n_305)
);

OAI32xp33_ASAP7_75t_L g307 ( 
.A1(n_271),
.A2(n_272),
.A3(n_286),
.B1(n_262),
.B2(n_283),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_177),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_273),
.A2(n_232),
.B1(n_234),
.B2(n_239),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_287),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_251),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_268),
.B(n_257),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_315),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_245),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_314),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_253),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_269),
.B(n_252),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_199),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_237),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_284),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_323),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_309),
.A2(n_262),
.B1(n_275),
.B2(n_274),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_320),
.A2(n_331),
.B1(n_337),
.B2(n_339),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_278),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_270),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_326),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_282),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_294),
.Y(n_329)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_329),
.Y(n_353)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_296),
.Y(n_330)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_330),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_309),
.A2(n_289),
.B1(n_288),
.B2(n_266),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_306),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_344),
.Y(n_352)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

XNOR2x1_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_341),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_300),
.A2(n_266),
.B1(n_281),
.B2(n_254),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_313),
.B(n_199),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_193),
.Y(n_367)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_307),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_304),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_308),
.A2(n_223),
.B1(n_161),
.B2(n_230),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_345),
.A2(n_223),
.B1(n_230),
.B2(n_226),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g346 ( 
.A(n_327),
.B(n_297),
.CI(n_301),
.CON(n_346),
.SN(n_346)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_360),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_323),
.C(n_327),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_354),
.C(n_356),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_338),
.A2(n_302),
.B(n_295),
.Y(n_350)
);

XOR2x2_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_162),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_340),
.B(n_293),
.C(n_315),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_355),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_342),
.C(n_326),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_316),
.C(n_303),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_357),
.B(n_167),
.C(n_191),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_324),
.A2(n_332),
.B1(n_306),
.B2(n_321),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_359),
.A2(n_362),
.B1(n_364),
.B2(n_344),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_322),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_320),
.A2(n_161),
.B1(n_230),
.B2(n_162),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_205),
.Y(n_366)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_366),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_335),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_318),
.B(n_226),
.Y(n_368)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_156),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_336),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_370),
.A2(n_381),
.B1(n_388),
.B2(n_363),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_361),
.B(n_337),
.Y(n_374)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_374),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_352),
.A2(n_336),
.B(n_334),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_376),
.Y(n_404)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_358),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_382),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_336),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_378),
.B(n_184),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_359),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_383),
.B(n_369),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_351),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_365),
.C(n_351),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_385),
.B(n_386),
.Y(n_399)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_365),
.B(n_135),
.C(n_147),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_363),
.C(n_364),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_366),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_393),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_402),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_356),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_357),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_396),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_373),
.A2(n_350),
.B(n_352),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_395),
.A2(n_384),
.B(n_374),
.Y(n_412)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_397),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_371),
.A2(n_353),
.B1(n_347),
.B2(n_346),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_400),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_347),
.B1(n_346),
.B2(n_367),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_187),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_401),
.B(n_403),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_185),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_116),
.C(n_160),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_151),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_399),
.B(n_380),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_417),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_387),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_409),
.B(n_419),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_412),
.A2(n_392),
.B(n_24),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_389),
.A2(n_372),
.B1(n_381),
.B2(n_376),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_413),
.B(n_415),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_404),
.A2(n_396),
.B1(n_403),
.B2(n_383),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_382),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_377),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_418),
.B(n_11),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_406),
.A2(n_402),
.B(n_392),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_425),
.B(n_12),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_391),
.Y(n_422)
);

AOI21xp33_ASAP7_75t_L g437 ( 
.A1(n_422),
.A2(n_12),
.B(n_3),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_12),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_410),
.A2(n_141),
.B(n_23),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_409),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_426),
.B(n_428),
.C(n_408),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_427),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_410),
.C(n_414),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_11),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_430),
.B(n_431),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_408),
.B(n_10),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_434),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_423),
.A2(n_419),
.B1(n_17),
.B2(n_37),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_435),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_437),
.Y(n_444)
);

XOR2x2_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_4),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_439),
.C(n_429),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_4),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_438),
.A2(n_429),
.B(n_37),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_445),
.Y(n_447)
);

A2O1A1O1Ixp25_ASAP7_75t_L g446 ( 
.A1(n_442),
.A2(n_433),
.B(n_440),
.C(n_436),
.D(n_37),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_446),
.A2(n_448),
.B(n_444),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_17),
.C(n_5),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_449),
.A2(n_450),
.B(n_14),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_447),
.A2(n_14),
.B(n_5),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_451),
.B(n_14),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_1),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_1),
.B(n_445),
.Y(n_454)
);


endmodule