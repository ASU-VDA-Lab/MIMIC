module fake_netlist_5_1981_n_1591 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_1591);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1591;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_144;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1565;
wire n_182;
wire n_143;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_146;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_338;
wire n_149;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_148;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_147;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_145;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_60),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_5),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_75),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_35),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_26),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_59),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_53),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_62),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_32),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_57),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_113),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_70),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_84),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_5),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_66),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_37),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_63),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_68),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_39),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_39),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_48),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_47),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_46),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_12),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_61),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_6),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_3),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_41),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_103),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_86),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_43),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_41),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_14),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_31),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_37),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_11),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_109),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_98),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_24),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_91),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_25),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_22),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_12),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_141),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_99),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_38),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_1),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_30),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_35),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_31),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_51),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_4),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_94),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_21),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_65),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_112),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_10),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_11),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_88),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_130),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_114),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_40),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_137),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_58),
.Y(n_225)
);

BUFx2_ASAP7_75t_SL g226 ( 
.A(n_90),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_93),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_67),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_46),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_138),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_0),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_116),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_4),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_14),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_97),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_102),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_139),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_126),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_89),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_96),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_33),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_45),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g243 ( 
.A(n_34),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_18),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_127),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_19),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_32),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_56),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_36),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_30),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_82),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_77),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_27),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_123),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_64),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_133),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_6),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_110),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_71),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_38),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_23),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_50),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_40),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_115),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_23),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_22),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_45),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_124),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_2),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_25),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_2),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_78),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_9),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_119),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_17),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_118),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_0),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_128),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_17),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_120),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_145),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_174),
.B(n_1),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_203),
.B(n_3),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_164),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_245),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_184),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_191),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_179),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_164),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_179),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_147),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_169),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_191),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_191),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_191),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_191),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_167),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_7),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_169),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_173),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_219),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_177),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_188),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_148),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_152),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_230),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_207),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_227),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_209),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_213),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_151),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_229),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_182),
.Y(n_315)
);

BUFx6f_ASAP7_75t_SL g316 ( 
.A(n_252),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_189),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_190),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_196),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_205),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_247),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_233),
.B(n_7),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_157),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_185),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_185),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_197),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_203),
.B(n_8),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_199),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_157),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_201),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_202),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_150),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_197),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_206),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_163),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_276),
.B(n_8),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_267),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_272),
.B(n_9),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_269),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_163),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_268),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_210),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_268),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_277),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_218),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_227),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_223),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_222),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_231),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_143),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_234),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_144),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_241),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_287),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_287),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_295),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_286),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_281),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_306),
.B(n_146),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_298),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_299),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_307),
.B(n_291),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_291),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_304),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_313),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_305),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_313),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_309),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_310),
.B(n_150),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_315),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_311),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_315),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_312),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_314),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_320),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_285),
.B(n_214),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_316),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_317),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_336),
.B(n_214),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_331),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_283),
.A2(n_232),
.B(n_156),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_332),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_342),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_344),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_288),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_290),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_293),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_351),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_294),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_317),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_323),
.B(n_232),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_318),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_321),
.B(n_233),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_282),
.B(n_176),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_319),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_330),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_300),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_340),
.A2(n_159),
.B(n_153),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_303),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_334),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_334),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_335),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_335),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_338),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_347),
.B(n_165),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_350),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_361),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_412),
.A2(n_393),
.B1(n_414),
.B2(n_406),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_324),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_350),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_390),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_401),
.Y(n_435)
);

BUFx10_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_352),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_397),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_308),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_417),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_417),
.B(n_324),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_391),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_401),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_406),
.B(n_414),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_402),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_411),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_361),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_366),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_406),
.B(n_412),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_352),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_333),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_419),
.Y(n_454)
);

AND3x1_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_246),
.C(n_215),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_393),
.A2(n_215),
.B1(n_244),
.B2(n_273),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_429),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_368),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_402),
.Y(n_460)
);

AO22x2_ASAP7_75t_L g461 ( 
.A1(n_425),
.A2(n_246),
.B1(n_149),
.B2(n_273),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_403),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_373),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_419),
.B(n_354),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_368),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_418),
.B(n_158),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_418),
.B(n_158),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_375),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_360),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_397),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_364),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_393),
.B(n_354),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_409),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_418),
.B(n_158),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_388),
.B(n_356),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_425),
.B(n_333),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_360),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_362),
.Y(n_479)
);

AND2x2_ASAP7_75t_SL g480 ( 
.A(n_409),
.B(n_158),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_393),
.B(n_178),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_405),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_409),
.B(n_356),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_369),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_427),
.B(n_339),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_362),
.B(n_358),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_418),
.B(n_178),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_L g492 ( 
.A(n_408),
.B(n_178),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_404),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_369),
.Y(n_494)
);

OR2x6_ASAP7_75t_L g495 ( 
.A(n_363),
.B(n_226),
.Y(n_495)
);

AO22x2_ASAP7_75t_L g496 ( 
.A1(n_404),
.A2(n_244),
.B1(n_149),
.B2(n_243),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_371),
.Y(n_497)
);

NAND2xp33_ASAP7_75t_L g498 ( 
.A(n_377),
.B(n_178),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_371),
.B(n_178),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_382),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_374),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_374),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_376),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_363),
.B(n_200),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_372),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_380),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_365),
.B(n_339),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_359),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_378),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_381),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_381),
.B(n_166),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_383),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_370),
.B(n_187),
.Y(n_514)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_372),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_365),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_383),
.B(n_170),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_385),
.B(n_395),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_394),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_384),
.B(n_386),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_394),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_395),
.Y(n_523)
);

BUFx4f_ASAP7_75t_L g524 ( 
.A(n_395),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_386),
.B(n_387),
.Y(n_525)
);

INVx5_ASAP7_75t_L g526 ( 
.A(n_396),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_392),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_398),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_407),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_389),
.B(n_187),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_399),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_400),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_400),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_396),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_410),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_396),
.B(n_171),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_415),
.B(n_353),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_416),
.B(n_224),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_422),
.A2(n_187),
.B1(n_235),
.B2(n_254),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_426),
.Y(n_541)
);

INVx3_ASAP7_75t_R g542 ( 
.A(n_423),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_424),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_361),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_363),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_390),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_367),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_411),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_390),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_390),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_411),
.B(n_183),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_361),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_379),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_367),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_397),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_413),
.B(n_316),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_390),
.Y(n_557)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_397),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_390),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_397),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_442),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_553),
.B(n_175),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_432),
.B(n_284),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_441),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_431),
.B(n_204),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_444),
.B(n_180),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_493),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_480),
.B(n_187),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_432),
.A2(n_348),
.B1(n_346),
.B2(n_337),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_449),
.B(n_198),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_480),
.B(n_187),
.Y(n_572)
);

OAI22x1_ASAP7_75t_SL g573 ( 
.A1(n_464),
.A2(n_193),
.B1(n_265),
.B2(n_192),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_503),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_446),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_440),
.B(n_211),
.Y(n_576)
);

O2A1O1Ixp33_ASAP7_75t_L g577 ( 
.A1(n_440),
.A2(n_248),
.B(n_280),
.C(n_274),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_548),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_431),
.B(n_225),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_433),
.B(n_154),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_437),
.B(n_154),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_452),
.A2(n_238),
.B1(n_258),
.B2(n_236),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_465),
.B(n_204),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_430),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_441),
.B(n_155),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_L g586 ( 
.A(n_481),
.B(n_204),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_524),
.B(n_204),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_453),
.A2(n_328),
.B1(n_327),
.B2(n_326),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_450),
.B(n_181),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_528),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_482),
.B(n_160),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_476),
.B(n_160),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_453),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_528),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_470),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_458),
.B(n_161),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_532),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_470),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_478),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_474),
.B(n_186),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_532),
.Y(n_601)
);

NAND2x1_ASAP7_75t_L g602 ( 
.A(n_462),
.B(n_49),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_439),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_524),
.B(n_451),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_435),
.Y(n_605)
);

INVx8_ASAP7_75t_L g606 ( 
.A(n_495),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_503),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_488),
.B(n_494),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_473),
.B(n_161),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_438),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_501),
.B(n_502),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_510),
.Y(n_612)
);

BUFx8_ASAP7_75t_L g613 ( 
.A(n_545),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_451),
.B(n_204),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_443),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_542),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_445),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_454),
.B(n_204),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_518),
.A2(n_194),
.B(n_195),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_507),
.B(n_289),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_511),
.B(n_513),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_454),
.B(n_204),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_460),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_477),
.B(n_489),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_544),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_477),
.B(n_249),
.C(n_250),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_497),
.B(n_292),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_544),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_463),
.Y(n_629)
);

NOR2x1p5_ASAP7_75t_L g630 ( 
.A(n_534),
.B(n_208),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_483),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_531),
.B(n_533),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_497),
.B(n_301),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_504),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_560),
.B(n_212),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_510),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_560),
.B(n_216),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_489),
.B(n_162),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_438),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_482),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_508),
.B(n_265),
.Y(n_641)
);

INVx6_ASAP7_75t_L g642 ( 
.A(n_534),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_552),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_487),
.B(n_162),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_484),
.Y(n_645)
);

AND2x6_ASAP7_75t_SL g646 ( 
.A(n_535),
.B(n_172),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_538),
.B(n_509),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_434),
.B(n_168),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_546),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_552),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_469),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_506),
.B(n_256),
.Y(n_652)
);

NOR2xp67_ASAP7_75t_L g653 ( 
.A(n_526),
.B(n_251),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_512),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_540),
.A2(n_168),
.B1(n_278),
.B2(n_239),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_534),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_549),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_519),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_457),
.A2(n_172),
.B1(n_192),
.B2(n_193),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_523),
.B(n_262),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_512),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_479),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_521),
.B(n_228),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_556),
.A2(n_264),
.B1(n_240),
.B2(n_217),
.Y(n_664)
);

O2A1O1Ixp5_ASAP7_75t_L g665 ( 
.A1(n_505),
.A2(n_255),
.B(n_237),
.C(n_220),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_521),
.B(n_221),
.Y(n_666)
);

AND2x2_ASAP7_75t_SL g667 ( 
.A(n_540),
.B(n_252),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_525),
.B(n_278),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_556),
.B(n_257),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g670 ( 
.A(n_526),
.B(n_74),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_523),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_522),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_522),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_550),
.B(n_252),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_534),
.B(n_10),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_520),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_448),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_490),
.B(n_279),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_508),
.B(n_275),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_448),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_523),
.B(n_275),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_479),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_557),
.B(n_271),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_559),
.B(n_271),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_500),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_457),
.B(n_270),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_436),
.B(n_208),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_523),
.B(n_55),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_517),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_527),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_456),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_516),
.B(n_69),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_517),
.Y(n_693)
);

BUFx6f_ASAP7_75t_SL g694 ( 
.A(n_527),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_436),
.B(n_13),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_547),
.B(n_15),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_526),
.B(n_72),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_547),
.B(n_15),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_561),
.B(n_486),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_455),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_456),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_459),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_496),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_554),
.B(n_16),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_459),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_554),
.B(n_16),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_466),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_624),
.A2(n_593),
.B1(n_580),
.B2(n_581),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_595),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_624),
.A2(n_467),
.B(n_491),
.C(n_468),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_580),
.B(n_505),
.Y(n_711)
);

BUFx4f_ASAP7_75t_L g712 ( 
.A(n_606),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_574),
.B(n_636),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_627),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_604),
.A2(n_558),
.B(n_462),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_565),
.B(n_529),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_634),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_662),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_604),
.A2(n_558),
.B(n_471),
.Y(n_719)
);

AND2x6_ASAP7_75t_L g720 ( 
.A(n_671),
.B(n_543),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_651),
.B(n_526),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_671),
.A2(n_471),
.B(n_475),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_576),
.B(n_475),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_607),
.B(n_467),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_620),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_656),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_659),
.A2(n_496),
.B1(n_461),
.B2(n_495),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_671),
.A2(n_555),
.B(n_485),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_671),
.A2(n_555),
.B(n_485),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_574),
.B(n_539),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_607),
.B(n_481),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_SL g732 ( 
.A1(n_644),
.A2(n_486),
.B(n_498),
.C(n_492),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_679),
.A2(n_514),
.B(n_530),
.C(n_541),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_585),
.B(n_481),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_662),
.Y(n_735)
);

BUFx8_ASAP7_75t_L g736 ( 
.A(n_694),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_585),
.B(n_481),
.Y(n_737)
);

BUFx4f_ASAP7_75t_L g738 ( 
.A(n_606),
.Y(n_738)
);

AO21x1_ASAP7_75t_L g739 ( 
.A1(n_688),
.A2(n_587),
.B(n_635),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_574),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_595),
.Y(n_741)
);

NAND3xp33_ASAP7_75t_L g742 ( 
.A(n_638),
.B(n_514),
.C(n_530),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_638),
.A2(n_495),
.B1(n_481),
.B2(n_541),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_609),
.B(n_496),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_633),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_659),
.A2(n_461),
.B1(n_536),
.B2(n_537),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_614),
.A2(n_555),
.B(n_438),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_636),
.B(n_485),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_618),
.A2(n_485),
.B(n_466),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_618),
.A2(n_447),
.B(n_515),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_609),
.B(n_461),
.Y(n_751)
);

O2A1O1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_681),
.A2(n_703),
.B(n_579),
.C(n_562),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_598),
.Y(n_753)
);

AOI21x1_ASAP7_75t_L g754 ( 
.A1(n_587),
.A2(n_536),
.B(n_515),
.Y(n_754)
);

AOI21x1_ASAP7_75t_L g755 ( 
.A1(n_622),
.A2(n_499),
.B(n_79),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_681),
.A2(n_19),
.B(n_20),
.C(n_24),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_682),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_647),
.B(n_687),
.Y(n_758)
);

O2A1O1Ixp5_ASAP7_75t_L g759 ( 
.A1(n_665),
.A2(n_499),
.B(n_81),
.C(n_85),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_613),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_636),
.B(n_499),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_663),
.B(n_499),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_666),
.B(n_499),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_622),
.A2(n_54),
.B(n_129),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_687),
.B(n_592),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_660),
.A2(n_52),
.B(n_122),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_660),
.A2(n_131),
.B(n_121),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_575),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_685),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_678),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_770)
);

BUFx12f_ASAP7_75t_L g771 ( 
.A(n_613),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_668),
.B(n_28),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_563),
.B(n_29),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_612),
.B(n_80),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_699),
.A2(n_87),
.B(n_105),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_641),
.B(n_34),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_644),
.B(n_36),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_678),
.B(n_42),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_610),
.A2(n_95),
.B(n_101),
.Y(n_779)
);

O2A1O1Ixp5_ASAP7_75t_L g780 ( 
.A1(n_569),
.A2(n_44),
.B(n_572),
.C(n_637),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_599),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_667),
.A2(n_686),
.B1(n_700),
.B2(n_688),
.Y(n_782)
);

BUFx6f_ASAP7_75t_L g783 ( 
.A(n_656),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_667),
.A2(n_44),
.B1(n_700),
.B2(n_592),
.Y(n_784)
);

AOI22x1_ASAP7_75t_L g785 ( 
.A1(n_605),
.A2(n_623),
.B1(n_629),
.B2(n_615),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_640),
.B(n_617),
.Y(n_786)
);

NOR2x1_ASAP7_75t_L g787 ( 
.A(n_690),
.B(n_626),
.Y(n_787)
);

AND2x2_ASAP7_75t_SL g788 ( 
.A(n_564),
.B(n_570),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_642),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_639),
.A2(n_583),
.B(n_652),
.Y(n_790)
);

INVx5_ASAP7_75t_L g791 ( 
.A(n_642),
.Y(n_791)
);

INVx5_ASAP7_75t_L g792 ( 
.A(n_642),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_603),
.B(n_669),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_631),
.B(n_645),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_608),
.B(n_611),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_635),
.A2(n_637),
.B(n_571),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_588),
.B(n_706),
.C(n_696),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_578),
.B(n_596),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_621),
.A2(n_632),
.B(n_567),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_569),
.A2(n_572),
.B(n_566),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_589),
.A2(n_600),
.B(n_619),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_577),
.A2(n_649),
.B(n_657),
.C(n_601),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_702),
.Y(n_803)
);

AOI21x1_ASAP7_75t_L g804 ( 
.A1(n_590),
.A2(n_594),
.B(n_597),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_612),
.B(n_661),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_602),
.Y(n_806)
);

OAI21xp33_ASAP7_75t_L g807 ( 
.A1(n_683),
.A2(n_684),
.B(n_706),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_696),
.B(n_698),
.Y(n_808)
);

NOR3xp33_ASAP7_75t_L g809 ( 
.A(n_698),
.B(n_695),
.C(n_704),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_591),
.B(n_654),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_648),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_692),
.A2(n_707),
.B(n_702),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_689),
.B(n_693),
.Y(n_813)
);

AOI21xp33_ASAP7_75t_L g814 ( 
.A1(n_582),
.A2(n_655),
.B(n_701),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_591),
.B(n_664),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_707),
.A2(n_705),
.B(n_691),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_676),
.B(n_568),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_658),
.B(n_673),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_648),
.A2(n_672),
.B1(n_677),
.B2(n_680),
.Y(n_819)
);

AO22x1_ASAP7_75t_L g820 ( 
.A1(n_674),
.A2(n_675),
.B1(n_646),
.B2(n_573),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_L g821 ( 
.A(n_586),
.B(n_584),
.C(n_650),
.Y(n_821)
);

OAI22xp33_ASAP7_75t_SL g822 ( 
.A1(n_675),
.A2(n_625),
.B1(n_643),
.B2(n_628),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_675),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_653),
.B(n_670),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_630),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_697),
.A2(n_606),
.B(n_620),
.Y(n_826)
);

AND2x2_ASAP7_75t_SL g827 ( 
.A(n_616),
.B(n_620),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_624),
.B(n_565),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_624),
.B(n_565),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_574),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_604),
.A2(n_524),
.B(n_671),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_593),
.B(n_442),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_624),
.B(n_565),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_574),
.Y(n_834)
);

AOI21xp33_ASAP7_75t_L g835 ( 
.A1(n_624),
.A2(n_432),
.B(n_585),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_624),
.B(n_444),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_587),
.A2(n_618),
.B(n_614),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_624),
.B(n_444),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_624),
.B(n_444),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_699),
.A2(n_618),
.B(n_614),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_604),
.A2(n_524),
.B(n_671),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_593),
.B(n_442),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_662),
.Y(n_843)
);

OAI21xp33_ASAP7_75t_L g844 ( 
.A1(n_679),
.A2(n_624),
.B(n_432),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_624),
.B(n_444),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_604),
.A2(n_524),
.B(n_671),
.Y(n_846)
);

OAI21xp33_ASAP7_75t_L g847 ( 
.A1(n_679),
.A2(n_624),
.B(n_432),
.Y(n_847)
);

CKINVDCx6p67_ASAP7_75t_R g848 ( 
.A(n_694),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_671),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_604),
.A2(n_524),
.B(n_671),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_595),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_624),
.B(n_444),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_604),
.A2(n_524),
.B(n_518),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_624),
.B(n_444),
.Y(n_854)
);

OAI321xp33_ASAP7_75t_L g855 ( 
.A1(n_624),
.A2(n_679),
.A3(n_565),
.B1(n_585),
.B2(n_417),
.C(n_576),
.Y(n_855)
);

NAND2x1p5_ASAP7_75t_L g856 ( 
.A(n_671),
.B(n_656),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_L g857 ( 
.A(n_651),
.B(n_526),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_595),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_574),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_624),
.B(n_444),
.Y(n_860)
);

AND2x2_ASAP7_75t_SL g861 ( 
.A(n_659),
.B(n_667),
.Y(n_861)
);

AOI21x1_ASAP7_75t_L g862 ( 
.A1(n_587),
.A2(n_618),
.B(n_614),
.Y(n_862)
);

INVx11_ASAP7_75t_L g863 ( 
.A(n_613),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_604),
.A2(n_524),
.B(n_518),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_662),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_595),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_835),
.B(n_708),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_768),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_849),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_803),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_804),
.A2(n_749),
.B(n_747),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_715),
.A2(n_719),
.B(n_831),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_832),
.B(n_842),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_841),
.A2(n_850),
.B(n_846),
.Y(n_875)
);

BUFx10_ASAP7_75t_L g876 ( 
.A(n_716),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_718),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_L g878 ( 
.A(n_765),
.B(n_847),
.C(n_844),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_849),
.Y(n_879)
);

INVx6_ASAP7_75t_SL g880 ( 
.A(n_805),
.Y(n_880)
);

AOI21xp33_ASAP7_75t_L g881 ( 
.A1(n_855),
.A2(n_861),
.B(n_778),
.Y(n_881)
);

OAI21x1_ASAP7_75t_L g882 ( 
.A1(n_722),
.A2(n_729),
.B(n_728),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_758),
.B(n_828),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_788),
.A2(n_829),
.B1(n_833),
.B2(n_808),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_801),
.A2(n_862),
.B(n_837),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_714),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_735),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_836),
.A2(n_839),
.B(n_838),
.Y(n_888)
);

OA21x2_ASAP7_75t_L g889 ( 
.A1(n_853),
.A2(n_864),
.B(n_800),
.Y(n_889)
);

OAI21x1_ASAP7_75t_L g890 ( 
.A1(n_816),
.A2(n_864),
.B(n_750),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_784),
.A2(n_782),
.B1(n_797),
.B2(n_777),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_714),
.Y(n_892)
);

AO21x2_ASAP7_75t_L g893 ( 
.A1(n_711),
.A2(n_737),
.B(n_734),
.Y(n_893)
);

AOI21xp33_ASAP7_75t_L g894 ( 
.A1(n_784),
.A2(n_782),
.B(n_772),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_785),
.A2(n_754),
.B(n_755),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_845),
.B(n_852),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_791),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_805),
.B(n_811),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_800),
.A2(n_724),
.B(n_748),
.Y(n_899)
);

AO31x2_ASAP7_75t_L g900 ( 
.A1(n_744),
.A2(n_802),
.A3(n_751),
.B(n_860),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_854),
.B(n_807),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_757),
.A2(n_865),
.B(n_843),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_752),
.A2(n_742),
.B(n_793),
.C(n_780),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_798),
.B(n_723),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_745),
.Y(n_905)
);

INVx5_ASAP7_75t_L g906 ( 
.A(n_720),
.Y(n_906)
);

OA21x2_ASAP7_75t_L g907 ( 
.A1(n_759),
.A2(n_762),
.B(n_763),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_709),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_794),
.B(n_741),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_710),
.A2(n_742),
.B(n_814),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_815),
.A2(n_824),
.B(n_731),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_745),
.Y(n_912)
);

AO21x2_ASAP7_75t_L g913 ( 
.A1(n_732),
.A2(n_814),
.B(n_809),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_753),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_713),
.A2(n_821),
.B(n_818),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_781),
.B(n_866),
.Y(n_916)
);

AOI211x1_ASAP7_75t_L g917 ( 
.A1(n_727),
.A2(n_746),
.B(n_776),
.C(n_820),
.Y(n_917)
);

AOI221xp5_ASAP7_75t_L g918 ( 
.A1(n_770),
.A2(n_746),
.B1(n_727),
.B2(n_756),
.C(n_773),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_851),
.B(n_858),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_743),
.A2(n_810),
.B(n_819),
.C(n_786),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_823),
.B(n_769),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_821),
.A2(n_817),
.B(n_822),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_740),
.B(n_834),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_740),
.B(n_834),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_856),
.A2(n_767),
.B(n_766),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_856),
.A2(n_859),
.B(n_830),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_787),
.A2(n_730),
.B1(n_813),
.B2(n_825),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_830),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_725),
.Y(n_929)
);

AOI21x1_ASAP7_75t_L g930 ( 
.A1(n_761),
.A2(n_774),
.B(n_764),
.Y(n_930)
);

CKINVDCx6p67_ASAP7_75t_R g931 ( 
.A(n_760),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_827),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_859),
.A2(n_775),
.B(n_779),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_822),
.A2(n_806),
.B(n_792),
.Y(n_934)
);

NOR2x1_ASAP7_75t_L g935 ( 
.A(n_721),
.B(n_857),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_792),
.A2(n_806),
.B(n_726),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_806),
.A2(n_720),
.B(n_792),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_720),
.A2(n_789),
.B(n_726),
.Y(n_938)
);

CKINVDCx16_ASAP7_75t_R g939 ( 
.A(n_771),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_783),
.A2(n_712),
.B(n_738),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_720),
.A2(n_712),
.B(n_738),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_783),
.B(n_789),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_848),
.B(n_736),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_863),
.B(n_736),
.Y(n_944)
);

OAI21x1_ASAP7_75t_L g945 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_714),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_769),
.Y(n_949)
);

AOI21x1_ASAP7_75t_L g950 ( 
.A1(n_804),
.A2(n_660),
.B(n_587),
.Y(n_950)
);

OAI21xp33_ASAP7_75t_L g951 ( 
.A1(n_844),
.A2(n_624),
.B(n_432),
.Y(n_951)
);

AO31x2_ASAP7_75t_L g952 ( 
.A1(n_739),
.A2(n_733),
.A3(n_782),
.B(n_711),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_836),
.B(n_838),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_799),
.A2(n_671),
.B(n_604),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_835),
.B(n_844),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_832),
.B(n_842),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_799),
.A2(n_796),
.B(n_795),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_768),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_804),
.A2(n_660),
.B(n_587),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_714),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_836),
.B(n_838),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_849),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_835),
.B(n_708),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_836),
.B(n_838),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_832),
.B(n_842),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_836),
.B(n_838),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_799),
.A2(n_796),
.B(n_795),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_718),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_836),
.B(n_838),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_805),
.B(n_811),
.Y(n_972)
);

AOI21x1_ASAP7_75t_L g973 ( 
.A1(n_804),
.A2(n_660),
.B(n_587),
.Y(n_973)
);

OAI21xp33_ASAP7_75t_L g974 ( 
.A1(n_844),
.A2(n_624),
.B(n_432),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_826),
.B(n_606),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_726),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_SL g978 ( 
.A(n_861),
.B(n_784),
.Y(n_978)
);

OR2x2_ASAP7_75t_L g979 ( 
.A(n_714),
.B(n_472),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_835),
.B(n_708),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_768),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_983)
);

AOI21x1_ASAP7_75t_L g984 ( 
.A1(n_804),
.A2(n_660),
.B(n_587),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_799),
.A2(n_671),
.B(n_604),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_835),
.A2(n_864),
.B(n_853),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_799),
.A2(n_796),
.B(n_795),
.Y(n_987)
);

AO31x2_ASAP7_75t_L g988 ( 
.A1(n_739),
.A2(n_733),
.A3(n_782),
.B(n_711),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_812),
.A2(n_840),
.B(n_790),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_791),
.B(n_792),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_836),
.B(n_838),
.Y(n_991)
);

AOI21x1_ASAP7_75t_L g992 ( 
.A1(n_804),
.A2(n_660),
.B(n_587),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_717),
.Y(n_993)
);

INVx5_ASAP7_75t_L g994 ( 
.A(n_906),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_979),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_883),
.B(n_896),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_940),
.B(n_975),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_874),
.B(n_958),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_978),
.A2(n_951),
.B1(n_974),
.B2(n_956),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_977),
.Y(n_1000)
);

AO221x2_ASAP7_75t_L g1001 ( 
.A1(n_878),
.A2(n_978),
.B1(n_910),
.B2(n_986),
.C(n_884),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_912),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_967),
.B(n_886),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_886),
.B(n_892),
.Y(n_1004)
);

BUFx10_ASAP7_75t_L g1005 ( 
.A(n_944),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_887),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_892),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_SL g1008 ( 
.A1(n_876),
.A2(n_905),
.B1(n_962),
.B2(n_947),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_905),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_897),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_959),
.A2(n_987),
.B(n_969),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_868),
.B(n_965),
.Y(n_1012)
);

NAND2x1p5_ASAP7_75t_L g1013 ( 
.A(n_897),
.B(n_906),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_940),
.B(n_975),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_932),
.B(n_891),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_896),
.B(n_953),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_L g1017 ( 
.A(n_894),
.B(n_980),
.C(n_918),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_876),
.B(n_921),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_954),
.A2(n_985),
.B(n_888),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_949),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_894),
.A2(n_991),
.B1(n_966),
.B2(n_971),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_953),
.A2(n_971),
.B1(n_963),
.B2(n_991),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_939),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_888),
.A2(n_911),
.B(n_968),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_911),
.A2(n_968),
.B(n_966),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_904),
.B(n_993),
.Y(n_1026)
);

OR2x6_ASAP7_75t_L g1027 ( 
.A(n_941),
.B(n_990),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_910),
.A2(n_904),
.B(n_903),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_929),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_941),
.B(n_990),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_880),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_869),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_970),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_975),
.B(n_960),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_901),
.A2(n_920),
.B1(n_917),
.B2(n_918),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_977),
.Y(n_1036)
);

OR2x6_ASAP7_75t_L g1037 ( 
.A(n_981),
.B(n_943),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_881),
.A2(n_898),
.B1(n_972),
.B2(n_913),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_908),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_SL g1040 ( 
.A1(n_906),
.A2(n_972),
.B1(n_898),
.B2(n_901),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_909),
.B(n_900),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_931),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_977),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_913),
.A2(n_986),
.B1(n_914),
.B2(n_880),
.Y(n_1044)
);

NAND2xp33_ASAP7_75t_L g1045 ( 
.A(n_906),
.B(n_935),
.Y(n_1045)
);

INVx5_ASAP7_75t_L g1046 ( 
.A(n_870),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_942),
.B(n_927),
.Y(n_1047)
);

AO31x2_ASAP7_75t_L g1048 ( 
.A1(n_922),
.A2(n_915),
.A3(n_934),
.B(n_952),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_900),
.B(n_942),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_871),
.Y(n_1050)
);

OR2x6_ASAP7_75t_L g1051 ( 
.A(n_936),
.B(n_937),
.Y(n_1051)
);

INVx3_ASAP7_75t_SL g1052 ( 
.A(n_870),
.Y(n_1052)
);

INVx3_ASAP7_75t_SL g1053 ( 
.A(n_879),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_879),
.B(n_964),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_900),
.B(n_919),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_964),
.B(n_938),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_926),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_915),
.A2(n_885),
.B(n_873),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_893),
.A2(n_925),
.B(n_875),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_928),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_923),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_924),
.B(n_952),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_952),
.B(n_988),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_988),
.B(n_893),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_988),
.B(n_889),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_899),
.Y(n_1066)
);

OR2x6_ASAP7_75t_L g1067 ( 
.A(n_930),
.B(n_933),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_907),
.B(n_890),
.Y(n_1068)
);

OA21x2_ASAP7_75t_L g1069 ( 
.A1(n_867),
.A2(n_957),
.B(n_989),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_895),
.A2(n_955),
.B(n_983),
.C(n_982),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_882),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_950),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_961),
.B(n_992),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_872),
.B(n_948),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_973),
.B(n_984),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_945),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_L g1077 ( 
.A(n_976),
.B(n_946),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_951),
.A2(n_835),
.B(n_847),
.C(n_844),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_883),
.B(n_828),
.Y(n_1079)
);

OAI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_891),
.A2(n_624),
.B(n_844),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_L g1081 ( 
.A(n_949),
.B(n_769),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_902),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_993),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_880),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_877),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_877),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_979),
.Y(n_1087)
);

AND2x6_ASAP7_75t_L g1088 ( 
.A(n_870),
.B(n_879),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_883),
.B(n_828),
.Y(n_1089)
);

O2A1O1Ixp5_ASAP7_75t_L g1090 ( 
.A1(n_881),
.A2(n_835),
.B(n_765),
.C(n_808),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_886),
.Y(n_1091)
);

AOI21xp33_ASAP7_75t_SL g1092 ( 
.A1(n_932),
.A2(n_432),
.B(n_624),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_979),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_978),
.A2(n_765),
.B1(n_564),
.B2(n_844),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_877),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_883),
.B(n_828),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_884),
.B(n_835),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_906),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_916),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_977),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_951),
.A2(n_835),
.B(n_847),
.C(n_844),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_949),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_902),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_993),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_978),
.A2(n_765),
.B1(n_564),
.B2(n_844),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_949),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_940),
.B(n_975),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_874),
.B(n_958),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_906),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_874),
.B(n_958),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_874),
.B(n_958),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_883),
.B(n_828),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_883),
.B(n_828),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_874),
.B(n_958),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_979),
.B(n_472),
.Y(n_1115)
);

BUFx2_ASAP7_75t_R g1116 ( 
.A(n_1102),
.Y(n_1116)
);

CKINVDCx11_ASAP7_75t_R g1117 ( 
.A(n_1023),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1097),
.B(n_1092),
.Y(n_1118)
);

INVxp67_ASAP7_75t_L g1119 ( 
.A(n_1009),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1094),
.A2(n_1105),
.B1(n_1016),
.B2(n_996),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1049),
.Y(n_1121)
);

INVx11_ASAP7_75t_L g1122 ( 
.A(n_1020),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1006),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1080),
.A2(n_1017),
.B1(n_1001),
.B2(n_1012),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_1001),
.A2(n_1015),
.B1(n_1035),
.B2(n_999),
.Y(n_1125)
);

INVx6_ASAP7_75t_L g1126 ( 
.A(n_994),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_1042),
.Y(n_1127)
);

BUFx2_ASAP7_75t_SL g1128 ( 
.A(n_1081),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1028),
.A2(n_1022),
.B1(n_1021),
.B2(n_1079),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_1070),
.A2(n_1019),
.B(n_1011),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_998),
.B(n_1108),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_SL g1132 ( 
.A1(n_1026),
.A2(n_1089),
.B1(n_1096),
.B2(n_1112),
.Y(n_1132)
);

OAI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1113),
.A2(n_1093),
.B1(n_995),
.B2(n_1087),
.Y(n_1133)
);

BUFx10_ASAP7_75t_L g1134 ( 
.A(n_1106),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1003),
.A2(n_1025),
.B1(n_1047),
.B2(n_1114),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1104),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1085),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1086),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1095),
.Y(n_1139)
);

BUFx2_ASAP7_75t_R g1140 ( 
.A(n_1050),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1039),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_994),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1109),
.Y(n_1143)
);

AO21x1_ASAP7_75t_SL g1144 ( 
.A1(n_1063),
.A2(n_1038),
.B(n_1055),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1091),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1047),
.A2(n_1110),
.B1(n_1111),
.B2(n_1041),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_1048),
.Y(n_1147)
);

CKINVDCx11_ASAP7_75t_R g1148 ( 
.A(n_1005),
.Y(n_1148)
);

INVx5_ASAP7_75t_L g1149 ( 
.A(n_1088),
.Y(n_1149)
);

NAND2x1p5_ASAP7_75t_L g1150 ( 
.A(n_1046),
.B(n_997),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1099),
.Y(n_1151)
);

OAI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1007),
.A2(n_1034),
.B1(n_1115),
.B2(n_1002),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_SL g1153 ( 
.A1(n_1018),
.A2(n_1107),
.B1(n_997),
.B2(n_1014),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1000),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1004),
.Y(n_1155)
);

INVx6_ASAP7_75t_L g1156 ( 
.A(n_1046),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1060),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1061),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1078),
.B(n_1101),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_SL g1160 ( 
.A1(n_1107),
.A2(n_1083),
.B1(n_1005),
.B2(n_1090),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1037),
.B(n_1036),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1031),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1008),
.A2(n_1024),
.B1(n_1040),
.B2(n_1044),
.Y(n_1163)
);

AOI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1076),
.A2(n_1064),
.B(n_1074),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1048),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1046),
.B(n_1098),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_SL g1167 ( 
.A1(n_1045),
.A2(n_1029),
.B1(n_1030),
.B2(n_1027),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1032),
.B(n_1037),
.Y(n_1168)
);

BUFx8_ASAP7_75t_L g1169 ( 
.A(n_1084),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1062),
.A2(n_1030),
.B1(n_1027),
.B2(n_1065),
.Y(n_1170)
);

INVx4_ASAP7_75t_L g1171 ( 
.A(n_1088),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_1051),
.B(n_1013),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1082),
.A2(n_1103),
.B1(n_1066),
.B2(n_1054),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_1000),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1054),
.A2(n_1052),
.B1(n_1053),
.B2(n_1010),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1048),
.B(n_1100),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1000),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1043),
.Y(n_1178)
);

AOI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1074),
.A2(n_1067),
.B(n_1068),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1056),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1043),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1043),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1100),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1100),
.B(n_1036),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_1056),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1072),
.A2(n_1088),
.B1(n_1051),
.B2(n_1067),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1057),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1057),
.A2(n_1071),
.B1(n_1069),
.B2(n_1077),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1069),
.A2(n_884),
.B1(n_765),
.B2(n_624),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1102),
.Y(n_1190)
);

BUFx8_ASAP7_75t_L g1191 ( 
.A(n_1020),
.Y(n_1191)
);

AO21x2_ASAP7_75t_L g1192 ( 
.A1(n_1070),
.A2(n_1058),
.B(n_1059),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1094),
.A2(n_765),
.B(n_432),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1049),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1094),
.A2(n_884),
.B1(n_765),
.B2(n_624),
.Y(n_1195)
);

BUFx12f_ASAP7_75t_L g1196 ( 
.A(n_1102),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_996),
.B(n_883),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1097),
.A2(n_861),
.B1(n_835),
.B2(n_847),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1075),
.A2(n_1073),
.B(n_1028),
.Y(n_1199)
);

INVx8_ASAP7_75t_L g1200 ( 
.A(n_994),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1097),
.A2(n_861),
.B1(n_978),
.B2(n_765),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1104),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1102),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_994),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1033),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1094),
.A2(n_978),
.B1(n_884),
.B2(n_784),
.Y(n_1206)
);

NAND2x1p5_ASAP7_75t_L g1207 ( 
.A(n_994),
.B(n_1109),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_1104),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1033),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1147),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1121),
.B(n_1194),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1121),
.B(n_1194),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1125),
.B(n_1144),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1165),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1125),
.B(n_1124),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1179),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1150),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1124),
.B(n_1180),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1164),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1185),
.B(n_1155),
.Y(n_1220)
);

AO21x2_ASAP7_75t_L g1221 ( 
.A1(n_1188),
.A2(n_1192),
.B(n_1130),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1185),
.B(n_1155),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1176),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1146),
.B(n_1129),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1172),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1193),
.A2(n_1195),
.B(n_1201),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1150),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1146),
.B(n_1129),
.Y(n_1228)
);

AO21x2_ASAP7_75t_L g1229 ( 
.A1(n_1188),
.A2(n_1192),
.B(n_1130),
.Y(n_1229)
);

INVx8_ASAP7_75t_L g1230 ( 
.A(n_1149),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1199),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1170),
.B(n_1151),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1170),
.B(n_1159),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1118),
.B(n_1135),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1120),
.B(n_1132),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1118),
.B(n_1135),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1186),
.A2(n_1187),
.B(n_1173),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1172),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1198),
.A2(n_1189),
.B(n_1206),
.Y(n_1239)
);

INVxp67_ASAP7_75t_R g1240 ( 
.A(n_1131),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1172),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1145),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1145),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1157),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1119),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1206),
.A2(n_1149),
.B(n_1198),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1123),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1197),
.B(n_1163),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1163),
.A2(n_1186),
.B(n_1137),
.Y(n_1249)
);

BUFx4f_ASAP7_75t_SL g1250 ( 
.A(n_1196),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1138),
.Y(n_1251)
);

INVxp33_ASAP7_75t_L g1252 ( 
.A(n_1202),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1139),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1141),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1205),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1209),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1171),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1119),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1158),
.Y(n_1259)
);

INVxp67_ASAP7_75t_SL g1260 ( 
.A(n_1152),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1153),
.B(n_1160),
.Y(n_1261)
);

OA21x2_ASAP7_75t_L g1262 ( 
.A1(n_1177),
.A2(n_1182),
.B(n_1178),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1152),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1223),
.B(n_1167),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1223),
.B(n_1181),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1235),
.A2(n_1133),
.B1(n_1175),
.B2(n_1140),
.Y(n_1266)
);

NOR2x1_ASAP7_75t_L g1267 ( 
.A(n_1219),
.B(n_1133),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1212),
.B(n_1168),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1210),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1211),
.B(n_1183),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1221),
.A2(n_1200),
.B(n_1207),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1210),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1232),
.B(n_1154),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1232),
.B(n_1154),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_1219),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1211),
.B(n_1136),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1221),
.B(n_1154),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1212),
.B(n_1142),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1241),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1239),
.A2(n_1161),
.B(n_1184),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1235),
.A2(n_1116),
.B1(n_1156),
.B2(n_1126),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1221),
.B(n_1154),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1221),
.B(n_1204),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1212),
.B(n_1204),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1229),
.B(n_1161),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1229),
.B(n_1166),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1229),
.B(n_1174),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1229),
.B(n_1143),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1214),
.B(n_1136),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1242),
.B(n_1208),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1251),
.B(n_1162),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1253),
.B(n_1162),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1216),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1253),
.B(n_1128),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1242),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1230),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1273),
.B(n_1234),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1272),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1266),
.A2(n_1226),
.B(n_1239),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1273),
.B(n_1234),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1268),
.B(n_1243),
.Y(n_1301)
);

AND2x2_ASAP7_75t_SL g1302 ( 
.A(n_1285),
.B(n_1241),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1266),
.A2(n_1226),
.B1(n_1263),
.B2(n_1248),
.Y(n_1303)
);

NAND3xp33_ASAP7_75t_L g1304 ( 
.A(n_1267),
.B(n_1263),
.C(n_1260),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1273),
.B(n_1236),
.Y(n_1305)
);

NAND3xp33_ASAP7_75t_L g1306 ( 
.A(n_1267),
.B(n_1260),
.C(n_1215),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1274),
.B(n_1236),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1274),
.B(n_1213),
.Y(n_1308)
);

NAND3xp33_ASAP7_75t_L g1309 ( 
.A(n_1281),
.B(n_1215),
.C(n_1248),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1281),
.A2(n_1246),
.B1(n_1233),
.B2(n_1261),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1274),
.B(n_1213),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1291),
.B(n_1244),
.Y(n_1312)
);

NOR3xp33_ASAP7_75t_L g1313 ( 
.A(n_1271),
.B(n_1233),
.C(n_1261),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1285),
.B(n_1218),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1290),
.B(n_1246),
.C(n_1245),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1292),
.B(n_1245),
.Y(n_1316)
);

NAND4xp25_ASAP7_75t_SL g1317 ( 
.A(n_1264),
.B(n_1224),
.C(n_1228),
.D(n_1218),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1285),
.B(n_1220),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1292),
.B(n_1294),
.Y(n_1319)
);

OAI221xp5_ASAP7_75t_L g1320 ( 
.A1(n_1290),
.A2(n_1238),
.B1(n_1225),
.B2(n_1258),
.C(n_1227),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1277),
.B(n_1220),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1277),
.B(n_1222),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1276),
.B(n_1252),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1276),
.B(n_1148),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1277),
.B(n_1222),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1282),
.B(n_1249),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1290),
.B(n_1259),
.C(n_1228),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1280),
.A2(n_1249),
.B1(n_1230),
.B2(n_1241),
.Y(n_1328)
);

NAND2xp33_ASAP7_75t_SL g1329 ( 
.A(n_1264),
.B(n_1241),
.Y(n_1329)
);

OAI221xp5_ASAP7_75t_L g1330 ( 
.A1(n_1271),
.A2(n_1238),
.B1(n_1225),
.B2(n_1227),
.C(n_1217),
.Y(n_1330)
);

NAND3xp33_ASAP7_75t_L g1331 ( 
.A(n_1289),
.B(n_1259),
.C(n_1249),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1289),
.B(n_1249),
.C(n_1264),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1283),
.A2(n_1237),
.B(n_1231),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1282),
.B(n_1262),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1280),
.B(n_1262),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1280),
.B(n_1262),
.Y(n_1336)
);

NAND3xp33_ASAP7_75t_L g1337 ( 
.A(n_1289),
.B(n_1255),
.C(n_1256),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1270),
.B(n_1254),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1270),
.B(n_1254),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1278),
.B(n_1247),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1334),
.B(n_1280),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1324),
.B(n_1148),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1326),
.B(n_1280),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1335),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1302),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1298),
.B(n_1295),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1336),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1337),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1340),
.B(n_1295),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1337),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1316),
.B(n_1278),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1339),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1329),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1302),
.B(n_1288),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1302),
.Y(n_1355)
);

AND2x4_ASAP7_75t_SL g1356 ( 
.A(n_1318),
.B(n_1296),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1333),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1314),
.B(n_1275),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1332),
.B(n_1279),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1333),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1314),
.B(n_1288),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1333),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1321),
.B(n_1287),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1323),
.B(n_1276),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1338),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1322),
.B(n_1286),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1332),
.B(n_1269),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1325),
.B(n_1286),
.Y(n_1368)
);

AND2x4_ASAP7_75t_SL g1369 ( 
.A(n_1313),
.B(n_1296),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1331),
.B(n_1279),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1299),
.A2(n_1240),
.B1(n_1238),
.B2(n_1284),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1319),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1301),
.B(n_1275),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1328),
.B(n_1293),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1352),
.B(n_1365),
.Y(n_1375)
);

NAND2xp67_ASAP7_75t_SL g1376 ( 
.A(n_1374),
.B(n_1265),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1345),
.B(n_1327),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1346),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1346),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1355),
.B(n_1354),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1352),
.B(n_1297),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1365),
.B(n_1364),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1373),
.B(n_1297),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1355),
.B(n_1308),
.Y(n_1384)
);

OR2x6_ASAP7_75t_L g1385 ( 
.A(n_1353),
.B(n_1304),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1354),
.B(n_1308),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1348),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1348),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1350),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1350),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1373),
.B(n_1300),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1349),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1349),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1351),
.B(n_1300),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1354),
.B(n_1311),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1358),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1358),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1361),
.B(n_1311),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1345),
.B(n_1327),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1361),
.B(n_1345),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1361),
.B(n_1366),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1342),
.B(n_1250),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1351),
.B(n_1305),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1369),
.A2(n_1306),
.B(n_1304),
.C(n_1309),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1372),
.B(n_1305),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1366),
.B(n_1307),
.Y(n_1406)
);

INVx3_ASAP7_75t_R g1407 ( 
.A(n_1353),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1359),
.B(n_1279),
.Y(n_1408)
);

INVxp33_ASAP7_75t_L g1409 ( 
.A(n_1371),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1367),
.B(n_1312),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1372),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1363),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1371),
.B(n_1306),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1343),
.B(n_1307),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1380),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1388),
.B(n_1367),
.Y(n_1416)
);

NAND2x1p5_ASAP7_75t_L g1417 ( 
.A(n_1413),
.B(n_1359),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1389),
.B(n_1343),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1401),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1390),
.B(n_1343),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1404),
.A2(n_1309),
.B1(n_1303),
.B2(n_1310),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1401),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1378),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1380),
.B(n_1341),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_1387),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1411),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1382),
.B(n_1341),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1392),
.B(n_1341),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1410),
.B(n_1367),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1385),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1379),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1385),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1385),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1400),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1410),
.B(n_1344),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1375),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1408),
.B(n_1400),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_L g1438 ( 
.A(n_1385),
.B(n_1315),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1393),
.B(n_1366),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1412),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_SL g1441 ( 
.A(n_1404),
.B(n_1413),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1381),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1396),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1397),
.B(n_1368),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1398),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1394),
.B(n_1368),
.Y(n_1446)
);

INVxp67_ASAP7_75t_L g1447 ( 
.A(n_1384),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1405),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1384),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1414),
.B(n_1344),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1408),
.B(n_1368),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1403),
.B(n_1344),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1407),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1406),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1406),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1383),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1398),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1453),
.B(n_1386),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1423),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1417),
.B(n_1386),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1415),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1441),
.Y(n_1462)
);

AO21x2_ASAP7_75t_L g1463 ( 
.A1(n_1430),
.A2(n_1362),
.B(n_1360),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1423),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1443),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1443),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1417),
.Y(n_1467)
);

INVxp67_ASAP7_75t_SL g1468 ( 
.A(n_1417),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1437),
.B(n_1395),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1431),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1426),
.B(n_1395),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1425),
.B(n_1409),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1440),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1421),
.B(n_1409),
.Y(n_1474)
);

CKINVDCx16_ASAP7_75t_R g1475 ( 
.A(n_1438),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1437),
.B(n_1377),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1415),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1416),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1451),
.B(n_1377),
.Y(n_1479)
);

CKINVDCx16_ASAP7_75t_R g1480 ( 
.A(n_1432),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1433),
.Y(n_1481)
);

INVx1_ASAP7_75t_SL g1482 ( 
.A(n_1429),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1419),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1419),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1447),
.B(n_1391),
.Y(n_1485)
);

CKINVDCx16_ASAP7_75t_R g1486 ( 
.A(n_1451),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1434),
.B(n_1377),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1416),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1429),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1445),
.B(n_1399),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1434),
.B(n_1399),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1442),
.B(n_1399),
.Y(n_1492)
);

INVxp67_ASAP7_75t_L g1493 ( 
.A(n_1436),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1475),
.A2(n_1462),
.B1(n_1474),
.B2(n_1486),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1468),
.A2(n_1436),
.B(n_1449),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1475),
.A2(n_1456),
.B1(n_1442),
.B2(n_1448),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1459),
.Y(n_1497)
);

OR3x1_ASAP7_75t_L g1498 ( 
.A(n_1477),
.B(n_1317),
.C(n_1402),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1486),
.A2(n_1480),
.B1(n_1472),
.B2(n_1467),
.Y(n_1499)
);

OAI221xp5_ASAP7_75t_L g1500 ( 
.A1(n_1481),
.A2(n_1448),
.B1(n_1456),
.B2(n_1422),
.C(n_1420),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1480),
.B(n_1454),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1459),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1458),
.B(n_1455),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1471),
.B(n_1445),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1467),
.B(n_1200),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1482),
.A2(n_1315),
.B(n_1359),
.Y(n_1506)
);

INVxp67_ASAP7_75t_SL g1507 ( 
.A(n_1467),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1458),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1464),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1464),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1465),
.Y(n_1511)
);

NOR4xp25_ASAP7_75t_L g1512 ( 
.A(n_1493),
.B(n_1418),
.C(n_1427),
.D(n_1428),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1465),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1460),
.A2(n_1369),
.B1(n_1359),
.B2(n_1370),
.Y(n_1514)
);

AOI211xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1461),
.A2(n_1330),
.B(n_1320),
.C(n_1424),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_L g1516 ( 
.A(n_1489),
.B(n_1117),
.C(n_1422),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1476),
.B(n_1457),
.Y(n_1517)
);

NOR2x1_ASAP7_75t_L g1518 ( 
.A(n_1466),
.B(n_1376),
.Y(n_1518)
);

INVx1_ASAP7_75t_SL g1519 ( 
.A(n_1476),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1508),
.B(n_1512),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1512),
.B(n_1519),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1503),
.B(n_1485),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1517),
.B(n_1469),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1516),
.A2(n_1460),
.B1(n_1485),
.B2(n_1479),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1497),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1502),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1501),
.B(n_1492),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1494),
.B(n_1477),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1509),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1499),
.B(n_1117),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1504),
.B(n_1478),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1496),
.B(n_1478),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1507),
.B(n_1469),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1495),
.B(n_1500),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1510),
.B(n_1470),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1505),
.B(n_1479),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1505),
.B(n_1490),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1511),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1505),
.Y(n_1539)
);

A2O1A1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1521),
.A2(n_1520),
.B(n_1534),
.C(n_1530),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_SL g1541 ( 
.A(n_1539),
.B(n_1506),
.Y(n_1541)
);

AOI221x1_ASAP7_75t_L g1542 ( 
.A1(n_1520),
.A2(n_1513),
.B1(n_1470),
.B2(n_1473),
.C(n_1466),
.Y(n_1542)
);

NAND4xp75_ASAP7_75t_L g1543 ( 
.A(n_1521),
.B(n_1518),
.C(n_1488),
.D(n_1514),
.Y(n_1543)
);

NOR4xp25_ASAP7_75t_L g1544 ( 
.A(n_1528),
.B(n_1488),
.C(n_1484),
.D(n_1483),
.Y(n_1544)
);

OAI211xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1532),
.A2(n_1527),
.B(n_1524),
.C(n_1533),
.Y(n_1545)
);

OAI21xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1523),
.A2(n_1490),
.B(n_1473),
.Y(n_1546)
);

AOI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1536),
.A2(n_1498),
.B1(n_1491),
.B2(n_1487),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1522),
.A2(n_1515),
.B1(n_1457),
.B2(n_1483),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1531),
.B(n_1537),
.Y(n_1549)
);

AOI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1525),
.A2(n_1484),
.B1(n_1487),
.B2(n_1491),
.C(n_1463),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1535),
.A2(n_1463),
.B(n_1487),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1548),
.A2(n_1539),
.B1(n_1491),
.B2(n_1487),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1540),
.A2(n_1535),
.B(n_1529),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1549),
.Y(n_1554)
);

OAI21xp33_ASAP7_75t_SL g1555 ( 
.A1(n_1543),
.A2(n_1538),
.B(n_1526),
.Y(n_1555)
);

NOR2x1p5_ASAP7_75t_SL g1556 ( 
.A(n_1544),
.B(n_1539),
.Y(n_1556)
);

NOR2xp67_ASAP7_75t_L g1557 ( 
.A(n_1546),
.B(n_1491),
.Y(n_1557)
);

NOR4xp25_ASAP7_75t_L g1558 ( 
.A(n_1545),
.B(n_1424),
.C(n_1435),
.D(n_1439),
.Y(n_1558)
);

NOR4xp25_ASAP7_75t_L g1559 ( 
.A(n_1550),
.B(n_1435),
.C(n_1444),
.D(n_1357),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1542),
.Y(n_1560)
);

O2A1O1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1560),
.A2(n_1541),
.B(n_1551),
.C(n_1463),
.Y(n_1561)
);

NOR4xp75_ASAP7_75t_L g1562 ( 
.A(n_1556),
.B(n_1547),
.C(n_1446),
.D(n_1191),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1553),
.A2(n_1203),
.B(n_1190),
.Y(n_1563)
);

NOR2x1_ASAP7_75t_L g1564 ( 
.A(n_1554),
.B(n_1127),
.Y(n_1564)
);

NAND4xp25_ASAP7_75t_L g1565 ( 
.A(n_1552),
.B(n_1359),
.C(n_1374),
.D(n_1452),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1564),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1563),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1561),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1565),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1562),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1565),
.A2(n_1555),
.B1(n_1557),
.B2(n_1558),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_SL g1572 ( 
.A(n_1571),
.B(n_1559),
.C(n_1191),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1569),
.Y(n_1573)
);

XOR2xp5_ASAP7_75t_L g1574 ( 
.A(n_1570),
.B(n_1122),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1566),
.B(n_1452),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1567),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1575),
.Y(n_1577)
);

NOR2x1_ASAP7_75t_L g1578 ( 
.A(n_1574),
.B(n_1568),
.Y(n_1578)
);

NAND4xp75_ASAP7_75t_L g1579 ( 
.A(n_1573),
.B(n_1567),
.C(n_1169),
.D(n_1134),
.Y(n_1579)
);

AO22x2_ASAP7_75t_L g1580 ( 
.A1(n_1579),
.A2(n_1576),
.B1(n_1572),
.B2(n_1169),
.Y(n_1580)
);

NAND3xp33_ASAP7_75t_L g1581 ( 
.A(n_1580),
.B(n_1578),
.C(n_1577),
.Y(n_1581)
);

OAI211xp5_ASAP7_75t_L g1582 ( 
.A1(n_1581),
.A2(n_1134),
.B(n_1362),
.C(n_1360),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1581),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1583),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1582),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1584),
.A2(n_1450),
.B(n_1357),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1585),
.A2(n_1450),
.B1(n_1369),
.B2(n_1347),
.Y(n_1587)
);

AOI21xp33_ASAP7_75t_L g1588 ( 
.A1(n_1586),
.A2(n_1357),
.B(n_1230),
.Y(n_1588)
);

XNOR2xp5_ASAP7_75t_L g1589 ( 
.A(n_1588),
.B(n_1587),
.Y(n_1589)
);

OAI221xp5_ASAP7_75t_R g1590 ( 
.A1(n_1589),
.A2(n_1230),
.B1(n_1347),
.B2(n_1370),
.C(n_1356),
.Y(n_1590)
);

AOI211xp5_ASAP7_75t_L g1591 ( 
.A1(n_1590),
.A2(n_1370),
.B(n_1374),
.C(n_1257),
.Y(n_1591)
);


endmodule