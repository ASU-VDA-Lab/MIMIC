module real_jpeg_19182_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_0),
.B(n_43),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_0),
.A2(n_42),
.B(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_0),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_0),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_0),
.A2(n_12),
.B(n_23),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_105),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_0),
.A2(n_81),
.B1(n_115),
.B2(n_116),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_0),
.B(n_69),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_1),
.A2(n_38),
.B1(n_43),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_52),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_52),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_38),
.B1(n_43),
.B2(n_76),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_25),
.Y(n_26)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_3),
.B(n_22),
.Y(n_132)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_5),
.A2(n_38),
.B1(n_43),
.B2(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_60),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_7),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_62),
.Y(n_101)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_11),
.A2(n_24),
.B1(n_34),
.B2(n_35),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_12),
.A2(n_34),
.B(n_56),
.C(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_34),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_12),
.A2(n_23),
.B1(n_25),
.B2(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_12),
.Y(n_58)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_92),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_91),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_63),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_18),
.B(n_63),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_45),
.C(n_53),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_19),
.A2(n_20),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_33),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_27),
.Y(n_21)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_25),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_26),
.B(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_26),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_26),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_30),
.A2(n_98),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_30),
.B(n_105),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.A3(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_49)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_40),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_35),
.A2(n_58),
.B(n_105),
.C(n_106),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_43),
.B(n_48),
.C(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_43),
.Y(n_48)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_45),
.A2(n_46),
.B1(n_53),
.B2(n_54),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_51),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_61),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_57),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_57),
.B(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_84),
.B2(n_85),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21x1_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_82),
.Y(n_78)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

XOR2x2_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_134),
.B(n_139),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_123),
.B(n_133),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_111),
.B(n_122),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_102),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_116),
.B(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_107),
.B2(n_108),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_107),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_117),
.B(n_121),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_125),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_130),
.C(n_131),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);


endmodule