module fake_jpeg_5349_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx6p67_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_34),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_0),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_15),
.B1(n_20),
.B2(n_16),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_25),
.B1(n_22),
.B2(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_27),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_26),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_15),
.B1(n_24),
.B2(n_19),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_16),
.B(n_27),
.C(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_38),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_19),
.B1(n_24),
.B2(n_20),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_55),
.B1(n_59),
.B2(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_60),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_25),
.B1(n_40),
.B2(n_17),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_49),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_22),
.B1(n_26),
.B2(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_21),
.B1(n_18),
.B2(n_4),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_39),
.B1(n_43),
.B2(n_21),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_71),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_21),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_66),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_51),
.C(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_89),
.Y(n_109)
);

AOI221xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_97),
.B1(n_81),
.B2(n_74),
.C(n_83),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_64),
.B(n_62),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_69),
.B(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_31),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_105),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_80),
.B1(n_74),
.B2(n_73),
.C(n_18),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_85),
.B1(n_90),
.B2(n_91),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_103),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_78),
.B(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_107),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_32),
.B(n_31),
.C(n_28),
.D(n_18),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_116),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_89),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_28),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_125),
.B1(n_113),
.B2(n_110),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_105),
.C(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_121),
.C(n_124),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_93),
.C(n_31),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_28),
.C(n_95),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_9),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_122),
.A2(n_111),
.B(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_128),
.B(n_7),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_116),
.B(n_123),
.C(n_4),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_130),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_134),
.B1(n_129),
.B2(n_8),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_6),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_136),
.A2(n_12),
.B(n_11),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_8),
.B(n_10),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_139),
.B(n_135),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_140),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_1),
.Y(n_142)
);


endmodule