module fake_netlist_1_9092_n_692 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_692);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_692;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g78 ( .A(n_67), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_16), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_19), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_57), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_22), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_30), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_16), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_70), .Y(n_85) );
BUFx2_ASAP7_75t_L g86 ( .A(n_9), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_52), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_65), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_19), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_53), .Y(n_90) );
HB1xp67_ASAP7_75t_L g91 ( .A(n_24), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_7), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_18), .Y(n_93) );
INVxp33_ASAP7_75t_SL g94 ( .A(n_51), .Y(n_94) );
INVxp67_ASAP7_75t_L g95 ( .A(n_50), .Y(n_95) );
CKINVDCx14_ASAP7_75t_R g96 ( .A(n_56), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_36), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_62), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_3), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_40), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_72), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_63), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_61), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_12), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_1), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_37), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_1), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_14), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_23), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_71), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_33), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_12), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_3), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_18), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_17), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_66), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_74), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_6), .Y(n_119) );
INVxp33_ASAP7_75t_L g120 ( .A(n_60), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_32), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_14), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_31), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_75), .Y(n_124) );
INVxp33_ASAP7_75t_SL g125 ( .A(n_42), .Y(n_125) );
AND2x2_ASAP7_75t_L g126 ( .A(n_86), .B(n_0), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_88), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_79), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_90), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_85), .B(n_0), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_80), .Y(n_143) );
INVx1_ASAP7_75t_SL g144 ( .A(n_87), .Y(n_144) );
OAI22xp33_ASAP7_75t_L g145 ( .A1(n_80), .A2(n_2), .B1(n_4), .B2(n_5), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_89), .B(n_84), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_107), .Y(n_147) );
AND2x6_ASAP7_75t_L g148 ( .A(n_98), .B(n_38), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_100), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_91), .B(n_2), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_109), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_100), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_101), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_101), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_108), .B(n_4), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_102), .Y(n_157) );
NAND2xp33_ASAP7_75t_L g158 ( .A(n_120), .B(n_77), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_84), .B(n_5), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_102), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_99), .B(n_6), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_103), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_108), .B(n_7), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_103), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_110), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_110), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_111), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_111), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_146), .B(n_116), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_152), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_159), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_152), .B(n_87), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_148), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_159), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_146), .B(n_116), .Y(n_175) );
AND2x4_ASAP7_75t_L g176 ( .A(n_146), .B(n_113), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_127), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_159), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_138), .B(n_119), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_138), .B(n_119), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
AND2x6_ASAP7_75t_L g185 ( .A(n_126), .B(n_112), .Y(n_185) );
OAI221xp5_ASAP7_75t_L g186 ( .A1(n_161), .A2(n_99), .B1(n_104), .B2(n_113), .C(n_122), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
AND2x6_ASAP7_75t_L g188 ( .A(n_126), .B(n_112), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_144), .B(n_96), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_144), .B(n_95), .Y(n_190) );
INVxp67_ASAP7_75t_SL g191 ( .A(n_141), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_149), .Y(n_192) );
OAI22xp33_ASAP7_75t_SL g193 ( .A1(n_141), .A2(n_105), .B1(n_106), .B2(n_93), .Y(n_193) );
INVxp33_ASAP7_75t_L g194 ( .A(n_156), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_128), .B(n_133), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_149), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_149), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_163), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_142), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_142), .Y(n_203) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_142), .Y(n_204) );
AO22x2_ASAP7_75t_L g205 ( .A1(n_163), .A2(n_121), .B1(n_124), .B2(n_123), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_128), .B(n_121), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_150), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_150), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_153), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_133), .B(n_122), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_135), .B(n_125), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_131), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_135), .B(n_124), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_153), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_136), .B(n_123), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_136), .B(n_104), .Y(n_218) );
BUFx10_ASAP7_75t_L g219 ( .A(n_148), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_137), .B(n_118), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_143), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_153), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_151), .A2(n_139), .B1(n_167), .B2(n_137), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_151), .Y(n_224) );
INVxp67_ASAP7_75t_L g225 ( .A(n_139), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_131), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_127), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_154), .B(n_118), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_154), .B(n_117), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_155), .Y(n_230) );
INVx4_ASAP7_75t_L g231 ( .A(n_148), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_196), .Y(n_232) );
INVx5_ASAP7_75t_L g233 ( .A(n_185), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_191), .B(n_162), .Y(n_234) );
INVxp67_ASAP7_75t_SL g235 ( .A(n_196), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_172), .B(n_160), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_207), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_218), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_169), .B(n_161), .Y(n_239) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_200), .Y(n_240) );
AND3x2_ASAP7_75t_SL g241 ( .A(n_221), .B(n_145), .C(n_92), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_173), .Y(n_242) );
BUFx3_ASAP7_75t_L g243 ( .A(n_173), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_171), .Y(n_244) );
OR2x6_ASAP7_75t_L g245 ( .A(n_205), .B(n_160), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_196), .Y(n_247) );
INVx3_ASAP7_75t_SL g248 ( .A(n_224), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_225), .B(n_167), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_170), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_207), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_207), .Y(n_252) );
INVx4_ASAP7_75t_L g253 ( .A(n_185), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_169), .B(n_164), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_212), .B(n_162), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_173), .Y(n_256) );
BUFx2_ASAP7_75t_SL g257 ( .A(n_185), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_218), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_169), .B(n_164), .Y(n_259) );
OR2x6_ASAP7_75t_L g260 ( .A(n_205), .B(n_195), .Y(n_260) );
INVxp67_ASAP7_75t_L g261 ( .A(n_182), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_231), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_184), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_224), .B(n_127), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_223), .B(n_168), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_175), .B(n_132), .Y(n_266) );
BUFx4f_ASAP7_75t_L g267 ( .A(n_185), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_175), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_219), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_231), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_185), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_220), .B(n_168), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_221), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_171), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_185), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_175), .B(n_132), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_188), .A2(n_158), .B1(n_148), .B2(n_94), .Y(n_277) );
INVx5_ASAP7_75t_L g278 ( .A(n_188), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_176), .Y(n_279) );
NAND2x1p5_ASAP7_75t_L g280 ( .A(n_231), .B(n_168), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_188), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_220), .B(n_166), .Y(n_282) );
OR2x2_ASAP7_75t_SL g283 ( .A(n_189), .B(n_114), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_219), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_207), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_219), .Y(n_286) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_174), .A2(n_117), .B(n_157), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_204), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_182), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_176), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_183), .Y(n_291) );
AOI22xp5_ASAP7_75t_SL g292 ( .A1(n_183), .A2(n_115), .B1(n_148), .B2(n_78), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_218), .Y(n_293) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_195), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_176), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_220), .B(n_166), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_188), .A2(n_148), .B1(n_166), .B2(n_157), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_211), .B(n_157), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_244), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_239), .B(n_188), .Y(n_300) );
AOI21x1_ASAP7_75t_L g301 ( .A1(n_265), .A2(n_181), .B(n_179), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_239), .B(n_188), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_233), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_244), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_236), .A2(n_171), .B(n_229), .C(n_228), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_253), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_253), .Y(n_307) );
AO32x2_ASAP7_75t_L g308 ( .A1(n_238), .A2(n_227), .A3(n_180), .B1(n_205), .B2(n_148), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_253), .B(n_211), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_244), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_233), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_239), .B(n_194), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_233), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_274), .Y(n_314) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_267), .B(n_205), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_274), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_235), .A2(n_194), .B1(n_186), .B2(n_190), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_232), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_297), .B(n_206), .C(n_214), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_247), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_298), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_245), .B(n_217), .Y(n_323) );
CKINVDCx5p33_ASAP7_75t_R g324 ( .A(n_248), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_240), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_254), .B(n_193), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_280), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_233), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_245), .B(n_155), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_250), .B(n_180), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_233), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_238), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_278), .B(n_155), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_298), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_261), .B(n_227), .Y(n_335) );
AND2x2_ASAP7_75t_SL g336 ( .A(n_267), .B(n_230), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_234), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_245), .A2(n_148), .B1(n_222), .B2(n_197), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_278), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_254), .B(n_210), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_280), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_242), .Y(n_342) );
BUFx12f_ASAP7_75t_L g343 ( .A(n_273), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_248), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_245), .A2(n_192), .B1(n_202), .B2(n_215), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_294), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_260), .B(n_289), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_260), .A2(n_208), .B1(n_198), .B2(n_209), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_260), .A2(n_134), .B1(n_147), .B2(n_140), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_260), .A2(n_165), .B1(n_147), .B2(n_140), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_337), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_329), .A2(n_267), .B1(n_293), .B2(n_258), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_337), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_315), .B(n_254), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_324), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_319), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_315), .A2(n_294), .B1(n_292), .B2(n_273), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_325), .B(n_278), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_310), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_344), .Y(n_360) );
AO222x2_ASAP7_75t_L g361 ( .A1(n_346), .A2(n_241), .B1(n_283), .B2(n_276), .C1(n_266), .C2(n_291), .Y(n_361) );
CKINVDCx12_ASAP7_75t_R g362 ( .A(n_329), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_312), .B(n_259), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_322), .B(n_259), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_329), .A2(n_296), .B1(n_272), .B2(n_282), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_329), .B(n_309), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_309), .B(n_278), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_348), .A2(n_257), .B1(n_293), .B2(n_258), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_326), .B(n_283), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_310), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
AOI21x1_ASAP7_75t_L g372 ( .A1(n_301), .A2(n_226), .B(n_213), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_314), .Y(n_373) );
NAND3xp33_ASAP7_75t_L g374 ( .A(n_305), .B(n_277), .C(n_131), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_306), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_309), .B(n_259), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_322), .B(n_278), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_323), .A2(n_271), .B1(n_275), .B2(n_281), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_347), .A2(n_271), .B1(n_275), .B2(n_268), .Y(n_379) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_336), .B(n_266), .Y(n_380) );
CKINVDCx6p67_ASAP7_75t_R g381 ( .A(n_343), .Y(n_381) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_318), .A2(n_255), .B(n_241), .C(n_264), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_347), .A2(n_295), .B1(n_290), .B2(n_279), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_359), .Y(n_384) );
INVx4_ASAP7_75t_L g385 ( .A(n_366), .Y(n_385) );
AOI332xp33_ASAP7_75t_L g386 ( .A1(n_361), .A2(n_129), .A3(n_130), .B1(n_132), .B2(n_334), .B3(n_134), .C1(n_147), .C2(n_140), .Y(n_386) );
OAI211xp5_ASAP7_75t_L g387 ( .A1(n_382), .A2(n_334), .B(n_335), .C(n_330), .Y(n_387) );
INVx1_ASAP7_75t_SL g388 ( .A(n_360), .Y(n_388) );
AOI222xp33_ASAP7_75t_L g389 ( .A1(n_369), .A2(n_343), .B1(n_321), .B2(n_323), .C1(n_263), .C2(n_276), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_357), .A2(n_300), .B1(n_302), .B2(n_276), .Y(n_391) );
OAI211xp5_ASAP7_75t_SL g392 ( .A1(n_382), .A2(n_350), .B(n_129), .C(n_130), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_351), .B(n_327), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_351), .A2(n_130), .B1(n_129), .B2(n_132), .C(n_321), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_380), .A2(n_324), .B1(n_345), .B2(n_349), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_353), .A2(n_130), .B1(n_129), .B2(n_266), .C(n_249), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_375), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_380), .A2(n_320), .B1(n_336), .B2(n_333), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_380), .A2(n_333), .B1(n_281), .B2(n_341), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_364), .B(n_327), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_356), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_359), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_356), .B(n_287), .Y(n_404) );
OAI211xp5_ASAP7_75t_L g405 ( .A1(n_383), .A2(n_340), .B(n_338), .C(n_341), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_363), .A2(n_134), .B1(n_332), .B2(n_304), .C(n_299), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
BUFx8_ASAP7_75t_SL g408 ( .A(n_355), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_365), .A2(n_304), .B1(n_299), .B2(n_316), .C(n_301), .Y(n_409) );
OA21x2_ASAP7_75t_L g410 ( .A1(n_372), .A2(n_226), .B(n_213), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_364), .B(n_308), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_384), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_402), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_393), .B(n_371), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_388), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_389), .A2(n_365), .B1(n_362), .B2(n_366), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_389), .A2(n_362), .B1(n_366), .B2(n_354), .Y(n_417) );
OAI31xp33_ASAP7_75t_L g418 ( .A1(n_392), .A2(n_368), .A3(n_354), .B(n_366), .Y(n_418) );
OA21x2_ASAP7_75t_L g419 ( .A1(n_409), .A2(n_372), .B(n_374), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_387), .A2(n_371), .B1(n_374), .B2(n_376), .C(n_368), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_393), .B(n_370), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_402), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_387), .A2(n_352), .B1(n_378), .B2(n_379), .Y(n_423) );
OAI31xp33_ASAP7_75t_SL g424 ( .A1(n_392), .A2(n_378), .A3(n_367), .B(n_377), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_384), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_393), .B(n_370), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_401), .B(n_373), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_395), .B(n_165), .C(n_131), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_395), .A2(n_373), .B1(n_381), .B2(n_281), .Y(n_429) );
OAI211xp5_ASAP7_75t_SL g430 ( .A1(n_388), .A2(n_97), .B(n_358), .C(n_381), .Y(n_430) );
NAND5xp2_ASAP7_75t_L g431 ( .A(n_386), .B(n_280), .C(n_316), .D(n_308), .E(n_281), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_396), .B(n_287), .Y(n_432) );
OAI33xp33_ASAP7_75t_L g433 ( .A1(n_396), .A2(n_187), .A3(n_177), .B1(n_178), .B2(n_201), .B3(n_203), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_391), .A2(n_377), .B1(n_367), .B2(n_287), .Y(n_434) );
AOI21xp33_ASAP7_75t_SL g435 ( .A1(n_386), .A2(n_8), .B(n_9), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_401), .B(n_373), .Y(n_436) );
BUFx3_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_397), .A2(n_377), .B1(n_367), .B2(n_333), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_397), .A2(n_377), .B1(n_367), .B2(n_317), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_385), .A2(n_314), .B1(n_317), .B2(n_281), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_398), .Y(n_441) );
AOI211xp5_ASAP7_75t_SL g442 ( .A1(n_409), .A2(n_375), .B(n_339), .C(n_311), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_406), .A2(n_375), .B1(n_306), .B2(n_307), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_390), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_390), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_399), .A2(n_165), .B1(n_375), .B2(n_331), .C(n_313), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_416), .A2(n_400), .B(n_394), .Y(n_447) );
AND2x2_ASAP7_75t_SL g448 ( .A(n_416), .B(n_385), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_414), .B(n_401), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_444), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_414), .B(n_385), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_435), .B(n_415), .C(n_428), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_435), .B(n_431), .Y(n_453) );
OAI33xp33_ASAP7_75t_L g454 ( .A1(n_413), .A2(n_404), .A3(n_10), .B1(n_11), .B2(n_13), .B3(n_15), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_444), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
CKINVDCx6p67_ASAP7_75t_R g457 ( .A(n_426), .Y(n_457) );
AOI33xp33_ASAP7_75t_L g458 ( .A1(n_422), .A2(n_411), .A3(n_394), .B1(n_13), .B2(n_15), .B3(n_17), .Y(n_458) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_428), .B(n_131), .C(n_404), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_445), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_430), .B(n_131), .C(n_411), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_427), .B(n_385), .Y(n_462) );
OAI221xp5_ASAP7_75t_SL g463 ( .A1(n_417), .A2(n_406), .B1(n_405), .B2(n_411), .C(n_407), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_422), .Y(n_464) );
OAI321xp33_ASAP7_75t_L g465 ( .A1(n_429), .A2(n_405), .A3(n_398), .B1(n_407), .B2(n_403), .C(n_390), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_421), .Y(n_466) );
INVx5_ASAP7_75t_L g467 ( .A(n_441), .Y(n_467) );
NAND2xp33_ASAP7_75t_R g468 ( .A(n_419), .B(n_410), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_437), .B(n_403), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_426), .B(n_403), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_420), .B(n_398), .C(n_204), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
OAI31xp33_ASAP7_75t_SL g473 ( .A1(n_443), .A2(n_407), .A3(n_408), .B(n_308), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_427), .Y(n_474) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_432), .A2(n_410), .B(n_187), .Y(n_475) );
AOI33xp33_ASAP7_75t_L g476 ( .A1(n_417), .A2(n_434), .A3(n_439), .B1(n_438), .B2(n_423), .B3(n_436), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_436), .B(n_398), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_445), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_412), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_412), .B(n_398), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_425), .B(n_398), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_437), .B(n_8), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_437), .B(n_398), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_425), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_418), .B(n_10), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_441), .Y(n_486) );
OAI33xp33_ASAP7_75t_L g487 ( .A1(n_418), .A2(n_177), .A3(n_178), .B1(n_201), .B2(n_203), .B3(n_308), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_423), .B(n_410), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_446), .A2(n_410), .B1(n_331), .B2(n_313), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_440), .B(n_20), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_424), .B(n_410), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_433), .B(n_199), .C(n_339), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_419), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_419), .Y(n_494) );
OAI21xp33_ASAP7_75t_SL g495 ( .A1(n_442), .A2(n_328), .B(n_308), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_419), .B(n_342), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_453), .A2(n_342), .B1(n_339), .B2(n_311), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_450), .B(n_204), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_450), .B(n_204), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_455), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_457), .B(n_21), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_473), .B(n_306), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_455), .B(n_204), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_456), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_464), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_453), .B(n_25), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_466), .B(n_26), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_460), .B(n_27), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_478), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_460), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_482), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_474), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_486), .B(n_216), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_449), .B(n_216), .Y(n_514) );
BUFx2_ASAP7_75t_L g515 ( .A(n_469), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_472), .B(n_28), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_448), .A2(n_342), .B1(n_311), .B2(n_303), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_488), .B(n_29), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_470), .B(n_216), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_479), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_469), .B(n_34), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_451), .B(n_216), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_494), .B(n_35), .Y(n_523) );
NOR3xp33_ASAP7_75t_SL g524 ( .A(n_454), .B(n_39), .C(n_41), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_490), .B(n_328), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_467), .B(n_43), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_484), .Y(n_527) );
AND2x4_ASAP7_75t_L g528 ( .A(n_467), .B(n_44), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_480), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_477), .B(n_216), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_462), .B(n_45), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_452), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_481), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_476), .B(n_46), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_458), .Y(n_535) );
NOR3xp33_ASAP7_75t_L g536 ( .A(n_461), .B(n_199), .C(n_328), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_475), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_491), .B(n_199), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_496), .B(n_47), .Y(n_539) );
INVx4_ASAP7_75t_L g540 ( .A(n_467), .Y(n_540) );
OAI222xp33_ASAP7_75t_L g541 ( .A1(n_463), .A2(n_303), .B1(n_49), .B2(n_54), .C1(n_55), .C2(n_58), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_475), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_496), .B(n_48), .Y(n_543) );
OAI33xp33_ASAP7_75t_L g544 ( .A1(n_489), .A2(n_59), .A3(n_64), .B1(n_68), .B2(n_69), .B3(n_73), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_458), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_485), .B(n_76), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_475), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_447), .B(n_342), .C(n_307), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_476), .B(n_342), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_448), .B(n_493), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_483), .B(n_307), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_467), .B(n_307), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_490), .A2(n_495), .B1(n_487), .B2(n_471), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_483), .B(n_307), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_529), .B(n_490), .Y(n_555) );
NOR2x1p5_ASAP7_75t_SL g556 ( .A(n_537), .B(n_468), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_510), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_529), .B(n_459), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_504), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_500), .B(n_468), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_500), .B(n_492), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_505), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_550), .B(n_492), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_509), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_512), .B(n_465), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_550), .B(n_237), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_532), .B(n_306), .Y(n_567) );
NAND4xp75_ASAP7_75t_L g568 ( .A(n_535), .B(n_306), .C(n_237), .D(n_285), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_511), .B(n_285), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_545), .B(n_252), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_520), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_533), .B(n_252), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_527), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_515), .B(n_251), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_538), .B(n_251), .Y(n_575) );
AO21x1_ASAP7_75t_L g576 ( .A1(n_502), .A2(n_246), .B(n_288), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_540), .Y(n_577) );
NOR2xp33_ASAP7_75t_R g578 ( .A(n_501), .B(n_242), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_513), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_506), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_513), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_519), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_518), .B(n_246), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_519), .Y(n_584) );
AND3x1_ASAP7_75t_L g585 ( .A(n_524), .B(n_288), .C(n_256), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_531), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_542), .B(n_288), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_547), .B(n_243), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_547), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g590 ( .A1(n_553), .A2(n_243), .B(n_256), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_530), .B(n_262), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_531), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_514), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_523), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_518), .B(n_262), .Y(n_595) );
NOR2x1_ASAP7_75t_L g596 ( .A(n_540), .B(n_270), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_549), .B(n_270), .Y(n_597) );
INVx4_ASAP7_75t_L g598 ( .A(n_540), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_522), .B(n_269), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_539), .B(n_269), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_539), .B(n_269), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_523), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_525), .B(n_269), .Y(n_603) );
XOR2x2_ASAP7_75t_L g604 ( .A(n_585), .B(n_525), .Y(n_604) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_598), .B(n_548), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_586), .B(n_543), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_584), .B(n_543), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_580), .B(n_534), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_559), .Y(n_609) );
NAND2xp33_ASAP7_75t_SL g610 ( .A(n_598), .B(n_502), .Y(n_610) );
AOI322xp5_ASAP7_75t_L g611 ( .A1(n_592), .A2(n_546), .A3(n_517), .B1(n_516), .B2(n_521), .C1(n_497), .C2(n_528), .Y(n_611) );
AOI211xp5_ASAP7_75t_SL g612 ( .A1(n_590), .A2(n_541), .B(n_528), .C(n_526), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_581), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_562), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_560), .Y(n_615) );
OA22x2_ASAP7_75t_L g616 ( .A1(n_598), .A2(n_577), .B1(n_563), .B2(n_564), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_565), .A2(n_544), .B(n_507), .C(n_536), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_571), .B(n_521), .Y(n_618) );
AO211x2_ASAP7_75t_L g619 ( .A1(n_573), .A2(n_526), .B(n_528), .C(n_508), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_573), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_577), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_557), .B(n_554), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_596), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_579), .B(n_554), .Y(n_624) );
XOR2xp5_ASAP7_75t_L g625 ( .A(n_563), .B(n_526), .Y(n_625) );
BUFx2_ASAP7_75t_L g626 ( .A(n_560), .Y(n_626) );
XOR2x2_ASAP7_75t_L g627 ( .A(n_568), .B(n_508), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_582), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_558), .Y(n_629) );
XOR2x2_ASAP7_75t_L g630 ( .A(n_568), .B(n_552), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_593), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_561), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_561), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_558), .B(n_498), .Y(n_634) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_603), .B(n_552), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_567), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_603), .Y(n_637) );
AOI321xp33_ASAP7_75t_L g638 ( .A1(n_555), .A2(n_499), .A3(n_503), .B1(n_552), .B2(n_551), .C(n_286), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_578), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_570), .B(n_499), .C(n_503), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_569), .B(n_284), .C(n_286), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_594), .A2(n_284), .B1(n_602), .B2(n_575), .C(n_589), .Y(n_642) );
INVx1_ASAP7_75t_SL g643 ( .A(n_566), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_602), .B(n_566), .Y(n_644) );
OAI211xp5_ASAP7_75t_SL g645 ( .A1(n_574), .A2(n_583), .B(n_597), .C(n_601), .Y(n_645) );
NAND4xp25_ASAP7_75t_L g646 ( .A(n_595), .B(n_591), .C(n_572), .D(n_600), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_600), .B(n_572), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_591), .A2(n_595), .B1(n_599), .B2(n_588), .Y(n_648) );
XNOR2x1_ASAP7_75t_L g649 ( .A(n_556), .B(n_599), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_576), .A2(n_532), .B1(n_580), .B2(n_145), .C(n_545), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_556), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g652 ( .A1(n_587), .A2(n_453), .A3(n_535), .B1(n_545), .B2(n_580), .C1(n_532), .C2(n_586), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_587), .B(n_588), .C(n_576), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_559), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_559), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_633), .Y(n_656) );
XNOR2x2_ASAP7_75t_L g657 ( .A(n_616), .B(n_639), .Y(n_657) );
INVx3_ASAP7_75t_L g658 ( .A(n_616), .Y(n_658) );
XNOR2x1_ASAP7_75t_L g659 ( .A(n_649), .B(n_619), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_649), .A2(n_608), .B1(n_629), .B2(n_632), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_620), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_650), .A2(n_629), .B1(n_631), .B2(n_626), .C(n_609), .Y(n_662) );
AOI32xp33_ASAP7_75t_L g663 ( .A1(n_612), .A2(n_610), .A3(n_605), .B1(n_637), .B2(n_651), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_655), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_654), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_612), .A2(n_652), .B(n_625), .Y(n_666) );
NAND4xp75_ASAP7_75t_L g667 ( .A(n_623), .B(n_635), .C(n_606), .D(n_642), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_617), .B(n_645), .C(n_641), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g669 ( .A1(n_611), .A2(n_646), .B(n_653), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_666), .A2(n_604), .B(n_621), .Y(n_670) );
AOI211xp5_ASAP7_75t_SL g671 ( .A1(n_669), .A2(n_648), .B(n_653), .C(n_636), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_656), .B(n_658), .Y(n_672) );
AO22x2_ASAP7_75t_L g673 ( .A1(n_658), .A2(n_614), .B1(n_637), .B2(n_613), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_660), .B(n_659), .Y(n_674) );
NAND4xp25_ASAP7_75t_SL g675 ( .A(n_663), .B(n_643), .C(n_607), .D(n_640), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_662), .A2(n_630), .B(n_627), .Y(n_676) );
OAI211xp5_ASAP7_75t_SL g677 ( .A1(n_668), .A2(n_638), .B(n_628), .C(n_634), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_670), .B(n_664), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_674), .B(n_657), .Y(n_679) );
NAND4xp25_ASAP7_75t_SL g680 ( .A(n_676), .B(n_667), .C(n_615), .D(n_634), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_671), .A2(n_665), .B1(n_661), .B2(n_618), .C(n_640), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_673), .A2(n_624), .B1(n_644), .B2(n_622), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_678), .B(n_672), .Y(n_683) );
AOI322xp5_ASAP7_75t_L g684 ( .A1(n_679), .A2(n_675), .A3(n_677), .B1(n_673), .B2(n_624), .C1(n_622), .C2(n_647), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_682), .Y(n_685) );
INVx3_ASAP7_75t_L g686 ( .A(n_683), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_685), .Y(n_687) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_687), .Y(n_688) );
AO21x2_ASAP7_75t_L g689 ( .A1(n_687), .A2(n_681), .B(n_686), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_688), .A2(n_686), .B(n_680), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_690), .A2(n_686), .B1(n_689), .B2(n_684), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_691), .A2(n_686), .B(n_689), .Y(n_692) );
endmodule