module fake_jpeg_28672_n_525 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_434;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_55),
.Y(n_144)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_56),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_62),
.Y(n_108)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_75),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_34),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_77),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_34),
.B(n_14),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_85),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx4f_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx5_ASAP7_75t_SL g132 ( 
.A(n_82),
.Y(n_132)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_86),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_20),
.B(n_15),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_89),
.B(n_93),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_20),
.B(n_15),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_27),
.Y(n_118)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_21),
.B(n_15),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_26),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_118),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_27),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_119),
.B(n_142),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_82),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_125),
.B(n_131),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_21),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_128),
.B(n_133),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_82),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_46),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_62),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_134),
.A2(n_157),
.B(n_50),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_90),
.A2(n_39),
.B1(n_50),
.B2(n_29),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_95),
.B1(n_39),
.B2(n_96),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_81),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_57),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_143),
.B(n_161),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_74),
.B(n_41),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_155),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_41),
.Y(n_155)
);

INVx2_ASAP7_75t_R g157 ( 
.A(n_67),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_22),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_166),
.A2(n_182),
.B1(n_185),
.B2(n_194),
.Y(n_224)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_170),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_129),
.B(n_149),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_134),
.C(n_48),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_39),
.B1(n_60),
.B2(n_38),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_186),
.B1(n_193),
.B2(n_215),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_204),
.Y(n_223)
);

CKINVDCx6p67_ASAP7_75t_R g179 ( 
.A(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_179),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_105),
.A2(n_87),
.B1(n_84),
.B2(n_80),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_181),
.A2(n_208),
.B1(n_152),
.B2(n_121),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_68),
.B1(n_92),
.B2(n_73),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_183),
.Y(n_256)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_71),
.B1(n_66),
.B2(n_59),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_120),
.A2(n_28),
.B1(n_40),
.B2(n_38),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_191),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_111),
.A2(n_44),
.B1(n_40),
.B2(n_48),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_140),
.A2(n_58),
.B1(n_24),
.B2(n_47),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_107),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_196),
.B(n_209),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_198),
.Y(n_253)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_200),
.Y(n_260)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_202),
.Y(n_254)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_137),
.A2(n_116),
.B(n_160),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_168),
.Y(n_228)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_141),
.A2(n_24),
.B1(n_47),
.B2(n_50),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_210),
.Y(n_255)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_212),
.B(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_99),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_218),
.Y(n_239)
);

CKINVDCx12_ASAP7_75t_R g214 ( 
.A(n_108),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_124),
.B1(n_127),
.B2(n_147),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_137),
.A2(n_47),
.B1(n_22),
.B2(n_43),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g216 ( 
.A(n_135),
.B(n_67),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_217),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_119),
.B(n_43),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_105),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_228),
.B(n_173),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_235),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_164),
.B(n_127),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_258),
.B(n_217),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_168),
.B(n_130),
.C(n_164),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_246),
.C(n_259),
.Y(n_283)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_245),
.A2(n_151),
.B1(n_219),
.B2(n_210),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_167),
.B(n_108),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_152),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_200),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_176),
.B(n_121),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_232),
.CI(n_240),
.CON(n_276),
.SN(n_276)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_172),
.A2(n_23),
.B(n_46),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_195),
.B(n_44),
.Y(n_259)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_216),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_262),
.A2(n_265),
.B(n_269),
.Y(n_304)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_264),
.B(n_282),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_224),
.A2(n_123),
.B1(n_151),
.B2(n_185),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_267),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_173),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_231),
.A2(n_183),
.B1(n_170),
.B2(n_204),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_268),
.A2(n_231),
.B1(n_226),
.B2(n_229),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_232),
.A2(n_197),
.B(n_207),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_169),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_270),
.B(n_271),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_192),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_222),
.A2(n_224),
.B1(n_234),
.B2(n_245),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_272),
.A2(n_274),
.B1(n_290),
.B2(n_180),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_288),
.B1(n_249),
.B2(n_261),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_247),
.A2(n_211),
.B1(n_136),
.B2(n_162),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_275),
.B(n_276),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_228),
.B(n_23),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_278),
.B(n_279),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_199),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_237),
.A2(n_189),
.B1(n_177),
.B2(n_136),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_280),
.B(n_284),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_179),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_293),
.C(n_227),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_252),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_188),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_236),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_286),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_250),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_287),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_258),
.A2(n_162),
.B1(n_190),
.B2(n_171),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_249),
.A2(n_203),
.B1(n_179),
.B2(n_175),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_220),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_291),
.B(n_295),
.Y(n_314)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_223),
.B(n_179),
.C(n_52),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_26),
.B(n_37),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_235),
.B(n_251),
.C(n_254),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_236),
.Y(n_294)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_52),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_302),
.A2(n_325),
.B1(n_331),
.B2(n_294),
.Y(n_358)
);

OAI32xp33_ASAP7_75t_L g307 ( 
.A1(n_270),
.A2(n_255),
.A3(n_221),
.B1(n_242),
.B2(n_227),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_329),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_309),
.A2(n_292),
.B1(n_282),
.B2(n_291),
.Y(n_344)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_311),
.Y(n_332)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_225),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_319),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_287),
.B(n_256),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_323),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_318),
.A2(n_286),
.B1(n_296),
.B2(n_277),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_265),
.A2(n_229),
.B(n_257),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_320),
.A2(n_269),
.B(n_289),
.Y(n_348)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_263),
.Y(n_322)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_322),
.Y(n_362)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_260),
.C(n_238),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_283),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_273),
.A2(n_238),
.B1(n_226),
.B2(n_241),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_288),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_295),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_266),
.A2(n_244),
.B1(n_233),
.B2(n_114),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_279),
.Y(n_335)
);

NOR4xp25_ASAP7_75t_L g366 ( 
.A(n_335),
.B(n_351),
.C(n_354),
.D(n_333),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_330),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_357),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_337),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_276),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_361),
.Y(n_388)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_262),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_343),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_317),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_341),
.B(n_348),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_313),
.Y(n_342)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_342),
.Y(n_369)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_262),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_344),
.A2(n_358),
.B1(n_359),
.B2(n_306),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_319),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_345),
.B(n_352),
.C(n_324),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_284),
.Y(n_346)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_303),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_267),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_278),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_328),
.A2(n_276),
.B1(n_293),
.B2(n_277),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_356),
.A2(n_360),
.B1(n_302),
.B2(n_309),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_312),
.A2(n_277),
.B1(n_294),
.B2(n_286),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_298),
.B(n_276),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_301),
.B(n_264),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_301),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_364),
.A2(n_358),
.B1(n_307),
.B2(n_310),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_363),
.B(n_314),
.Y(n_371)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_355),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_372),
.B(n_380),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_314),
.Y(n_375)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_375),
.Y(n_402)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_342),
.Y(n_376)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_332),
.Y(n_377)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_395),
.C(n_350),
.Y(n_397)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_379),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_362),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_347),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_382),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_339),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_383),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_384),
.B(n_322),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_346),
.B(n_299),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_386),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_326),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_344),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_338),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_389),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_338),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_390),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_311),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_391),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_361),
.B(n_310),
.Y(n_392)
);

AOI21xp33_ASAP7_75t_L g419 ( 
.A1(n_392),
.A2(n_393),
.B(n_305),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_348),
.B(n_308),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_298),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_394),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_320),
.C(n_321),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_397),
.B(n_399),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_373),
.A2(n_334),
.B(n_336),
.Y(n_399)
);

BUFx12f_ASAP7_75t_SL g405 ( 
.A(n_393),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_405),
.A2(n_411),
.B(n_388),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_350),
.C(n_395),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_408),
.B(n_409),
.C(n_388),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_387),
.B(n_356),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_364),
.A2(n_331),
.B1(n_325),
.B2(n_334),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_410),
.A2(n_416),
.B1(n_421),
.B2(n_380),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_367),
.A2(n_343),
.B(n_340),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_417),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_374),
.Y(n_415)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_415),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_419),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_368),
.A2(n_305),
.B1(n_303),
.B2(n_327),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_388),
.B(n_124),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_385),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_405),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_427),
.Y(n_450)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_384),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_407),
.Y(n_428)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_428),
.Y(n_459)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_420),
.Y(n_430)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_430),
.Y(n_465)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_420),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_435),
.Y(n_455)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_406),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_432),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_402),
.B(n_365),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_433),
.B(n_442),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_396),
.A2(n_368),
.B1(n_376),
.B2(n_369),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_434),
.A2(n_441),
.B1(n_444),
.B2(n_416),
.Y(n_447)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

AO21x1_ASAP7_75t_L g458 ( 
.A1(n_438),
.A2(n_423),
.B(n_414),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_411),
.A2(n_373),
.B(n_394),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_439),
.A2(n_403),
.B(n_410),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_445),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_404),
.A2(n_390),
.B1(n_389),
.B2(n_369),
.Y(n_441)
);

BUFx24_ASAP7_75t_SL g442 ( 
.A(n_403),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_414),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_443),
.A2(n_377),
.B1(n_382),
.B2(n_374),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_370),
.B1(n_386),
.B2(n_379),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_445),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_447),
.B(n_462),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_437),
.B(n_397),
.C(n_408),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_457),
.C(n_461),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_441),
.A2(n_423),
.B(n_399),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_452),
.A2(n_454),
.B(n_458),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_409),
.C(n_417),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_444),
.A2(n_370),
.B1(n_413),
.B2(n_400),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_460),
.A2(n_463),
.B1(n_425),
.B2(n_432),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_440),
.B(n_412),
.C(n_422),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_436),
.A2(n_381),
.B1(n_244),
.B2(n_233),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_464),
.B(n_438),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_467),
.B(n_461),
.Y(n_487)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_468),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_449),
.A2(n_428),
.B1(n_426),
.B2(n_434),
.Y(n_469)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_469),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_439),
.Y(n_470)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_458),
.A2(n_429),
.B(n_148),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_471),
.A2(n_478),
.B(n_3),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_456),
.B(n_429),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_475),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_178),
.C(n_124),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_476),
.C(n_477),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_178),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_37),
.C(n_50),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_50),
.C(n_42),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_454),
.A2(n_0),
.B(n_1),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_447),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_482),
.C(n_3),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_452),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_481),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_455),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_467),
.A2(n_465),
.B1(n_451),
.B2(n_463),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_487),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_451),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_485),
.A2(n_488),
.B(n_482),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_459),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_8),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_491),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_480),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_492),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_473),
.B(n_6),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_8),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_502),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_499),
.A2(n_501),
.B(n_487),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_473),
.C(n_479),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_500),
.B(n_505),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_496),
.A2(n_474),
.B(n_476),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_484),
.A2(n_477),
.B(n_10),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_503),
.B(n_506),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_42),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_493),
.A2(n_11),
.B(n_13),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_507),
.B(n_491),
.Y(n_508)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_508),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_509),
.B(n_513),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_495),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_500),
.A2(n_486),
.B1(n_13),
.B2(n_42),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_497),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_SL g519 ( 
.A1(n_515),
.A2(n_512),
.B(n_510),
.C(n_508),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_511),
.A2(n_504),
.B(n_486),
.Y(n_516)
);

AOI31xp33_ASAP7_75t_L g520 ( 
.A1(n_516),
.A2(n_506),
.A3(n_498),
.B(n_13),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_519),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_518),
.B1(n_517),
.B2(n_520),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_522),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_42),
.C(n_26),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_42),
.Y(n_525)
);


endmodule