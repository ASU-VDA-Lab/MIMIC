module fake_jpeg_28625_n_486 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_486);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_486;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_60),
.Y(n_148)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_61),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_16),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_63),
.B(n_72),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_74),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_15),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_1),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_20),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_1),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_77),
.B(n_93),
.Y(n_140)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_34),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_44),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_45),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_27),
.B(n_3),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_97),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_17),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

BUFx6f_ASAP7_75t_SL g147 ( 
.A(n_99),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_34),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_105),
.B(n_137),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_55),
.A2(n_32),
.B1(n_42),
.B2(n_31),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_110),
.A2(n_125),
.B1(n_126),
.B2(n_129),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_53),
.A2(n_40),
.B1(n_32),
.B2(n_31),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_54),
.B1(n_94),
.B2(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_60),
.A2(n_40),
.B1(n_32),
.B2(n_46),
.Y(n_129)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_78),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_70),
.A2(n_31),
.B1(n_42),
.B2(n_40),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_154),
.B1(n_28),
.B2(n_22),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_57),
.A2(n_42),
.B1(n_45),
.B2(n_29),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_91),
.B1(n_75),
.B2(n_56),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_78),
.B(n_29),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_151),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_47),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_152),
.B(n_79),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_71),
.A2(n_36),
.B1(n_47),
.B2(n_46),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_61),
.A2(n_36),
.B1(n_48),
.B2(n_41),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_99),
.B1(n_68),
.B2(n_48),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_158),
.Y(n_211)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_159),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_147),
.Y(n_160)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_162),
.Y(n_242)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_106),
.B(n_80),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_199),
.C(n_120),
.Y(n_209)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_166),
.A2(n_171),
.B1(n_201),
.B2(n_207),
.Y(n_221)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g241 ( 
.A(n_167),
.B(n_203),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

AO22x2_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_69),
.B1(n_98),
.B2(n_84),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_103),
.B1(n_130),
.B2(n_143),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_172),
.Y(n_231)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_39),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_39),
.B(n_37),
.C(n_28),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_176),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_101),
.B(n_37),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_22),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_180),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_138),
.B(n_21),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_181),
.B(n_185),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_184),
.A2(n_111),
.B1(n_139),
.B2(n_148),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_149),
.B(n_21),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

BUFx4f_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_140),
.A2(n_48),
.B(n_96),
.C(n_92),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_187),
.A2(n_110),
.B(n_145),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_190),
.Y(n_234)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_135),
.B(n_81),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_191),
.B(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_140),
.B(n_99),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_108),
.B(n_85),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_200),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_156),
.A2(n_83),
.B(n_59),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_65),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_103),
.A2(n_41),
.B1(n_87),
.B2(n_58),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_202),
.Y(n_226)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_206),
.Y(n_224)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_117),
.B(n_41),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_209),
.B(n_210),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_190),
.A2(n_124),
.B1(n_139),
.B2(n_111),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_222),
.A2(n_158),
.B(n_172),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_164),
.B(n_131),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_235),
.C(n_170),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_225),
.A2(n_229),
.B1(n_236),
.B2(n_247),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_164),
.B1(n_183),
.B2(n_166),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_128),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_174),
.B(n_133),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_245),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_179),
.A2(n_155),
.B(n_143),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_244),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_178),
.B(n_133),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_187),
.A2(n_126),
.B1(n_148),
.B2(n_153),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_224),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_249),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_218),
.B(n_163),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_252),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_176),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_240),
.B(n_157),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_253),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_220),
.A2(n_199),
.B1(n_170),
.B2(n_169),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_254),
.A2(n_257),
.B1(n_259),
.B2(n_266),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_204),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_255),
.B(n_256),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_223),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_221),
.A2(n_229),
.B1(n_235),
.B2(n_210),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_170),
.B1(n_175),
.B2(n_153),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_209),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_261),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_262),
.A2(n_213),
.B(n_228),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_195),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_263),
.Y(n_295)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_219),
.B(n_215),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_267),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_159),
.B1(n_173),
.B2(n_189),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_165),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_227),
.B(n_206),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_268),
.B(n_276),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_195),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_269),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_203),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_270),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_224),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_271),
.A2(n_232),
.B(n_242),
.Y(n_303)
);

AO22x1_ASAP7_75t_SL g272 ( 
.A1(n_227),
.A2(n_197),
.B1(n_186),
.B2(n_168),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_222),
.A2(n_161),
.B1(n_134),
.B2(n_132),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_275),
.A2(n_282),
.B1(n_211),
.B2(n_121),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_224),
.B(n_182),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_217),
.Y(n_279)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_238),
.B(n_182),
.Y(n_281)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_241),
.A2(n_202),
.B1(n_167),
.B2(n_104),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_228),
.B1(n_213),
.B2(n_211),
.Y(n_286)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_217),
.Y(n_284)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_284),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_286),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_287),
.A2(n_291),
.B1(n_307),
.B2(n_275),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_288),
.A2(n_296),
.B(n_303),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_257),
.A2(n_239),
.B1(n_243),
.B2(n_214),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_274),
.A2(n_213),
.B(n_242),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_274),
.A2(n_231),
.B(n_226),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_305),
.A2(n_306),
.B(n_313),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_274),
.A2(n_208),
.B(n_232),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_239),
.B1(n_243),
.B2(n_231),
.Y(n_307)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_270),
.A2(n_262),
.B(n_282),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_280),
.A2(n_177),
.B(n_208),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_315),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_261),
.A2(n_160),
.B(n_216),
.Y(n_315)
);

AO22x1_ASAP7_75t_L g316 ( 
.A1(n_259),
.A2(n_252),
.B1(n_278),
.B2(n_271),
.Y(n_316)
);

AO22x1_ASAP7_75t_L g344 ( 
.A1(n_316),
.A2(n_272),
.B1(n_216),
.B2(n_264),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_260),
.A2(n_230),
.B(n_216),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_318),
.B(n_249),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_256),
.C(n_251),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_325),
.C(n_346),
.Y(n_350)
);

XNOR2x1_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_251),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_320),
.B(n_288),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_253),
.Y(n_323)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_255),
.Y(n_324)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_324),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_267),
.C(n_265),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_293),
.Y(n_326)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_327),
.A2(n_313),
.B(n_314),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_297),
.B(n_304),
.Y(n_328)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_328),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_329),
.A2(n_334),
.B1(n_344),
.B2(n_292),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_305),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_338),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_290),
.B(n_250),
.Y(n_331)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_277),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_332),
.B(n_337),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_291),
.A2(n_278),
.B1(n_276),
.B2(n_268),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_293),
.Y(n_335)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_316),
.A2(n_266),
.B1(n_281),
.B2(n_272),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_336),
.A2(n_289),
.B1(n_285),
.B2(n_130),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_290),
.B(n_301),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_308),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_310),
.Y(n_339)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_339),
.Y(n_361)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_341),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_299),
.A2(n_284),
.B1(n_279),
.B2(n_269),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_342),
.A2(n_286),
.B(n_309),
.Y(n_370)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_343),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_294),
.B(n_263),
.C(n_258),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_295),
.B(n_188),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_349),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_294),
.B(n_104),
.C(n_188),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_296),
.C(n_306),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_272),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_302),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_364),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_357),
.A2(n_368),
.B1(n_336),
.B2(n_349),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_316),
.B(n_315),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_375),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_339),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_325),
.B(n_302),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_374),
.Y(n_401)
);

AOI21xp33_ASAP7_75t_L g363 ( 
.A1(n_323),
.A2(n_301),
.B(n_307),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_363),
.B(n_331),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_317),
.C(n_318),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_366),
.B(n_348),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_334),
.A2(n_292),
.B1(n_299),
.B2(n_303),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_369),
.B(n_333),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_370),
.A2(n_371),
.B(n_345),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_333),
.A2(n_340),
.B(n_322),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_320),
.B(n_311),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_340),
.A2(n_311),
.B(n_309),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_378),
.A2(n_329),
.B1(n_344),
.B2(n_342),
.Y(n_381)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_381),
.A2(n_399),
.B1(n_359),
.B2(n_370),
.Y(n_408)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_361),
.Y(n_382)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_383),
.B(n_386),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_324),
.Y(n_384)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_384),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_385),
.B(n_391),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_376),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_372),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_388),
.Y(n_404)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_398),
.C(n_377),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_357),
.A2(n_344),
.B1(n_327),
.B2(n_337),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_383),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_395),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_371),
.A2(n_328),
.B(n_330),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_394),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_376),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_396),
.B(n_403),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_343),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_374),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_373),
.B(n_338),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_368),
.A2(n_341),
.B1(n_335),
.B2(n_326),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_402),
.A2(n_356),
.B(n_375),
.Y(n_413)
);

FAx1_ASAP7_75t_SL g403 ( 
.A(n_369),
.B(n_321),
.CI(n_285),
.CON(n_403),
.SN(n_403)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_408),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_350),
.C(n_366),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_411),
.C(n_414),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_401),
.C(n_364),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_413),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_360),
.C(n_353),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_381),
.A2(n_367),
.B1(n_362),
.B2(n_365),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_415),
.A2(n_417),
.B1(n_418),
.B2(n_407),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_382),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_401),
.B(n_358),
.C(n_378),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_400),
.C(n_385),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_422),
.A2(n_379),
.B1(n_403),
.B2(n_392),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_405),
.A2(n_400),
.B(n_384),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_423),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_438),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_427),
.A2(n_212),
.B1(n_5),
.B2(n_6),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_380),
.C(n_402),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_428),
.B(n_429),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_380),
.C(n_394),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_380),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_431),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_420),
.A2(n_421),
.B(n_419),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_395),
.C(n_403),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_434),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_422),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_410),
.B(n_377),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_289),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_437),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_391),
.C(n_351),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_446),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_435),
.A2(n_413),
.B1(n_352),
.B2(n_351),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_445),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_406),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_406),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_321),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_449),
.A2(n_450),
.B1(n_4),
.B2(n_5),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_435),
.A2(n_432),
.B1(n_424),
.B2(n_426),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_212),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_5),
.C(n_6),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_448),
.B(n_424),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_456),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_452),
.A2(n_447),
.B(n_441),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_454),
.A2(n_7),
.B(n_8),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_442),
.B(n_4),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_461),
.Y(n_469)
);

AND2x2_ASAP7_75t_SL g458 ( 
.A(n_446),
.B(n_4),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_459),
.Y(n_471)
);

INVx11_ASAP7_75t_L g461 ( 
.A(n_442),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_5),
.C(n_6),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_463),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_439),
.A2(n_440),
.B1(n_444),
.B2(n_451),
.Y(n_463)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_454),
.A2(n_7),
.B(n_10),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_466),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_455),
.A2(n_11),
.B(n_12),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_470),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_460),
.A2(n_11),
.B(n_12),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_460),
.B(n_12),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_473),
.B(n_462),
.C(n_459),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_476),
.A2(n_477),
.B(n_472),
.Y(n_479)
);

AO21x1_ASAP7_75t_L g477 ( 
.A1(n_468),
.A2(n_464),
.B(n_461),
.Y(n_477)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_479),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_477),
.A2(n_469),
.B(n_471),
.Y(n_480)
);

AOI221xp5_ASAP7_75t_L g482 ( 
.A1(n_480),
.A2(n_481),
.B1(n_458),
.B2(n_13),
.C(n_14),
.Y(n_482)
);

AOI321xp33_ASAP7_75t_L g481 ( 
.A1(n_474),
.A2(n_458),
.A3(n_478),
.B1(n_475),
.B2(n_13),
.C(n_14),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_482),
.B(n_14),
.Y(n_484)
);

FAx1_ASAP7_75t_SL g485 ( 
.A(n_484),
.B(n_483),
.CI(n_14),
.CON(n_485),
.SN(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_485),
.B(n_384),
.Y(n_486)
);


endmodule