module fake_jpeg_5609_n_143 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_11),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_12),
.B1(n_19),
.B2(n_18),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_35),
.B1(n_16),
.B2(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_37),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_12),
.B1(n_19),
.B2(n_18),
.Y(n_35)
);

CKINVDCx12_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_27),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_20),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_12),
.B1(n_35),
.B2(n_29),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_46),
.B1(n_37),
.B2(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_52),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_20),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_17),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_54),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_57),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_31),
.B1(n_35),
.B2(n_52),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_53),
.B1(n_63),
.B2(n_55),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_63),
.B(n_42),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_49),
.B1(n_51),
.B2(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_75),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_45),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_73),
.C(n_56),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_49),
.C(n_40),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_55),
.B1(n_61),
.B2(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_60),
.Y(n_81)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

OAI22x1_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_62),
.B1(n_59),
.B2(n_56),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_32),
.B(n_17),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_82),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_33),
.B(n_53),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_60),
.C(n_61),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_74),
.C(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_91),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_93),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_32),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_8),
.Y(n_97)
);

BUFx12f_ASAP7_75t_SL g100 ( 
.A(n_97),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_77),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_79),
.B1(n_32),
.B2(n_13),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_102),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_13),
.B1(n_14),
.B2(n_27),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_9),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_17),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_89),
.C(n_96),
.Y(n_111)
);

OAI321xp33_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_14),
.A3(n_13),
.B1(n_10),
.B2(n_6),
.C(n_8),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_6),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_0),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_7),
.B1(n_9),
.B2(n_13),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_104),
.B1(n_2),
.B2(n_3),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_14),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_100),
.B(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_111),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_99),
.B1(n_105),
.B2(n_3),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_113),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_10),
.B(n_2),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_115),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_129),
.B(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_1),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_1),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_1),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_122),
.B1(n_121),
.B2(n_120),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_135),
.C(n_4),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_122),
.B(n_2),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_4),
.B(n_5),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_137),
.B(n_5),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_134),
.B1(n_5),
.B2(n_10),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_141),
.C(n_5),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_10),
.Y(n_143)
);


endmodule