module fake_jpeg_20055_n_40 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx12f_ASAP7_75t_SL g12 ( 
.A(n_5),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_19),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_7),
.B1(n_15),
.B2(n_16),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_13),
.Y(n_28)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_19),
.B(n_18),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_28),
.B1(n_15),
.B2(n_14),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_30),
.B(n_16),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_26),
.B1(n_20),
.B2(n_13),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_25),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_9),
.B(n_10),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_33),
.C(n_23),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_26),
.B1(n_9),
.B2(n_10),
.Y(n_39)
);

FAx1_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_37),
.CI(n_28),
.CON(n_40),
.SN(n_40)
);


endmodule