module real_aes_4712_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_1032, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_1032;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_666;
wire n_320;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_1025;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_523;
wire n_298;
wire n_996;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_1003;
wire n_1028;
wire n_533;
wire n_1000;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_649;
wire n_358;
wire n_293;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
HB1xp67_ASAP7_75t_L g292 ( .A(n_0), .Y(n_292) );
AND2x4_ASAP7_75t_L g786 ( .A(n_0), .B(n_787), .Y(n_786) );
AND2x4_ASAP7_75t_L g794 ( .A(n_0), .B(n_270), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_1), .A2(n_164), .B1(n_358), .B2(n_367), .Y(n_357) );
AO22x1_ASAP7_75t_L g829 ( .A1(n_2), .A2(n_3), .B1(n_793), .B2(n_811), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_4), .A2(n_204), .B1(n_783), .B2(n_790), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_5), .A2(n_35), .B1(n_503), .B2(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_6), .A2(n_279), .B1(n_540), .B2(n_541), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_7), .A2(n_188), .B1(n_387), .B2(n_477), .Y(n_476) );
AOI22x1_ASAP7_75t_L g1012 ( .A1(n_8), .A2(n_142), .B1(n_404), .B2(n_624), .Y(n_1012) );
CKINVDCx5p33_ASAP7_75t_R g665 ( .A(n_9), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_10), .A2(n_242), .B1(n_480), .B2(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_11), .A2(n_159), .B1(n_450), .B2(n_451), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_12), .A2(n_276), .B1(n_447), .B2(n_448), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_13), .A2(n_140), .B1(n_507), .B2(n_509), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_14), .A2(n_136), .B1(n_342), .B2(n_647), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_15), .Y(n_678) );
AO22x1_ASAP7_75t_L g745 ( .A1(n_16), .A2(n_24), .B1(n_746), .B2(n_747), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_17), .A2(n_122), .B1(n_820), .B2(n_835), .Y(n_834) );
AOI211xp5_ASAP7_75t_L g1002 ( .A1(n_18), .A2(n_1003), .B(n_1005), .C(n_1009), .Y(n_1002) );
XNOR2x1_ASAP7_75t_L g704 ( .A(n_19), .B(n_705), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g1006 ( .A1(n_20), .A2(n_36), .B1(n_342), .B2(n_424), .Y(n_1006) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_21), .A2(n_133), .B1(n_416), .B2(n_532), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_22), .A2(n_268), .B1(n_419), .B2(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_23), .A2(n_79), .B1(n_453), .B2(n_456), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_25), .A2(n_66), .B1(n_397), .B2(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g753 ( .A(n_26), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_27), .A2(n_174), .B1(n_490), .B2(n_491), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_28), .A2(n_72), .B1(n_585), .B2(n_586), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_29), .A2(n_94), .B1(n_465), .B2(n_466), .Y(n_707) );
INVx1_ASAP7_75t_L g768 ( .A(n_30), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_31), .A2(n_113), .B1(n_416), .B2(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g568 ( .A(n_32), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_33), .A2(n_182), .B1(n_399), .B2(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_34), .A2(n_46), .B1(n_624), .B2(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_37), .B(n_208), .Y(n_290) );
INVx1_ASAP7_75t_L g324 ( .A(n_37), .Y(n_324) );
INVxp67_ASAP7_75t_L g366 ( .A(n_37), .Y(n_366) );
OA22x2_ASAP7_75t_L g443 ( .A1(n_38), .A2(n_444), .B1(n_470), .B2(n_471), .Y(n_443) );
INVx1_ASAP7_75t_L g471 ( .A(n_38), .Y(n_471) );
INVx1_ASAP7_75t_L g487 ( .A(n_39), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_40), .A2(n_210), .B1(n_465), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_41), .A2(n_130), .B1(n_592), .B2(n_593), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_42), .A2(n_54), .B1(n_402), .B2(n_404), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_43), .A2(n_151), .B1(n_377), .B2(n_690), .Y(n_689) );
AOI21xp33_ASAP7_75t_SL g485 ( .A1(n_44), .A2(n_304), .B(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_45), .A2(n_103), .B1(n_624), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_47), .A2(n_138), .B1(n_469), .B2(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_48), .B(n_424), .Y(n_505) );
INVx1_ASAP7_75t_L g734 ( .A(n_49), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_50), .A2(n_468), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_51), .B(n_309), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_52), .A2(n_112), .B1(n_649), .B2(n_651), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_53), .A2(n_235), .B1(n_416), .B2(n_417), .Y(n_515) );
INVx1_ASAP7_75t_L g766 ( .A(n_55), .Y(n_766) );
INVx1_ASAP7_75t_L g335 ( .A(n_56), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_57), .A2(n_218), .B1(n_460), .B2(n_466), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_58), .A2(n_176), .B1(n_799), .B2(n_811), .Y(n_825) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_59), .A2(n_567), .B(n_733), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_60), .A2(n_134), .B1(n_397), .B2(n_399), .Y(n_396) );
INVx2_ASAP7_75t_L g287 ( .A(n_61), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_62), .A2(n_101), .B1(n_387), .B2(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g327 ( .A(n_63), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_64), .A2(n_172), .B1(n_465), .B2(n_469), .Y(n_730) );
INVx1_ASAP7_75t_L g785 ( .A(n_65), .Y(n_785) );
AND2x4_ASAP7_75t_L g791 ( .A(n_65), .B(n_287), .Y(n_791) );
INVx1_ASAP7_75t_SL g833 ( .A(n_65), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g1013 ( .A1(n_67), .A2(n_236), .B1(n_651), .B2(n_1014), .C(n_1015), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_68), .A2(n_195), .B1(n_793), .B2(n_795), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_69), .A2(n_98), .B1(n_465), .B2(n_466), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_70), .A2(n_201), .B1(n_404), .B2(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g770 ( .A(n_71), .Y(n_770) );
INVx1_ASAP7_75t_L g499 ( .A(n_73), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_74), .A2(n_249), .B1(n_421), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_75), .A2(n_180), .B1(n_793), .B2(n_811), .Y(n_842) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_76), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_77), .A2(n_85), .B1(n_416), .B2(n_417), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_78), .A2(n_216), .B1(n_450), .B2(n_451), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_80), .A2(n_194), .B1(n_421), .B2(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g762 ( .A(n_81), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_82), .A2(n_260), .B1(n_460), .B2(n_469), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_83), .A2(n_280), .B1(n_447), .B2(n_456), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_84), .A2(n_165), .B1(n_783), .B2(n_818), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_86), .A2(n_169), .B1(n_413), .B2(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_87), .A2(n_135), .B1(n_377), .B2(n_413), .Y(n_626) );
INVx1_ASAP7_75t_L g712 ( .A(n_88), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_89), .A2(n_238), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_90), .A2(n_119), .B1(n_453), .B2(n_456), .Y(n_557) );
INVx1_ASAP7_75t_L g313 ( .A(n_91), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_91), .B(n_207), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_92), .A2(n_269), .B1(n_387), .B2(n_414), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_93), .A2(n_267), .B1(n_593), .B2(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g671 ( .A(n_95), .Y(n_671) );
AO22x1_ASAP7_75t_L g614 ( .A1(n_96), .A2(n_118), .B1(n_480), .B2(n_504), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_97), .A2(n_252), .B1(n_448), .B2(n_457), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_99), .A2(n_155), .B1(n_543), .B2(n_545), .C(n_547), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_100), .A2(n_145), .B1(n_460), .B2(n_469), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_102), .A2(n_612), .B(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_104), .A2(n_202), .B1(n_387), .B2(n_414), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_105), .A2(n_173), .B1(n_783), .B2(n_788), .Y(n_797) );
INVx2_ASAP7_75t_R g298 ( .A(n_106), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_107), .A2(n_272), .B1(n_447), .B2(n_448), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_108), .A2(n_120), .B1(n_783), .B2(n_790), .Y(n_843) );
AOI221xp5_ASAP7_75t_SL g458 ( .A1(n_109), .A2(n_244), .B1(n_459), .B2(n_460), .C(n_461), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_110), .B(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_111), .A2(n_154), .B1(n_530), .B2(n_532), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_114), .A2(n_237), .B1(n_404), .B2(n_419), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_115), .A2(n_222), .B1(n_429), .B2(n_1008), .Y(n_1007) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_116), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_117), .A2(n_183), .B1(n_465), .B2(n_466), .C(n_467), .Y(n_464) );
CKINVDCx14_ASAP7_75t_R g1000 ( .A(n_120), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_120), .A2(n_1022), .B1(n_1024), .B2(n_1028), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_121), .A2(n_209), .B1(n_781), .B2(n_788), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_123), .B(n_595), .Y(n_729) );
INVx1_ASAP7_75t_L g681 ( .A(n_124), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_125), .A2(n_185), .B1(n_595), .B2(n_597), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_126), .A2(n_259), .B1(n_783), .B2(n_790), .Y(n_826) );
INVx1_ASAP7_75t_L g409 ( .A(n_127), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_128), .A2(n_158), .B1(n_456), .B2(n_457), .Y(n_455) );
NAND2xp33_ASAP7_75t_L g580 ( .A(n_129), .B(n_541), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_131), .A2(n_193), .B1(n_450), .B2(n_451), .Y(n_739) );
INVx1_ASAP7_75t_L g656 ( .A(n_132), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_137), .A2(n_219), .B1(n_601), .B2(n_621), .Y(n_749) );
AO22x1_ASAP7_75t_L g1015 ( .A1(n_139), .A2(n_196), .B1(n_377), .B2(n_758), .Y(n_1015) );
INVx1_ASAP7_75t_L g761 ( .A(n_141), .Y(n_761) );
AO22x1_ASAP7_75t_L g1009 ( .A1(n_143), .A2(n_256), .B1(n_387), .B2(n_477), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_144), .A2(n_149), .B1(n_413), .B2(n_414), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_146), .A2(n_212), .B1(n_447), .B2(n_448), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_147), .A2(n_192), .B1(n_453), .B2(n_454), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g376 ( .A1(n_148), .A2(n_200), .B1(n_377), .B2(n_382), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_150), .A2(n_254), .B1(n_790), .B2(n_832), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_152), .A2(n_251), .B1(n_416), .B2(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g302 ( .A(n_153), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_156), .A2(n_1025), .B1(n_1026), .B2(n_1027), .Y(n_1024) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_156), .Y(n_1025) );
AO22x1_ASAP7_75t_L g467 ( .A1(n_157), .A2(n_234), .B1(n_468), .B2(n_469), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_160), .A2(n_220), .B1(n_696), .B2(n_698), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_161), .A2(n_239), .B1(n_454), .B2(n_457), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_162), .A2(n_177), .B1(n_429), .B2(n_480), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_163), .A2(n_243), .B1(n_454), .B2(n_457), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_166), .A2(n_168), .B1(n_397), .B2(n_399), .Y(n_475) );
INVx1_ASAP7_75t_L g340 ( .A(n_167), .Y(n_340) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_170), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_171), .A2(n_221), .B1(n_799), .B2(n_820), .Y(n_819) );
XOR2x2_ASAP7_75t_L g742 ( .A(n_173), .B(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_175), .B(n_597), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_178), .A2(n_258), .B1(n_377), .B2(n_413), .Y(n_638) );
AO221x2_ASAP7_75t_L g828 ( .A1(n_179), .A2(n_230), .B1(n_783), .B2(n_818), .C(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g427 ( .A(n_181), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_184), .A2(n_241), .B1(n_304), .B2(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_186), .A2(n_248), .B1(n_621), .B2(n_693), .Y(n_692) );
OA22x2_ASAP7_75t_L g307 ( .A1(n_187), .A2(n_208), .B1(n_308), .B2(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g348 ( .A(n_187), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_189), .A2(n_206), .B1(n_494), .B2(n_601), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_190), .A2(n_226), .B1(n_424), .B2(n_425), .C(n_426), .Y(n_423) );
INVx1_ASAP7_75t_L g565 ( .A(n_191), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_197), .A2(n_266), .B1(n_795), .B2(n_799), .Y(n_798) );
AOI221x1_ASAP7_75t_L g581 ( .A1(n_198), .A2(n_247), .B1(n_540), .B2(n_551), .C(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g1010 ( .A1(n_199), .A2(n_213), .B1(n_621), .B2(n_640), .C(n_1011), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_203), .A2(n_271), .B1(n_799), .B2(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_205), .A2(n_245), .B1(n_397), .B2(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g326 ( .A(n_207), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_207), .B(n_346), .Y(n_373) );
OAI21xp33_ASAP7_75t_L g349 ( .A1(n_208), .A2(n_224), .B(n_350), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g608 ( .A(n_209), .Y(n_608) );
AND2x2_ASAP7_75t_L g582 ( .A(n_211), .B(n_531), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g472 ( .A(n_214), .B(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_215), .A2(n_227), .B1(n_342), .B2(n_618), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_217), .A2(n_246), .B1(n_402), .B2(n_404), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_223), .A2(n_233), .B1(n_431), .B2(n_432), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_224), .B(n_262), .Y(n_291) );
INVx1_ASAP7_75t_L g315 ( .A(n_224), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_225), .A2(n_257), .B1(n_450), .B2(n_451), .Y(n_558) );
INVx1_ASAP7_75t_L g548 ( .A(n_228), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_229), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g726 ( .A(n_230), .Y(n_726) );
XNOR2x1_ASAP7_75t_L g526 ( .A(n_231), .B(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_232), .A2(n_275), .B1(n_431), .B2(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g352 ( .A(n_240), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_250), .B(n_425), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_253), .A2(n_265), .B1(n_419), .B2(n_520), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g578 ( .A(n_254), .B(n_579), .C(n_583), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_254), .A2(n_583), .B1(n_590), .B2(n_1032), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_254), .A2(n_579), .B(n_599), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_255), .A2(n_273), .B1(n_304), .B2(n_342), .Y(n_434) );
INVx1_ASAP7_75t_L g756 ( .A(n_261), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_262), .B(n_319), .Y(n_318) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_263), .A2(n_460), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_264), .B(n_490), .Y(n_709) );
INVx1_ASAP7_75t_L g787 ( .A(n_270), .Y(n_787) );
INVx1_ASAP7_75t_L g701 ( .A(n_274), .Y(n_701) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_277), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_278), .A2(n_612), .B(n_614), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_293), .B(n_776), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx4_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
NAND3xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .C(n_292), .Y(n_284) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_285), .B(n_1019), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_285), .B(n_1020), .Y(n_1023) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OA21x2_ASAP7_75t_L g1029 ( .A1(n_286), .A2(n_833), .B(n_1030), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g784 ( .A(n_287), .B(n_785), .Y(n_784) );
AND3x4_ASAP7_75t_L g832 ( .A(n_287), .B(n_786), .C(n_833), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_288), .B(n_1020), .Y(n_1019) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AO21x2_ASAP7_75t_L g370 ( .A1(n_289), .A2(n_371), .B(n_372), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_L g1020 ( .A(n_292), .Y(n_1020) );
XNOR2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_523), .Y(n_293) );
OA22x2_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_439), .B1(n_521), .B2(n_522), .Y(n_294) );
INVx1_ASAP7_75t_L g522 ( .A(n_295), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_407), .B1(n_435), .B2(n_436), .Y(n_295) );
INVx2_ASAP7_75t_L g435 ( .A(n_296), .Y(n_435) );
HB1xp67_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
XNOR2x1_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_374), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_334), .C(n_351), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B1(n_327), .B2(n_328), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_303), .A2(n_665), .B1(n_666), .B2(n_667), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_303), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
INVx4_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g508 ( .A(n_305), .Y(n_508) );
BUFx3_ASAP7_75t_L g592 ( .A(n_305), .Y(n_592) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_316), .Y(n_305) );
AND2x4_ASAP7_75t_L g337 ( .A(n_306), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g460 ( .A(n_306), .B(n_316), .Y(n_460) );
AND2x2_ASAP7_75t_L g567 ( .A(n_306), .B(n_338), .Y(n_567) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_310), .Y(n_306) );
AND2x2_ASAP7_75t_L g333 ( .A(n_307), .B(n_311), .Y(n_333) );
AND2x2_ASAP7_75t_L g364 ( .A(n_307), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g390 ( .A(n_307), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_308), .B(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp33_ASAP7_75t_L g312 ( .A(n_309), .B(n_313), .Y(n_312) );
INVx3_ASAP7_75t_L g319 ( .A(n_309), .Y(n_319) );
NAND2xp33_ASAP7_75t_L g325 ( .A(n_309), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g350 ( .A(n_309), .Y(n_350) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_309), .Y(n_362) );
AND2x4_ASAP7_75t_L g389 ( .A(n_310), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_313), .B(n_348), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_315), .A2(n_350), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g332 ( .A(n_316), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g398 ( .A(n_316), .B(n_389), .Y(n_398) );
AND2x4_ASAP7_75t_L g450 ( .A(n_316), .B(n_389), .Y(n_450) );
AND2x4_ASAP7_75t_L g465 ( .A(n_316), .B(n_333), .Y(n_465) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_321), .Y(n_316) );
INVx2_ASAP7_75t_L g339 ( .A(n_317), .Y(n_339) );
AND2x2_ASAP7_75t_L g360 ( .A(n_317), .B(n_361), .Y(n_360) );
AND2x4_ASAP7_75t_L g379 ( .A(n_317), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g385 ( .A(n_317), .B(n_381), .Y(n_385) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_319), .B(n_324), .Y(n_323) );
INVxp67_ASAP7_75t_L g346 ( .A(n_319), .Y(n_346) );
NAND3xp33_ASAP7_75t_L g372 ( .A(n_320), .B(n_345), .C(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g338 ( .A(n_321), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g381 ( .A(n_322), .Y(n_381) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g616 ( .A(n_330), .Y(n_616) );
INVx2_ASAP7_75t_L g764 ( .A(n_330), .Y(n_764) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g431 ( .A(n_331), .Y(n_431) );
INVx2_ASAP7_75t_L g585 ( .A(n_331), .Y(n_585) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_332), .Y(n_511) );
BUFx3_ASAP7_75t_L g669 ( .A(n_332), .Y(n_669) );
AND2x2_ASAP7_75t_L g356 ( .A(n_333), .B(n_338), .Y(n_356) );
AND2x2_ASAP7_75t_L g378 ( .A(n_333), .B(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g383 ( .A(n_333), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g447 ( .A(n_333), .B(n_379), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_333), .B(n_391), .Y(n_448) );
AND2x2_ASAP7_75t_L g468 ( .A(n_333), .B(n_338), .Y(n_468) );
AND2x2_ASAP7_75t_L g531 ( .A(n_333), .B(n_379), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_340), .B2(n_341), .Y(n_334) );
INVx3_ASAP7_75t_L g424 ( .A(n_336), .Y(n_424) );
INVx2_ASAP7_75t_L g618 ( .A(n_336), .Y(n_618) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_337), .Y(n_459) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_337), .Y(n_490) );
INVx2_ASAP7_75t_L g544 ( .A(n_337), .Y(n_544) );
BUFx3_ASAP7_75t_L g588 ( .A(n_337), .Y(n_588) );
AND2x4_ASAP7_75t_L g343 ( .A(n_338), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g400 ( .A(n_338), .B(n_389), .Y(n_400) );
AND2x4_ASAP7_75t_L g451 ( .A(n_338), .B(n_389), .Y(n_451) );
AND2x4_ASAP7_75t_L g469 ( .A(n_338), .B(n_344), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_341), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_765) );
INVx4_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g492 ( .A(n_343), .Y(n_492) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_343), .Y(n_586) );
AND2x4_ASAP7_75t_L g394 ( .A(n_344), .B(n_391), .Y(n_394) );
AND2x4_ASAP7_75t_L g406 ( .A(n_344), .B(n_379), .Y(n_406) );
AND2x4_ASAP7_75t_L g456 ( .A(n_344), .B(n_379), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_344), .B(n_391), .Y(n_457) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B(n_357), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx3_ASAP7_75t_SL g425 ( .A(n_355), .Y(n_425) );
INVx2_ASAP7_75t_L g503 ( .A(n_355), .Y(n_503) );
INVx2_ASAP7_75t_L g1004 ( .A(n_355), .Y(n_1004) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx3_ASAP7_75t_L g561 ( .A(n_356), .Y(n_561) );
INVx2_ASAP7_75t_L g596 ( .A(n_356), .Y(n_596) );
BUFx4f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx5_ASAP7_75t_L g433 ( .A(n_359), .Y(n_433) );
BUFx2_ASAP7_75t_L g480 ( .A(n_359), .Y(n_480) );
BUFx2_ASAP7_75t_L g655 ( .A(n_359), .Y(n_655) );
AND2x4_ASAP7_75t_L g359 ( .A(n_360), .B(n_364), .Y(n_359) );
AND2x2_ASAP7_75t_L g466 ( .A(n_360), .B(n_364), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g371 ( .A(n_362), .Y(n_371) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx4_ASAP7_75t_L g429 ( .A(n_368), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_368), .B(n_734), .Y(n_733) );
INVx4_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx3_ASAP7_75t_L g488 ( .A(n_369), .Y(n_488) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_370), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_395), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_386), .Y(n_375) );
BUFx8_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
AND2x4_ASAP7_75t_L g403 ( .A(n_379), .B(n_389), .Y(n_403) );
AND2x4_ASAP7_75t_L g453 ( .A(n_379), .B(n_389), .Y(n_453) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx3_ASAP7_75t_L g690 ( .A(n_382), .Y(n_690) );
BUFx12f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_383), .Y(n_413) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_383), .Y(n_482) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_383), .Y(n_532) );
BUFx3_ASAP7_75t_L g758 ( .A(n_383), .Y(n_758) );
AND2x4_ASAP7_75t_L g454 ( .A(n_384), .B(n_389), .Y(n_454) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g391 ( .A(n_385), .Y(n_391) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_388), .Y(n_417) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_388), .Y(n_540) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_388), .Y(n_697) );
AND2x4_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g477 ( .A(n_393), .Y(n_477) );
INVx3_ASAP7_75t_L g514 ( .A(n_393), .Y(n_514) );
INVx5_ASAP7_75t_L g541 ( .A(n_393), .Y(n_541) );
INVx2_ASAP7_75t_L g700 ( .A(n_393), .Y(n_700) );
INVx6_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx12f_ASAP7_75t_L g414 ( .A(n_394), .Y(n_414) );
NAND2xp33_ASAP7_75t_L g395 ( .A(n_396), .B(n_401), .Y(n_395) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx3_ASAP7_75t_L g518 ( .A(n_398), .Y(n_518) );
BUFx12f_ASAP7_75t_L g551 ( .A(n_398), .Y(n_551) );
BUFx5_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_400), .Y(n_421) );
BUFx3_ASAP7_75t_L g601 ( .A(n_400), .Y(n_601) );
INVx1_ASAP7_75t_L g642 ( .A(n_400), .Y(n_642) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx12f_ASAP7_75t_L g416 ( .A(n_403), .Y(n_416) );
INVx4_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx4_ASAP7_75t_L g494 ( .A(n_405), .Y(n_494) );
INVx2_ASAP7_75t_L g520 ( .A(n_405), .Y(n_520) );
INVx2_ASAP7_75t_SL g534 ( .A(n_405), .Y(n_534) );
INVx4_ASAP7_75t_L g688 ( .A(n_405), .Y(n_688) );
INVx1_ASAP7_75t_L g751 ( .A(n_405), .Y(n_751) );
INVx8_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g438 ( .A(n_408), .Y(n_438) );
XNOR2x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
NOR2x1_ASAP7_75t_L g410 ( .A(n_411), .B(n_422), .Y(n_410) );
NAND4xp25_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .C(n_418), .D(n_420), .Y(n_411) );
BUFx12f_ASAP7_75t_L g624 ( .A(n_416), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_430), .C(n_434), .Y(n_422) );
INVx1_ASAP7_75t_L g771 ( .A(n_425), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g536 ( .A(n_433), .Y(n_536) );
INVx4_ASAP7_75t_L g593 ( .A(n_433), .Y(n_593) );
INVx3_ASAP7_75t_L g1008 ( .A(n_433), .Y(n_1008) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g521 ( .A(n_439), .Y(n_521) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
XOR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_496), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B1(n_472), .B2(n_495), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g470 ( .A(n_444), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_458), .C(n_464), .Y(n_444) );
AND4x1_ASAP7_75t_L g445 ( .A(n_446), .B(n_449), .C(n_452), .D(n_455), .Y(n_445) );
BUFx3_ASAP7_75t_L g647 ( .A(n_459), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g504 ( .A(n_462), .Y(n_504) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_462), .Y(n_549) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_462), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_462), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g546 ( .A(n_468), .Y(n_546) );
INVx1_ASAP7_75t_L g495 ( .A(n_472), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .C(n_483), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_479), .B(n_481), .Y(n_478) );
NAND4xp25_ASAP7_75t_SL g483 ( .A(n_484), .B(n_485), .C(n_489), .D(n_493), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_488), .B(n_565), .Y(n_564) );
INVx4_ASAP7_75t_L g676 ( .A(n_488), .Y(n_676) );
BUFx3_ASAP7_75t_L g680 ( .A(n_490), .Y(n_680) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g509 ( .A(n_492), .Y(n_509) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
XNOR2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
NOR2x1_ASAP7_75t_L g500 ( .A(n_501), .B(n_512), .Y(n_500) );
NAND4xp25_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .C(n_506), .D(n_510), .Y(n_501) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g512 ( .A(n_513), .B(n_515), .C(n_516), .D(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g622 ( .A(n_518), .Y(n_622) );
XNOR2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_629), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_571), .B1(n_627), .B2(n_628), .Y(n_524) );
INVx2_ASAP7_75t_L g627 ( .A(n_525), .Y(n_627) );
OA22x2_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_552), .B1(n_569), .B2(n_570), .Y(n_525) );
INVx1_ASAP7_75t_L g569 ( .A(n_526), .Y(n_569) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_538), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .C(n_535), .D(n_537), .Y(n_528) );
BUFx4f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_531), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .C(n_550), .Y(n_538) );
BUFx3_ASAP7_75t_L g746 ( .A(n_540), .Y(n_746) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g570 ( .A(n_552), .Y(n_570) );
XOR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_568), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g553 ( .A(n_554), .B(n_559), .Y(n_553) );
NAND4xp25_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .C(n_557), .D(n_558), .Y(n_554) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .C(n_563), .D(n_566), .Y(n_559) );
INVx1_ASAP7_75t_L g613 ( .A(n_561), .Y(n_613) );
INVx1_ASAP7_75t_L g628 ( .A(n_571), .Y(n_628) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_606), .B2(n_607), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AO22x2_ASAP7_75t_L g722 ( .A1(n_577), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_577), .Y(n_723) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_589), .B(n_603), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_584), .B(n_587), .Y(n_583) );
BUFx3_ASAP7_75t_L g651 ( .A(n_585), .Y(n_651) );
BUFx3_ASAP7_75t_L g683 ( .A(n_586), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_599), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
INVx2_ASAP7_75t_L g650 ( .A(n_592), .Y(n_650) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_592), .Y(n_1014) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_596), .Y(n_674) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NAND2x1_ASAP7_75t_SL g599 ( .A(n_600), .B(n_602), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
XNOR2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g609 ( .A(n_610), .B(n_619), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_615), .C(n_617), .Y(n_610) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .C(n_625), .D(n_626), .Y(n_619) );
BUFx4f_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_719), .B1(n_720), .B2(n_775), .Y(n_629) );
INVx1_ASAP7_75t_L g775 ( .A(n_630), .Y(n_775) );
XNOR2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_659), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AO21x2_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_658), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g658 ( .A(n_633), .B(n_636), .C(n_645), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_644), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND4xp25_ASAP7_75t_SL g636 ( .A(n_637), .B(n_638), .C(n_639), .D(n_643), .Y(n_636) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g694 ( .A(n_641), .Y(n_694) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .C(n_652), .Y(n_645) );
INVx1_ASAP7_75t_L g767 ( .A(n_647), .Y(n_767) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_656), .B(n_657), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_702), .B2(n_718), .Y(n_659) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
XOR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_701), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_684), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_670), .C(n_677), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI21xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B(n_675), .Y(n_670) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_681), .B2(n_682), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NOR2xp67_ASAP7_75t_L g684 ( .A(n_685), .B(n_691), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .Y(n_685) );
BUFx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_695), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_700), .Y(n_747) );
INVx1_ASAP7_75t_L g718 ( .A(n_702), .Y(n_718) );
HB1xp67_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_713), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .C(n_709), .D(n_710), .Y(n_706) );
NAND4xp25_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .C(n_716), .D(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_741), .B1(n_773), .B2(n_774), .Y(n_720) );
INVx1_ASAP7_75t_L g773 ( .A(n_721), .Y(n_773) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AO21x2_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_740), .Y(n_725) );
NOR3xp33_ASAP7_75t_SL g740 ( .A(n_726), .B(n_728), .C(n_735), .Y(n_740) );
OR2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_735), .Y(n_727) );
NAND4xp75_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .C(n_731), .D(n_732), .Y(n_728) );
NAND4xp25_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .C(n_738), .D(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g774 ( .A(n_741), .Y(n_774) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_759), .Y(n_743) );
NOR3xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_748), .C(n_752), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_756), .B2(n_757), .Y(n_752) );
INVxp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_765), .C(n_769), .Y(n_759) );
INVxp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OAI21xp33_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B(n_772), .Y(n_769) );
OAI221xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_996), .B1(n_998), .B2(n_1016), .C(n_1021), .Y(n_776) );
AOI211xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_800), .B(n_868), .C(n_962), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_779), .B(n_796), .Y(n_778) );
AOI221xp5_ASAP7_75t_L g894 ( .A1(n_779), .A2(n_837), .B1(n_895), .B2(n_897), .C(n_920), .Y(n_894) );
CKINVDCx5p33_ASAP7_75t_R g922 ( .A(n_779), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_779), .B(n_839), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_779), .A2(n_896), .B1(n_904), .B2(n_909), .C(n_969), .Y(n_968) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_792), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_784), .B(n_786), .Y(n_783) );
AND2x4_ASAP7_75t_L g793 ( .A(n_784), .B(n_794), .Y(n_793) );
AND2x2_ASAP7_75t_L g799 ( .A(n_784), .B(n_794), .Y(n_799) );
AND2x2_ASAP7_75t_L g835 ( .A(n_784), .B(n_794), .Y(n_835) );
AND2x4_ASAP7_75t_L g790 ( .A(n_786), .B(n_791), .Y(n_790) );
AND2x4_ASAP7_75t_L g818 ( .A(n_786), .B(n_791), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_786), .B(n_791), .Y(n_997) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_786), .Y(n_1030) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
AND2x4_ASAP7_75t_L g795 ( .A(n_791), .B(n_794), .Y(n_795) );
AND2x2_ASAP7_75t_L g811 ( .A(n_791), .B(n_794), .Y(n_811) );
AND2x2_ASAP7_75t_L g820 ( .A(n_791), .B(n_794), .Y(n_820) );
INVx1_ASAP7_75t_L g893 ( .A(n_796), .Y(n_893) );
INVx4_ASAP7_75t_L g900 ( .A(n_796), .Y(n_900) );
AND2x2_ASAP7_75t_L g904 ( .A(n_796), .B(n_841), .Y(n_904) );
NAND3xp33_ASAP7_75t_L g906 ( .A(n_796), .B(n_856), .C(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g909 ( .A(n_796), .B(n_910), .Y(n_909) );
AND2x2_ASAP7_75t_L g961 ( .A(n_796), .B(n_891), .Y(n_961) );
AND2x2_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
NAND4xp25_ASAP7_75t_L g800 ( .A(n_801), .B(n_836), .C(n_858), .D(n_864), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_813), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g946 ( .A(n_804), .B(n_904), .Y(n_946) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g860 ( .A(n_805), .Y(n_860) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_806), .Y(n_881) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OR2x2_ASAP7_75t_L g892 ( .A(n_808), .B(n_840), .Y(n_892) );
INVx2_ASAP7_75t_L g910 ( .A(n_808), .Y(n_910) );
INVx4_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
OR2x2_ASAP7_75t_L g866 ( .A(n_809), .B(n_840), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_809), .B(n_878), .Y(n_877) );
OR2x2_ASAP7_75t_L g901 ( .A(n_809), .B(n_841), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g907 ( .A(n_809), .B(n_824), .Y(n_907) );
AND2x2_ASAP7_75t_L g953 ( .A(n_809), .B(n_840), .Y(n_953) );
AND2x2_ASAP7_75t_L g809 ( .A(n_810), .B(n_812), .Y(n_809) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_821), .Y(n_814) );
AND2x2_ASAP7_75t_L g848 ( .A(n_815), .B(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_815), .B(n_856), .Y(n_855) );
AND2x2_ASAP7_75t_L g874 ( .A(n_815), .B(n_824), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_815), .B(n_857), .Y(n_912) );
AND2x2_ASAP7_75t_L g914 ( .A(n_815), .B(n_883), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_815), .B(n_850), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_815), .B(n_944), .Y(n_965) );
AND2x2_ASAP7_75t_L g979 ( .A(n_815), .B(n_828), .Y(n_979) );
CKINVDCx6p67_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g852 ( .A(n_816), .B(n_830), .Y(n_852) );
AND2x2_ASAP7_75t_L g862 ( .A(n_816), .B(n_822), .Y(n_862) );
AND2x2_ASAP7_75t_L g872 ( .A(n_816), .B(n_849), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_816), .B(n_857), .Y(n_888) );
AND2x2_ASAP7_75t_L g896 ( .A(n_816), .B(n_883), .Y(n_896) );
AND2x2_ASAP7_75t_L g903 ( .A(n_816), .B(n_863), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_816), .B(n_828), .Y(n_933) );
AND2x2_ASAP7_75t_L g943 ( .A(n_816), .B(n_944), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_816), .B(n_850), .Y(n_955) );
AND2x2_ASAP7_75t_L g816 ( .A(n_817), .B(n_819), .Y(n_816) );
INVx1_ASAP7_75t_L g993 ( .A(n_821), .Y(n_993) );
NOR2x1_ASAP7_75t_L g821 ( .A(n_822), .B(n_827), .Y(n_821) );
AND2x2_ASAP7_75t_L g853 ( .A(n_822), .B(n_854), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g976 ( .A(n_822), .B(n_952), .Y(n_976) );
INVx3_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g844 ( .A(n_823), .B(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_823), .B(n_848), .Y(n_885) );
AND2x2_ASAP7_75t_L g939 ( .A(n_823), .B(n_940), .Y(n_939) );
AND2x2_ASAP7_75t_L g944 ( .A(n_823), .B(n_863), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_823), .B(n_955), .Y(n_954) );
INVx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g878 ( .A(n_824), .Y(n_878) );
INVx2_ASAP7_75t_L g890 ( .A(n_824), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_824), .B(n_933), .Y(n_932) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_824), .B(n_936), .Y(n_935) );
AND2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
INVx1_ASAP7_75t_L g883 ( .A(n_827), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g983 ( .A(n_827), .B(n_878), .Y(n_983) );
OR2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_830), .Y(n_827) );
AND2x2_ASAP7_75t_L g849 ( .A(n_828), .B(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g857 ( .A(n_828), .Y(n_857) );
AND2x2_ASAP7_75t_L g863 ( .A(n_828), .B(n_830), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_828), .B(n_862), .Y(n_921) );
INVx1_ASAP7_75t_L g850 ( .A(n_830), .Y(n_850) );
AND2x2_ASAP7_75t_L g856 ( .A(n_830), .B(n_857), .Y(n_856) );
OAI21xp33_ASAP7_75t_L g974 ( .A1(n_830), .A2(n_975), .B(n_977), .Y(n_974) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_834), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_844), .B2(n_853), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
OAI21xp33_ASAP7_75t_L g884 ( .A1(n_838), .A2(n_885), .B(n_886), .Y(n_884) );
INVx3_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
AOI21xp33_ASAP7_75t_L g879 ( .A1(n_839), .A2(n_861), .B(n_880), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_839), .B(n_900), .Y(n_981) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVxp67_ASAP7_75t_L g917 ( .A(n_840), .Y(n_917) );
AND2x2_ASAP7_75t_L g973 ( .A(n_840), .B(n_900), .Y(n_973) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_SL g846 ( .A(n_847), .B(n_851), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_848), .B(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g936 ( .A(n_849), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_849), .B(n_862), .Y(n_970) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_852), .B(n_890), .Y(n_919) );
OAI221xp5_ASAP7_75t_L g923 ( .A1(n_853), .A2(n_924), .B1(n_930), .B2(n_937), .C(n_941), .Y(n_923) );
INVx2_ASAP7_75t_L g867 ( .A(n_854), .Y(n_867) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_856), .B(n_899), .Y(n_898) );
AOI221xp5_ASAP7_75t_L g982 ( .A1(n_856), .A2(n_862), .B1(n_876), .B2(n_948), .C(n_983), .Y(n_982) );
INVxp67_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_860), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
AND2x2_ASAP7_75t_L g882 ( .A(n_862), .B(n_883), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_863), .B(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g948 ( .A(n_863), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g990 ( .A1(n_863), .A2(n_950), .B(n_991), .Y(n_990) );
INVxp67_ASAP7_75t_SL g864 ( .A(n_865), .Y(n_864) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
A2O1A1Ixp33_ASAP7_75t_L g870 ( .A1(n_866), .A2(n_871), .B(n_873), .C(n_875), .Y(n_870) );
AOI211xp5_ASAP7_75t_L g920 ( .A1(n_866), .A2(n_885), .B(n_921), .C(n_922), .Y(n_920) );
INVx1_ASAP7_75t_L g940 ( .A(n_866), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_866), .B(n_967), .Y(n_966) );
NAND4xp25_ASAP7_75t_L g868 ( .A(n_869), .B(n_894), .C(n_923), .D(n_942), .Y(n_868) );
OAI31xp33_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_879), .A3(n_884), .B(n_893), .Y(n_869) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g959 ( .A(n_873), .Y(n_959) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
AND2x2_ASAP7_75t_L g895 ( .A(n_878), .B(n_896), .Y(n_895) );
AND2x2_ASAP7_75t_L g978 ( .A(n_878), .B(n_979), .Y(n_978) );
OAI211xp5_ASAP7_75t_SL g924 ( .A1(n_880), .A2(n_925), .B(n_926), .C(n_929), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_883), .B(n_939), .Y(n_938) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_887), .B(n_889), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_888), .A2(n_960), .B1(n_965), .B2(n_966), .C(n_968), .Y(n_964) );
AND2x2_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
OAI21xp33_ASAP7_75t_L g911 ( .A1(n_890), .A2(n_912), .B(n_913), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_890), .B(n_927), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g950 ( .A(n_890), .B(n_901), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_890), .B(n_928), .Y(n_957) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g930 ( .A1(n_892), .A2(n_901), .B1(n_922), .B2(n_931), .C(n_934), .Y(n_930) );
O2A1O1Ixp33_ASAP7_75t_SL g962 ( .A1(n_893), .A2(n_963), .B(n_971), .C(n_985), .Y(n_962) );
INVx1_ASAP7_75t_L g984 ( .A(n_895), .Y(n_984) );
NOR2xp33_ASAP7_75t_SL g958 ( .A(n_896), .B(n_959), .Y(n_958) );
NAND3xp33_ASAP7_75t_L g897 ( .A(n_898), .B(n_902), .C(n_908), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
OR2x2_ASAP7_75t_L g916 ( .A(n_900), .B(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g967 ( .A(n_900), .Y(n_967) );
AND2x2_ASAP7_75t_L g972 ( .A(n_900), .B(n_910), .Y(n_972) );
NOR2xp33_ASAP7_75t_L g987 ( .A(n_900), .B(n_922), .Y(n_987) );
OAI221xp5_ASAP7_75t_L g992 ( .A1(n_901), .A2(n_952), .B1(n_993), .B2(n_994), .C(n_995), .Y(n_992) );
AOI21xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B(n_905), .Y(n_902) );
INVx1_ASAP7_75t_L g989 ( .A(n_903), .Y(n_989) );
INVxp67_ASAP7_75t_SL g905 ( .A(n_906), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_911), .B1(n_915), .B2(n_918), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_910), .B(n_957), .Y(n_956) );
A2O1A1Ixp33_ASAP7_75t_L g988 ( .A1(n_910), .A2(n_919), .B(n_989), .C(n_990), .Y(n_988) );
INVx1_ASAP7_75t_L g991 ( .A(n_912), .Y(n_991) );
AOI21xp33_ASAP7_75t_L g947 ( .A1(n_913), .A2(n_948), .B(n_949), .Y(n_947) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_918), .B(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx2_ASAP7_75t_L g929 ( .A(n_922), .Y(n_929) );
AOI221xp5_ASAP7_75t_L g942 ( .A1(n_922), .A2(n_943), .B1(n_945), .B2(n_947), .C(n_951), .Y(n_942) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OAI322xp33_ASAP7_75t_L g951 ( .A1(n_929), .A2(n_941), .A3(n_952), .B1(n_954), .B2(n_956), .C1(n_958), .C2(n_960), .Y(n_951) );
OAI211xp5_ASAP7_75t_L g980 ( .A1(n_929), .A2(n_981), .B(n_982), .C(n_984), .Y(n_980) );
INVx1_ASAP7_75t_L g994 ( .A(n_932), .Y(n_994) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVxp67_ASAP7_75t_SL g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_953), .B(n_969), .Y(n_995) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVxp67_ASAP7_75t_SL g963 ( .A(n_964), .Y(n_963) );
AOI211xp5_ASAP7_75t_SL g985 ( .A1(n_964), .A2(n_986), .B(n_988), .C(n_992), .Y(n_985) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
O2A1O1Ixp33_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .B(n_974), .C(n_980), .Y(n_971) );
INVxp33_ASAP7_75t_SL g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
BUFx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVxp67_ASAP7_75t_SL g998 ( .A(n_999), .Y(n_998) );
XNOR2x2_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1001), .Y(n_999) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_1001), .Y(n_1026) );
NAND3xp33_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1010), .C(n_1013), .Y(n_1001) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1007), .Y(n_1005) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
HB1xp67_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
BUFx2_ASAP7_75t_SL g1022 ( .A(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1026), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
endmodule