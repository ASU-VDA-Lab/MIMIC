module fake_jpeg_1496_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_0),
.B(n_2),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_8),
.B(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_18),
.A2(n_19),
.B1(n_7),
.B2(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_5),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_16),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_10),
.C(n_11),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_26),
.C(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_15),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_30),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_13),
.B1(n_18),
.B2(n_7),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_0),
.B(n_13),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_0),
.Y(n_37)
);


endmodule