module fake_netlist_5_1777_n_2100 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2100);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2100;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1951;
wire n_1825;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_368;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_29),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_73),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_7),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_189),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_148),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_115),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_77),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_125),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_47),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_102),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_39),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_81),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_153),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_107),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_45),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_19),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_134),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_137),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_135),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_109),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_136),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_64),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_196),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_63),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_10),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_127),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_56),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_101),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_7),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_39),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_13),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_61),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_26),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_50),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_9),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_1),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_140),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_113),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_187),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_1),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_123),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_4),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_24),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_75),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_154),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_25),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_192),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_144),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_164),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_71),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_13),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_60),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_89),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_74),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_61),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_149),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_8),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_25),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_117),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_180),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_146),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_171),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_193),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_150),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_108),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_31),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_93),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_106),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_99),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_72),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_63),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_24),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_100),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_188),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_128),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_181),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_139),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_82),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_84),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_178),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_64),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_183),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_10),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_85),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_96),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_97),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_55),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_62),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_6),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_38),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_155),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_71),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_42),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_28),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_95),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_33),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_30),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_62),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_50),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_91),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_132),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_31),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_37),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_75),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_76),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_174),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_2),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_12),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_38),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_34),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_160),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_168),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_141),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_77),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_170),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_65),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_0),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_41),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_161),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_37),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_156),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_182),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_112),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_28),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_118),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_23),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_138),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_58),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_65),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_5),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_116),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_147),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_120),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_70),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_53),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_45),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_11),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_74),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_152),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_176),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_19),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_124),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_16),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_8),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_12),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_0),
.Y(n_356)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_53),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_121),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_88),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_67),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_72),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_51),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_5),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_15),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_83),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_111),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_162),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_119),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_143),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_20),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_167),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_46),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_52),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_103),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_79),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_49),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_33),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_26),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_18),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_36),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_165),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_56),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_51),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_27),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_104),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_29),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_86),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_59),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_131),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_57),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_172),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_133),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_220),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_260),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_357),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_260),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_197),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_197),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_229),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_288),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_223),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_311),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_358),
.B(n_374),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_332),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_202),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_202),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_205),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_260),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_221),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_260),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_358),
.B(n_2),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_198),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_260),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_221),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_287),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_287),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_260),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_200),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_199),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_329),
.B(n_3),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_205),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_209),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_200),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_206),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_387),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_233),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_233),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_201),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_203),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_204),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_206),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_261),
.B(n_3),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_231),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_367),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_237),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_208),
.Y(n_436)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_200),
.B(n_4),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_240),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_376),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_207),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_210),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_L g442 ( 
.A(n_239),
.B(n_6),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_242),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_211),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_207),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_217),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_374),
.B(n_11),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_243),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_244),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_217),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_367),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_245),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_224),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_224),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_232),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_367),
.B(n_14),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_215),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_232),
.B(n_14),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_234),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_222),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_234),
.B(n_15),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_226),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_235),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_376),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_212),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_249),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_250),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_252),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_253),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_255),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_250),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_246),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_257),
.B(n_16),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_239),
.B(n_17),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_239),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_257),
.B(n_17),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_259),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_263),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_251),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_247),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_254),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_256),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_262),
.B(n_18),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_258),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_251),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_271),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_272),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_251),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_280),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_280),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_273),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_262),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_394),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_396),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_401),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_396),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_394),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_401),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_428),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_401),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_413),
.B(n_218),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_408),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_410),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_434),
.B(n_370),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_429),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_423),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_423),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_418),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_409),
.B(n_227),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_399),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_397),
.B(n_218),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_418),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_430),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_436),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_488),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_441),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_444),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_475),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_451),
.B(n_447),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_492),
.B(n_370),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_475),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_400),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_479),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_457),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_403),
.B(n_213),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_460),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_479),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_420),
.B(n_241),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_485),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_439),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_485),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_462),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_488),
.B(n_381),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_489),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_R g542 ( 
.A(n_412),
.B(n_274),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_398),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_402),
.Y(n_544)
);

NOR2x1_ASAP7_75t_L g545 ( 
.A(n_488),
.B(n_218),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_489),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_405),
.B(n_275),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_406),
.B(n_278),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_490),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_466),
.Y(n_550)
);

XNOR2x2_ASAP7_75t_L g551 ( 
.A(n_411),
.B(n_334),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_464),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_407),
.B(n_370),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_421),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_458),
.B(n_223),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_490),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_424),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_456),
.A2(n_268),
.B(n_248),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_412),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_431),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_440),
.B(n_280),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_445),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_461),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_446),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_404),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_450),
.B(n_283),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_453),
.B(n_248),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_454),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_455),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_459),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_419),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_493),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_493),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_493),
.Y(n_575)
);

INVxp67_ASAP7_75t_SL g576 ( 
.A(n_495),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_498),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_503),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_508),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_513),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_561),
.B(n_269),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_508),
.B(n_471),
.Y(n_582)
);

AND2x6_ASAP7_75t_L g583 ( 
.A(n_508),
.B(n_248),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_498),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_513),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_503),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_SL g587 ( 
.A(n_535),
.B(n_414),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_513),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_496),
.Y(n_589)
);

NOR2x1p5_ASAP7_75t_L g590 ( 
.A(n_526),
.B(n_393),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_543),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_496),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_532),
.B(n_465),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_503),
.Y(n_594)
);

OAI21xp33_ASAP7_75t_L g595 ( 
.A1(n_532),
.A2(n_476),
.B(n_473),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_529),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_543),
.Y(n_597)
);

NOR2x1p5_ASAP7_75t_L g598 ( 
.A(n_526),
.B(n_393),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_504),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_542),
.B(n_416),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_496),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_513),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_513),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_496),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_563),
.B(n_425),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_504),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_513),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_527),
.B(n_419),
.Y(n_608)
);

AND2x6_ASAP7_75t_L g609 ( 
.A(n_504),
.B(n_268),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_563),
.B(n_395),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_496),
.Y(n_611)
);

XNOR2x2_ASAP7_75t_L g612 ( 
.A(n_551),
.B(n_334),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_542),
.B(n_395),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_498),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_516),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_527),
.B(n_422),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_504),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_547),
.B(n_422),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_535),
.A2(n_472),
.B1(n_480),
.B2(n_463),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_496),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_550),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_504),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_513),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_547),
.B(n_481),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_561),
.B(n_269),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_510),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_522),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_572),
.B(n_426),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_494),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_537),
.Y(n_630)
);

NOR2x1p5_ASAP7_75t_L g631 ( 
.A(n_500),
.B(n_281),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_496),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_499),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_543),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_561),
.B(n_270),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_554),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_494),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_548),
.B(n_433),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_548),
.B(n_482),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_497),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_499),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_566),
.B(n_484),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_510),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_566),
.B(n_433),
.Y(n_644)
);

OR2x6_ASAP7_75t_L g645 ( 
.A(n_558),
.B(n_268),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_537),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_499),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_497),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_502),
.Y(n_649)
);

INVx4_ASAP7_75t_SL g650 ( 
.A(n_555),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_509),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_499),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_522),
.B(n_435),
.Y(n_653)
);

AND2x6_ASAP7_75t_L g654 ( 
.A(n_518),
.B(n_285),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_555),
.A2(n_483),
.B1(n_442),
.B2(n_474),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_502),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_510),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_505),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_505),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_552),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_527),
.B(n_435),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_550),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_507),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_520),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_507),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_552),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_499),
.Y(n_667)
);

AO21x2_ASAP7_75t_L g668 ( 
.A1(n_558),
.A2(n_277),
.B(n_270),
.Y(n_668)
);

BUFx6f_ASAP7_75t_SL g669 ( 
.A(n_572),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_522),
.B(n_438),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_511),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_522),
.B(n_438),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_522),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_559),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_554),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_555),
.A2(n_437),
.B1(n_336),
.B2(n_356),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_551),
.B(n_427),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_499),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_511),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_557),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_512),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_512),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_555),
.B(n_443),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_499),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_562),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_515),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_555),
.B(n_443),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_562),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_501),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_572),
.B(n_448),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_559),
.B(n_486),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_554),
.B(n_487),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_564),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_564),
.B(n_491),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_556),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_568),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_568),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_557),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_501),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_570),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_555),
.A2(n_281),
.B1(n_330),
.B2(n_336),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_557),
.Y(n_702)
);

AND2x6_ASAP7_75t_L g703 ( 
.A(n_518),
.B(n_285),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_553),
.B(n_277),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_557),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_570),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_515),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_515),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_519),
.Y(n_709)
);

BUFx8_ASAP7_75t_SL g710 ( 
.A(n_517),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_569),
.B(n_448),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_557),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_555),
.B(n_449),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_553),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_569),
.B(n_449),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_501),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_557),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_557),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_560),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_560),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_560),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_553),
.B(n_569),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_551),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_555),
.B(n_452),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_SL g725 ( 
.A(n_521),
.B(n_415),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_595),
.A2(n_579),
.B(n_714),
.C(n_582),
.Y(n_726)
);

NAND2x1p5_ASAP7_75t_L g727 ( 
.A(n_627),
.B(n_558),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_579),
.B(n_555),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_627),
.B(n_572),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_627),
.B(n_673),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_714),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_627),
.B(n_572),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_595),
.A2(n_583),
.B1(n_625),
.B2(n_581),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_722),
.B(n_560),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_599),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_599),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_606),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_610),
.B(n_452),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_722),
.B(n_560),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_606),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_605),
.B(n_468),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_593),
.B(n_560),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_593),
.B(n_560),
.Y(n_743)
);

NOR2x1_ASAP7_75t_L g744 ( 
.A(n_690),
.B(n_216),
.Y(n_744)
);

NAND2x1_ASAP7_75t_L g745 ( 
.A(n_673),
.B(n_495),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_618),
.B(n_468),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_653),
.B(n_571),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_670),
.B(n_571),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_617),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_672),
.B(n_571),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_673),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_617),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_583),
.A2(n_567),
.B1(n_518),
.B2(n_285),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_711),
.B(n_571),
.Y(n_754)
);

XOR2x2_ASAP7_75t_SL g755 ( 
.A(n_612),
.B(n_212),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_582),
.B(n_704),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_723),
.A2(n_432),
.B(n_214),
.C(n_228),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_665),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_622),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_660),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_L g761 ( 
.A(n_619),
.B(n_662),
.Y(n_761)
);

NOR2x1p5_ASAP7_75t_L g762 ( 
.A(n_638),
.B(n_523),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_715),
.B(n_571),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_673),
.B(n_683),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_631),
.B(n_704),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_624),
.A2(n_469),
.B1(n_477),
.B2(n_470),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_576),
.A2(n_501),
.B(n_506),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_622),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_644),
.B(n_571),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_685),
.B(n_571),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_685),
.B(n_518),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_639),
.B(n_469),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_665),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_688),
.B(n_518),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_642),
.B(n_694),
.Y(n_775)
);

AND2x2_ASAP7_75t_SL g776 ( 
.A(n_723),
.B(n_310),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_688),
.B(n_567),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_681),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_693),
.B(n_567),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_660),
.B(n_470),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_693),
.B(n_567),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_SL g782 ( 
.A1(n_615),
.A2(n_516),
.B1(n_517),
.B2(n_266),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_696),
.B(n_567),
.Y(n_783)
);

AND2x6_ASAP7_75t_SL g784 ( 
.A(n_691),
.B(n_214),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_621),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_666),
.B(n_477),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_681),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_687),
.A2(n_330),
.B(n_360),
.C(n_356),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_696),
.B(n_540),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_697),
.B(n_700),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_609),
.Y(n_791)
);

NOR3xp33_ASAP7_75t_L g792 ( 
.A(n_587),
.B(n_478),
.C(n_524),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_697),
.B(n_540),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_583),
.A2(n_478),
.B1(n_213),
.B2(n_225),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_608),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_700),
.B(n_556),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_704),
.B(n_525),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_SL g798 ( 
.A(n_590),
.B(n_598),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_706),
.B(n_556),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_706),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_713),
.B(n_223),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_629),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_666),
.B(n_531),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_629),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_581),
.A2(n_338),
.B(n_219),
.C(n_228),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_637),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_583),
.B(n_223),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_637),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_583),
.B(n_556),
.Y(n_809)
);

HB1xp67_ASAP7_75t_SL g810 ( 
.A(n_651),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_724),
.B(n_223),
.Y(n_811)
);

NOR3xp33_ASAP7_75t_L g812 ( 
.A(n_628),
.B(n_539),
.C(n_533),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_640),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_583),
.B(n_556),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_583),
.B(n_495),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_640),
.B(n_495),
.Y(n_816)
);

O2A1O1Ixp5_ASAP7_75t_L g817 ( 
.A1(n_573),
.A2(n_578),
.B(n_575),
.C(n_574),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_692),
.B(n_544),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_621),
.B(n_565),
.Y(n_819)
);

A2O1A1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_581),
.A2(n_219),
.B(n_236),
.C(n_238),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_674),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_590),
.A2(n_265),
.B1(n_279),
.B2(n_342),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_648),
.Y(n_823)
);

NAND2x1_ASAP7_75t_L g824 ( 
.A(n_609),
.B(n_495),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_581),
.A2(n_236),
.B(n_238),
.C(n_373),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_646),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_650),
.B(n_223),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_625),
.A2(n_310),
.B1(n_292),
.B2(n_294),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_648),
.B(n_506),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_L g830 ( 
.A(n_609),
.B(n_365),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_695),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_608),
.B(n_353),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_616),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_SL g834 ( 
.A(n_598),
.B(n_230),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_591),
.Y(n_835)
);

AND2x6_ASAP7_75t_SL g836 ( 
.A(n_616),
.B(n_300),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_649),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_649),
.B(n_506),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_656),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_661),
.A2(n_631),
.B1(n_704),
.B2(n_635),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_656),
.B(n_514),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_655),
.A2(n_310),
.B1(n_305),
.B2(n_392),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_625),
.A2(n_292),
.B1(n_321),
.B2(n_305),
.Y(n_843)
);

OAI221xp5_ASAP7_75t_L g844 ( 
.A1(n_676),
.A2(n_336),
.B1(n_281),
.B2(n_356),
.C(n_360),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_658),
.B(n_659),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_661),
.A2(n_352),
.B1(n_284),
.B2(n_325),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_658),
.B(n_514),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_659),
.B(n_286),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_663),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_663),
.B(n_286),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_671),
.B(n_294),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_671),
.B(n_321),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_L g853 ( 
.A(n_609),
.B(n_365),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_613),
.B(n_353),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_600),
.B(n_264),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_679),
.B(n_337),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_679),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_682),
.B(n_573),
.Y(n_858)
);

OR2x6_ASAP7_75t_L g859 ( 
.A(n_625),
.B(n_337),
.Y(n_859)
);

NOR2x1p5_ASAP7_75t_L g860 ( 
.A(n_677),
.B(n_664),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_591),
.B(n_267),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_635),
.A2(n_369),
.B1(n_289),
.B2(n_322),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_682),
.B(n_575),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_SL g864 ( 
.A(n_669),
.B(n_304),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_574),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_650),
.B(n_365),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_635),
.A2(n_385),
.B1(n_392),
.B2(n_365),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_635),
.A2(n_385),
.B1(n_365),
.B2(n_360),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_578),
.B(n_525),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_591),
.B(n_530),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_597),
.B(n_530),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_677),
.B(n_300),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_597),
.B(n_634),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_654),
.A2(n_365),
.B1(n_330),
.B2(n_545),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_597),
.A2(n_359),
.B1(n_290),
.B2(n_333),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_R g876 ( 
.A(n_596),
.B(n_295),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_646),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_634),
.B(n_534),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_634),
.B(n_534),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_654),
.A2(n_545),
.B1(n_386),
.B2(n_384),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_586),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_586),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_630),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_636),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_636),
.B(n_536),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_636),
.Y(n_886)
);

AOI221xp5_ASAP7_75t_L g887 ( 
.A1(n_612),
.A2(n_378),
.B1(n_379),
.B2(n_320),
.C(n_324),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_695),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_695),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_675),
.B(n_536),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_675),
.B(n_538),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_594),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_675),
.B(n_538),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_594),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_654),
.A2(n_350),
.B1(n_296),
.B2(n_301),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_669),
.B(n_276),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_654),
.A2(n_703),
.B1(n_609),
.B2(n_701),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_791),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_810),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_756),
.B(n_668),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_735),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_798),
.B(n_725),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_742),
.B(n_654),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_826),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_751),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_743),
.B(n_654),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_751),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_736),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_802),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_756),
.B(n_650),
.Y(n_910)
);

BUFx8_ASAP7_75t_L g911 ( 
.A(n_795),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_835),
.B(n_650),
.Y(n_912)
);

NAND2x1p5_ASAP7_75t_L g913 ( 
.A(n_791),
.B(n_698),
.Y(n_913)
);

AOI21x1_ASAP7_75t_L g914 ( 
.A1(n_801),
.A2(n_717),
.B(n_712),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_731),
.B(n_775),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_R g916 ( 
.A(n_798),
.B(n_669),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_R g917 ( 
.A(n_834),
.B(n_669),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_835),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_877),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_737),
.Y(n_920)
);

INVx3_ASAP7_75t_SL g921 ( 
.A(n_776),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_740),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_749),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_802),
.Y(n_924)
);

NOR3xp33_ASAP7_75t_SL g925 ( 
.A(n_887),
.B(n_291),
.C(n_282),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_876),
.Y(n_926)
);

OAI22xp33_ASAP7_75t_L g927 ( 
.A1(n_840),
.A2(n_645),
.B1(n_362),
.B2(n_328),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_731),
.B(n_654),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_760),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_776),
.A2(n_703),
.B1(n_609),
.B2(n_719),
.Y(n_930)
);

BUFx10_ASAP7_75t_L g931 ( 
.A(n_803),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_752),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_759),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_772),
.B(n_703),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_768),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_813),
.Y(n_936)
);

NOR3xp33_ASAP7_75t_SL g937 ( 
.A(n_834),
.B(n_297),
.C(n_293),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_813),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_797),
.B(n_703),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_823),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_823),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_R g942 ( 
.A(n_864),
.B(n_609),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_797),
.B(n_703),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_751),
.A2(n_680),
.B(n_585),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_795),
.A2(n_703),
.B1(n_720),
.B2(n_719),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_837),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_837),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_746),
.B(n_710),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_857),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_857),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_791),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_832),
.B(n_668),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_758),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_758),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_785),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_800),
.B(n_703),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_773),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_773),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_804),
.B(n_592),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_733),
.B(n_650),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_842),
.A2(n_645),
.B1(n_668),
.B2(n_707),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_806),
.B(n_592),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_SL g963 ( 
.A1(n_782),
.A2(n_345),
.B1(n_298),
.B2(n_302),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_883),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_808),
.B(n_592),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_791),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_778),
.Y(n_967)
);

NAND2x1p5_ASAP7_75t_L g968 ( 
.A(n_791),
.B(n_698),
.Y(n_968)
);

BUFx10_ASAP7_75t_L g969 ( 
.A(n_818),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_833),
.B(n_839),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_778),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_824),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_787),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_R g974 ( 
.A(n_819),
.B(n_316),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_738),
.B(n_299),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_784),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_765),
.B(n_645),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_849),
.B(n_592),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_824),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_787),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_R g981 ( 
.A(n_741),
.B(n_323),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_865),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_821),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_790),
.B(n_611),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_836),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_884),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_765),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_765),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_726),
.B(n_611),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_755),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_780),
.B(n_303),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_786),
.B(n_645),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_865),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_881),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_888),
.Y(n_995)
);

NAND2xp33_ASAP7_75t_SL g996 ( 
.A(n_897),
.B(n_589),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_845),
.B(n_611),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_761),
.A2(n_721),
.B1(n_720),
.B2(n_718),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_SL g999 ( 
.A(n_762),
.B(n_589),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_769),
.B(n_611),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_745),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_789),
.B(n_793),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_745),
.Y(n_1003)
);

NAND2xp33_ASAP7_75t_SL g1004 ( 
.A(n_730),
.B(n_589),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_881),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_882),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_859),
.Y(n_1007)
);

XOR2xp5_ASAP7_75t_L g1008 ( 
.A(n_766),
.B(n_306),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_765),
.B(n_886),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_888),
.Y(n_1010)
);

BUFx10_ASAP7_75t_L g1011 ( 
.A(n_896),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_882),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_892),
.Y(n_1013)
);

BUFx10_ASAP7_75t_L g1014 ( 
.A(n_854),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_755),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_858),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_882),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_892),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_894),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_860),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_859),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_872),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_873),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_815),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_894),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_734),
.B(n_620),
.Y(n_1026)
);

OR2x4_ASAP7_75t_L g1027 ( 
.A(n_872),
.B(n_312),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_859),
.A2(n_645),
.B1(n_686),
.B2(n_707),
.Y(n_1028)
);

INVxp67_ASAP7_75t_SL g1029 ( 
.A(n_730),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_739),
.B(n_620),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_859),
.B(n_686),
.Y(n_1031)
);

AO22x1_ASAP7_75t_L g1032 ( 
.A1(n_855),
.A2(n_363),
.B1(n_307),
.B2(n_390),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_863),
.B(n_620),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_757),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_809),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_889),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_889),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_727),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_817),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_861),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_754),
.B(n_620),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_870),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_763),
.B(n_633),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_871),
.B(n_633),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_757),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_829),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_838),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_822),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_878),
.B(n_633),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_869),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_SL g1051 ( 
.A(n_805),
.B(n_309),
.C(n_308),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_771),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_830),
.B(n_331),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_846),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_744),
.B(n_314),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_727),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_814),
.Y(n_1057)
);

CKINVDCx6p67_ASAP7_75t_R g1058 ( 
.A(n_848),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_879),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_885),
.B(n_633),
.Y(n_1060)
);

BUFx8_ASAP7_75t_L g1061 ( 
.A(n_812),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_727),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_850),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_890),
.B(n_652),
.Y(n_1064)
);

BUFx8_ASAP7_75t_L g1065 ( 
.A(n_792),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_774),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_891),
.B(n_652),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_777),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_893),
.Y(n_1069)
);

NOR3xp33_ASAP7_75t_SL g1070 ( 
.A(n_805),
.B(n_317),
.C(n_315),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_841),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_820),
.B(n_825),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_851),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_728),
.B(n_721),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_830),
.B(n_335),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_794),
.B(n_718),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_847),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_729),
.B(n_732),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_852),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_816),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_779),
.Y(n_1081)
);

AND2x6_ASAP7_75t_SL g1082 ( 
.A(n_856),
.B(n_312),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_875),
.Y(n_1083)
);

HB1xp67_ASAP7_75t_L g1084 ( 
.A(n_820),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_781),
.B(n_717),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_825),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_783),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_753),
.B(n_712),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_729),
.B(n_698),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_853),
.B(n_341),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_SL g1091 ( 
.A(n_862),
.B(n_340),
.C(n_318),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_915),
.B(n_732),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_914),
.A2(n_748),
.B(n_747),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_909),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_921),
.B(n_796),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_929),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1050),
.B(n_843),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_L g1098 ( 
.A(n_975),
.B(n_844),
.C(n_853),
.Y(n_1098)
);

NAND2x1p5_ASAP7_75t_L g1099 ( 
.A(n_1007),
.B(n_827),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1071),
.B(n_828),
.Y(n_1100)
);

INVxp67_ASAP7_75t_SL g1101 ( 
.A(n_905),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_900),
.A2(n_906),
.B(n_903),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_909),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_921),
.A2(n_807),
.B1(n_895),
.B2(n_764),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_987),
.B(n_831),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_900),
.A2(n_811),
.B(n_801),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_SL g1107 ( 
.A1(n_930),
.A2(n_788),
.B(n_799),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1022),
.B(n_1040),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_991),
.B(n_233),
.Y(n_1109)
);

AO22x2_ASAP7_75t_L g1110 ( 
.A1(n_1008),
.A2(n_386),
.B1(n_313),
.B2(n_338),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_987),
.B(n_764),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1078),
.A2(n_811),
.B(n_750),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_924),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_989),
.A2(n_770),
.B(n_767),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1077),
.B(n_868),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_924),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1038),
.A2(n_866),
.B(n_827),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1038),
.A2(n_866),
.B(n_603),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_905),
.A2(n_807),
.B(n_680),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1038),
.A2(n_607),
.B(n_603),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_990),
.A2(n_867),
.B(n_874),
.C(n_880),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1062),
.A2(n_602),
.B(n_607),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1062),
.A2(n_602),
.B(n_652),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_990),
.A2(n_313),
.B(n_348),
.C(n_373),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_936),
.Y(n_1125)
);

BUFx10_ASAP7_75t_L g1126 ( 
.A(n_899),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_952),
.A2(n_348),
.B(n_377),
.C(n_384),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_905),
.A2(n_680),
.B(n_580),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1079),
.B(n_708),
.Y(n_1129)
);

BUFx5_ASAP7_75t_L g1130 ( 
.A(n_1056),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_929),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1062),
.A2(n_684),
.B(n_652),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1016),
.B(n_708),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_904),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1039),
.A2(n_699),
.B(n_684),
.Y(n_1135)
);

AOI21xp33_ASAP7_75t_L g1136 ( 
.A1(n_927),
.A2(n_326),
.B(n_327),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1039),
.A2(n_699),
.B(n_684),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1016),
.B(n_709),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1015),
.B(n_319),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_946),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_944),
.A2(n_699),
.B(n_684),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1063),
.B(n_1073),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1015),
.B(n_339),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1059),
.B(n_709),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_946),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1034),
.A2(n_643),
.A3(n_657),
.B(n_626),
.Y(n_1146)
);

INVxp67_ASAP7_75t_SL g1147 ( 
.A(n_907),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1074),
.A2(n_699),
.B(n_689),
.Y(n_1148)
);

INVx5_ASAP7_75t_L g1149 ( 
.A(n_898),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_SL g1150 ( 
.A(n_1007),
.B(n_343),
.Y(n_1150)
);

INVx5_ASAP7_75t_L g1151 ( 
.A(n_898),
.Y(n_1151)
);

CKINVDCx16_ASAP7_75t_R g1152 ( 
.A(n_1020),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_907),
.A2(n_680),
.B(n_580),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_907),
.A2(n_588),
.B(n_580),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_904),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_952),
.A2(n_377),
.B(n_361),
.C(n_364),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_1034),
.A2(n_643),
.A3(n_626),
.B(n_657),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1029),
.A2(n_705),
.B1(n_702),
.B2(n_678),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_899),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_970),
.B(n_233),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1069),
.B(n_678),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1052),
.B(n_678),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_970),
.B(n_344),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1052),
.B(n_678),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1074),
.A2(n_1030),
.B(n_1026),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1048),
.B(n_346),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1045),
.A2(n_643),
.A3(n_584),
.B(n_577),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1000),
.A2(n_689),
.B(n_584),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_950),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_950),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1057),
.B(n_702),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1066),
.B(n_689),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1066),
.B(n_689),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_981),
.B(n_388),
.C(n_355),
.Y(n_1174)
);

AOI21xp33_ASAP7_75t_L g1175 ( 
.A1(n_1048),
.A2(n_354),
.B(n_351),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_992),
.A2(n_702),
.B1(n_705),
.B2(n_368),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_912),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1041),
.A2(n_577),
.B(n_614),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_931),
.B(n_347),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_961),
.A2(n_577),
.B(n_614),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_992),
.A2(n_705),
.B1(n_391),
.B2(n_389),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1043),
.A2(n_549),
.B(n_528),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1068),
.B(n_549),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_926),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1068),
.B(n_580),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_912),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_995),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1081),
.B(n_585),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1085),
.A2(n_519),
.B(n_528),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1081),
.B(n_585),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_996),
.A2(n_588),
.B(n_585),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_931),
.B(n_372),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1010),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1044),
.A2(n_519),
.B(n_528),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_939),
.A2(n_588),
.B(n_623),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1057),
.B(n_589),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_951),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_943),
.A2(n_588),
.B(n_623),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1036),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1006),
.A2(n_541),
.B(n_546),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1087),
.B(n_1002),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1087),
.B(n_623),
.Y(n_1202)
);

AO21x1_ASAP7_75t_L g1203 ( 
.A1(n_1004),
.A2(n_623),
.B(n_541),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_951),
.Y(n_1204)
);

AOI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1076),
.A2(n_546),
.B(n_541),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1045),
.A2(n_382),
.B(n_380),
.C(n_383),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_938),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_996),
.A2(n_716),
.B(n_667),
.Y(n_1208)
);

BUFx12f_ASAP7_75t_L g1209 ( 
.A(n_1020),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1037),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1046),
.B(n_349),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_911),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1004),
.A2(n_716),
.B(n_667),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1047),
.B(n_366),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_925),
.A2(n_371),
.B(n_546),
.C(n_375),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_931),
.B(n_241),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1042),
.B(n_589),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_926),
.Y(n_1218)
);

AO22x2_ASAP7_75t_L g1219 ( 
.A1(n_1008),
.A2(n_1072),
.B1(n_977),
.B2(n_960),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1042),
.B(n_589),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_901),
.B(n_632),
.Y(n_1221)
);

OR2x6_ASAP7_75t_L g1222 ( 
.A(n_977),
.B(n_632),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1049),
.A2(n_716),
.B(n_667),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_919),
.Y(n_1224)
);

AO21x1_ASAP7_75t_L g1225 ( 
.A1(n_1076),
.A2(n_241),
.B(n_375),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_940),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1006),
.A2(n_716),
.B(n_667),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_908),
.B(n_632),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_920),
.B(n_632),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1006),
.A2(n_716),
.B(n_667),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1014),
.B(n_983),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_960),
.A2(n_716),
.B1(n_667),
.B2(n_632),
.Y(n_1232)
);

INVxp67_ASAP7_75t_SL g1233 ( 
.A(n_898),
.Y(n_1233)
);

O2A1O1Ixp5_ASAP7_75t_L g1234 ( 
.A1(n_934),
.A2(n_241),
.B(n_375),
.C(n_78),
.Y(n_1234)
);

O2A1O1Ixp5_ASAP7_75t_L g1235 ( 
.A1(n_999),
.A2(n_375),
.B(n_80),
.C(n_142),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1061),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1037),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1060),
.A2(n_641),
.B(n_632),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1083),
.A2(n_641),
.B1(n_647),
.B2(n_604),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_922),
.B(n_641),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_988),
.B(n_151),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1064),
.A2(n_641),
.B(n_647),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1055),
.B(n_641),
.C(n_501),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_SL g1244 ( 
.A1(n_966),
.A2(n_186),
.B(n_185),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_923),
.B(n_641),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1014),
.B(n_20),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_964),
.Y(n_1247)
);

NOR2x1_ASAP7_75t_SL g1248 ( 
.A(n_898),
.B(n_951),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_932),
.B(n_21),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_928),
.A2(n_647),
.B(n_604),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1088),
.A2(n_997),
.B(n_984),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_983),
.B(n_21),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1014),
.B(n_22),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1067),
.A2(n_647),
.B(n_604),
.Y(n_1254)
);

NAND2x1p5_ASAP7_75t_L g1255 ( 
.A(n_1007),
.B(n_647),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1177),
.B(n_988),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1120),
.A2(n_962),
.B(n_959),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1103),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1120),
.A2(n_978),
.B(n_965),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1134),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1166),
.A2(n_1054),
.B1(n_948),
.B2(n_969),
.Y(n_1261)
);

BUFx2_ASAP7_75t_SL g1262 ( 
.A(n_1149),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1177),
.Y(n_1263)
);

CKINVDCx16_ASAP7_75t_R g1264 ( 
.A(n_1152),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1219),
.B(n_1086),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1103),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1122),
.A2(n_1033),
.B(n_1037),
.Y(n_1267)
);

AO21x2_ASAP7_75t_L g1268 ( 
.A1(n_1203),
.A2(n_998),
.B(n_1088),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1219),
.B(n_1086),
.Y(n_1269)
);

OR2x6_ASAP7_75t_L g1270 ( 
.A(n_1219),
.B(n_1056),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1098),
.A2(n_999),
.B(n_1054),
.C(n_1091),
.Y(n_1271)
);

AOI222xp33_ASAP7_75t_L g1272 ( 
.A1(n_1110),
.A2(n_1143),
.B1(n_1139),
.B2(n_1166),
.C1(n_963),
.C2(n_1109),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1122),
.A2(n_941),
.B(n_947),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1149),
.Y(n_1274)
);

AO31x2_ASAP7_75t_L g1275 ( 
.A1(n_1127),
.A2(n_949),
.A3(n_1080),
.B(n_958),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1116),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1135),
.A2(n_1025),
.B(n_994),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1112),
.A2(n_956),
.B(n_1089),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1135),
.A2(n_1025),
.B(n_994),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1092),
.A2(n_1028),
.B(n_1084),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1182),
.A2(n_1194),
.B(n_1178),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1187),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1102),
.A2(n_1031),
.B(n_945),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1247),
.Y(n_1284)
);

BUFx2_ASAP7_75t_SL g1285 ( 
.A(n_1149),
.Y(n_1285)
);

BUFx10_ASAP7_75t_L g1286 ( 
.A(n_1184),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1149),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1131),
.B(n_969),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1155),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1247),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1193),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1186),
.B(n_1009),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1209),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1182),
.A2(n_1089),
.B(n_1070),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1127),
.A2(n_967),
.A3(n_980),
.B(n_954),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1116),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1201),
.B(n_1072),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1199),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1096),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1159),
.Y(n_1300)
);

OA21x2_ASAP7_75t_L g1301 ( 
.A1(n_1194),
.A2(n_1013),
.B(n_1005),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_SL g1302 ( 
.A1(n_1244),
.A2(n_986),
.B(n_933),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1125),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1104),
.A2(n_1097),
.B1(n_1105),
.B2(n_1100),
.Y(n_1304)
);

OR2x2_ASAP7_75t_L g1305 ( 
.A(n_1095),
.B(n_935),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1106),
.A2(n_1031),
.B(n_1089),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1125),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1111),
.B(n_977),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1137),
.A2(n_1025),
.B(n_1019),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1145),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1137),
.A2(n_982),
.B(n_1018),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1205),
.A2(n_982),
.B(n_1018),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1142),
.B(n_969),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1136),
.A2(n_1021),
.B1(n_1009),
.B2(n_974),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1159),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1224),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1156),
.A2(n_937),
.B(n_1051),
.C(n_1009),
.Y(n_1317)
);

AOI221xp5_ASAP7_75t_L g1318 ( 
.A1(n_1175),
.A2(n_1032),
.B1(n_976),
.B2(n_902),
.C(n_955),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1207),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1145),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1163),
.B(n_1058),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1178),
.A2(n_993),
.B(n_1019),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1094),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1110),
.A2(n_1061),
.B1(n_942),
.B2(n_976),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1223),
.A2(n_1005),
.B(n_1013),
.Y(n_1325)
);

OAI21xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1115),
.A2(n_986),
.B(n_966),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1251),
.A2(n_973),
.B(n_957),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1121),
.A2(n_973),
.B(n_957),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1186),
.B(n_1160),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1121),
.A2(n_1165),
.B(n_1234),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1139),
.A2(n_1058),
.B1(n_1011),
.B2(n_1057),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1241),
.B(n_918),
.Y(n_1332)
);

BUFx5_ASAP7_75t_L g1333 ( 
.A(n_1111),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1191),
.A2(n_1003),
.B(n_1001),
.Y(n_1334)
);

AOI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1168),
.A2(n_993),
.B(n_971),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1224),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1238),
.A2(n_953),
.B(n_971),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1123),
.A2(n_953),
.B(n_913),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1095),
.B(n_1023),
.Y(n_1339)
);

OAI31xp33_ASAP7_75t_L g1340 ( 
.A1(n_1143),
.A2(n_1072),
.A3(n_918),
.B(n_1027),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_SL g1341 ( 
.A1(n_1107),
.A2(n_966),
.B(n_916),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1210),
.Y(n_1342)
);

AOI21xp33_ASAP7_75t_SL g1343 ( 
.A1(n_1110),
.A2(n_985),
.B(n_1027),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1126),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1113),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1195),
.A2(n_1003),
.B(n_1001),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1141),
.A2(n_968),
.B(n_913),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1210),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1126),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1237),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1236),
.A2(n_985),
.B1(n_1007),
.B2(n_1057),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1105),
.A2(n_1007),
.B1(n_1057),
.B2(n_1035),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1129),
.B(n_1023),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1237),
.Y(n_1354)
);

AO22x2_ASAP7_75t_L g1355 ( 
.A1(n_1111),
.A2(n_1171),
.B1(n_1243),
.B2(n_1226),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1141),
.A2(n_968),
.B(n_1017),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1140),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1254),
.A2(n_1012),
.B(n_1017),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1198),
.A2(n_1003),
.B(n_1001),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1169),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1126),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1170),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1168),
.A2(n_1012),
.B(n_1023),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1144),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1174),
.A2(n_1011),
.B1(n_1035),
.B2(n_1024),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1222),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1211),
.B(n_1023),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1236),
.A2(n_1035),
.B1(n_1024),
.B2(n_1001),
.Y(n_1368)
);

INVx6_ASAP7_75t_L g1369 ( 
.A(n_1151),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1108),
.B(n_1011),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1132),
.A2(n_1001),
.B(n_1003),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1225),
.A2(n_1090),
.B(n_1053),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1231),
.B(n_1179),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1132),
.A2(n_1003),
.B(n_1035),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1105),
.A2(n_1241),
.B1(n_1246),
.B2(n_1253),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1180),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_1184),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1241),
.A2(n_1024),
.B1(n_1061),
.B2(n_1065),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1180),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_SL g1380 ( 
.A1(n_1215),
.A2(n_917),
.B(n_1075),
.C(n_911),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1151),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1183),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1222),
.Y(n_1383)
);

NAND2x1_ASAP7_75t_L g1384 ( 
.A(n_1197),
.B(n_898),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1180),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1222),
.B(n_951),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1156),
.A2(n_1082),
.A3(n_979),
.B(n_972),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1118),
.A2(n_979),
.B(n_972),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1171),
.B(n_910),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1151),
.B(n_979),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1118),
.A2(n_979),
.B(n_972),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1227),
.A2(n_911),
.B(n_1065),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1214),
.B(n_910),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1248),
.A2(n_1065),
.B(n_910),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1133),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1239),
.A2(n_1151),
.B1(n_1231),
.B2(n_1233),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1138),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1206),
.B(n_912),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1162),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1167),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1119),
.A2(n_647),
.B(n_604),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1230),
.A2(n_604),
.B(n_601),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1164),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1197),
.Y(n_1404)
);

OAI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1206),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.C(n_30),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1208),
.A2(n_604),
.B(n_601),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1200),
.A2(n_601),
.B(n_129),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1249),
.B(n_32),
.Y(n_1408)
);

INVx6_ASAP7_75t_L g1409 ( 
.A(n_1130),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1114),
.A2(n_601),
.B(n_130),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1114),
.A2(n_601),
.B(n_126),
.Y(n_1411)
);

CKINVDCx6p67_ASAP7_75t_R g1412 ( 
.A(n_1209),
.Y(n_1412)
);

BUFx2_ASAP7_75t_L g1413 ( 
.A(n_1204),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1204),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1124),
.A2(n_32),
.B(n_34),
.C(n_35),
.Y(n_1415)
);

INVx4_ASAP7_75t_L g1416 ( 
.A(n_1130),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1185),
.A2(n_601),
.B(n_177),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1188),
.A2(n_173),
.B(n_169),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1093),
.A2(n_166),
.B(n_157),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1192),
.B(n_35),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1213),
.A2(n_110),
.B(n_145),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1189),
.A2(n_122),
.B(n_114),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1221),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1189),
.A2(n_94),
.B(n_92),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1289),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1260),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1260),
.Y(n_1427)
);

CKINVDCx14_ASAP7_75t_R g1428 ( 
.A(n_1293),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1297),
.B(n_1216),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1332),
.B(n_1212),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1282),
.Y(n_1431)
);

NAND2xp33_ASAP7_75t_R g1432 ( 
.A(n_1315),
.B(n_1218),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1330),
.A2(n_1093),
.B(n_1196),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1291),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1339),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1297),
.B(n_1124),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1272),
.A2(n_1181),
.B1(n_1252),
.B2(n_1212),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1346),
.A2(n_1196),
.B(n_1190),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1409),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1369),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1298),
.Y(n_1441)
);

NOR2x1_ASAP7_75t_R g1442 ( 
.A(n_1293),
.B(n_1218),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1319),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1405),
.A2(n_1130),
.B1(n_1099),
.B2(n_1117),
.Y(n_1444)
);

NOR2xp67_ASAP7_75t_L g1445 ( 
.A(n_1284),
.B(n_1176),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1316),
.Y(n_1446)
);

AOI21xp33_ASAP7_75t_L g1447 ( 
.A1(n_1304),
.A2(n_1215),
.B(n_1161),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1360),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1323),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1409),
.Y(n_1450)
);

OAI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1261),
.A2(n_1202),
.B1(n_1173),
.B2(n_1172),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1345),
.Y(n_1452)
);

BUFx2_ASAP7_75t_L g1453 ( 
.A(n_1336),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1340),
.A2(n_1150),
.B1(n_1130),
.B2(n_1217),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1332),
.B(n_1101),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1290),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1373),
.A2(n_1130),
.B1(n_1220),
.B2(n_1245),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1375),
.A2(n_1099),
.B1(n_1147),
.B2(n_1228),
.Y(n_1458)
);

NAND2xp33_ASAP7_75t_SL g1459 ( 
.A(n_1315),
.B(n_1229),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1420),
.A2(n_1240),
.B1(n_1158),
.B2(n_1232),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1398),
.A2(n_1130),
.B1(n_1117),
.B2(n_1148),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1382),
.B(n_1157),
.Y(n_1462)
);

OAI211xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1318),
.A2(n_1235),
.B(n_1154),
.C(n_1153),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1377),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1359),
.A2(n_1334),
.B(n_1417),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1321),
.A2(n_1128),
.B1(n_1250),
.B2(n_1255),
.Y(n_1466)
);

INVx5_ASAP7_75t_SL g1467 ( 
.A(n_1412),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1329),
.B(n_1157),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1398),
.A2(n_1242),
.B1(n_1255),
.B2(n_501),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1274),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1410),
.A2(n_1157),
.B(n_1146),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1314),
.A2(n_1242),
.B1(n_1157),
.B2(n_1146),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1332),
.B(n_1146),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1313),
.B(n_1146),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1377),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_SL g1476 ( 
.A1(n_1265),
.A2(n_1242),
.B1(n_40),
.B2(n_41),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1382),
.B(n_1167),
.Y(n_1477)
);

CKINVDCx16_ASAP7_75t_R g1478 ( 
.A(n_1264),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1357),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1265),
.A2(n_36),
.B1(n_40),
.B2(n_42),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1329),
.B(n_1167),
.Y(n_1481)
);

OAI211xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1415),
.A2(n_1408),
.B(n_1324),
.C(n_1271),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1357),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1280),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1274),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1258),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1256),
.B(n_1167),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1269),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1327),
.A2(n_501),
.B(n_90),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1395),
.B(n_48),
.Y(n_1490)
);

NAND2x1_ASAP7_75t_L g1491 ( 
.A(n_1409),
.B(n_87),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1305),
.B(n_48),
.Y(n_1492)
);

OAI222xp33_ASAP7_75t_L g1493 ( 
.A1(n_1270),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.C1(n_55),
.C2(n_57),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1367),
.A2(n_54),
.B(n_58),
.Y(n_1494)
);

NOR2xp67_ASAP7_75t_SL g1495 ( 
.A(n_1262),
.B(n_59),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1308),
.B(n_60),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1256),
.B(n_66),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1331),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1286),
.Y(n_1499)
);

BUFx8_ASAP7_75t_SL g1500 ( 
.A(n_1300),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1286),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1362),
.Y(n_1502)
);

AOI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1343),
.A2(n_1370),
.B1(n_1288),
.B2(n_1317),
.C(n_1364),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1269),
.A2(n_68),
.B1(n_69),
.B2(n_73),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1397),
.B(n_69),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1300),
.Y(n_1506)
);

AOI222xp33_ASAP7_75t_L g1507 ( 
.A1(n_1418),
.A2(n_76),
.B1(n_1393),
.B2(n_1283),
.C1(n_1378),
.C2(n_1364),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1365),
.A2(n_1308),
.B1(n_1305),
.B2(n_1368),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1362),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1270),
.A2(n_1333),
.B1(n_1306),
.B2(n_1355),
.Y(n_1510)
);

AOI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1380),
.A2(n_1351),
.B1(n_1299),
.B2(n_1355),
.C(n_1328),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1308),
.A2(n_1270),
.B1(n_1333),
.B2(n_1339),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1308),
.B(n_1292),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1262),
.B(n_1285),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1256),
.B(n_1292),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1386),
.A2(n_1352),
.B1(n_1361),
.B2(n_1349),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1386),
.A2(n_1361),
.B1(n_1349),
.B2(n_1344),
.Y(n_1517)
);

OAI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1386),
.A2(n_1344),
.B1(n_1383),
.B2(n_1270),
.Y(n_1518)
);

AOI21xp33_ASAP7_75t_L g1519 ( 
.A1(n_1372),
.A2(n_1353),
.B(n_1278),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1371),
.A2(n_1388),
.B(n_1391),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1326),
.A2(n_1396),
.B(n_1423),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_SL g1522 ( 
.A1(n_1384),
.A2(n_1366),
.B(n_1403),
.C(n_1399),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1399),
.A2(n_1403),
.B1(n_1333),
.B2(n_1372),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_L g1524 ( 
.A(n_1292),
.B(n_1389),
.C(n_1366),
.Y(n_1524)
);

INVx6_ASAP7_75t_L g1525 ( 
.A(n_1286),
.Y(n_1525)
);

AOI221xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1383),
.A2(n_1400),
.B1(n_1296),
.B2(n_1404),
.C(n_1413),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1333),
.A2(n_1412),
.B1(n_1389),
.B2(n_1372),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1333),
.A2(n_1389),
.B1(n_1263),
.B2(n_1294),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1263),
.B(n_1333),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1386),
.A2(n_1389),
.B1(n_1355),
.B2(n_1369),
.Y(n_1530)
);

OR2x6_ASAP7_75t_L g1531 ( 
.A(n_1285),
.B(n_1394),
.Y(n_1531)
);

CKINVDCx6p67_ASAP7_75t_R g1532 ( 
.A(n_1414),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1266),
.B(n_1276),
.Y(n_1533)
);

AOI222xp33_ASAP7_75t_L g1534 ( 
.A1(n_1266),
.A2(n_1310),
.B1(n_1276),
.B2(n_1303),
.C1(n_1307),
.C2(n_1320),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1355),
.A2(n_1369),
.B1(n_1263),
.B2(n_1413),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1303),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1394),
.B(n_1341),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1333),
.A2(n_1268),
.B1(n_1278),
.B2(n_1341),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_SL g1539 ( 
.A1(n_1404),
.A2(n_1414),
.B1(n_1369),
.B2(n_1384),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1333),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1275),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1310),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1414),
.B(n_1416),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1320),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1342),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1294),
.A2(n_1278),
.B1(n_1302),
.B2(n_1268),
.Y(n_1546)
);

CKINVDCx16_ASAP7_75t_R g1547 ( 
.A(n_1414),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1348),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1348),
.B(n_1350),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1268),
.A2(n_1294),
.B1(n_1350),
.B2(n_1354),
.Y(n_1550)
);

CKINVDCx9p33_ASAP7_75t_R g1551 ( 
.A(n_1354),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1295),
.Y(n_1552)
);

NAND2xp33_ASAP7_75t_SL g1553 ( 
.A(n_1274),
.B(n_1287),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1387),
.B(n_1275),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1295),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1387),
.B(n_1275),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1414),
.B(n_1416),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1371),
.A2(n_1388),
.B(n_1391),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1302),
.A2(n_1419),
.B1(n_1400),
.B2(n_1376),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1257),
.A2(n_1259),
.B(n_1273),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1416),
.B(n_1392),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1419),
.A2(n_1392),
.B1(n_1421),
.B2(n_1376),
.Y(n_1562)
);

INVx8_ASAP7_75t_L g1563 ( 
.A(n_1274),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1387),
.B(n_1275),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1295),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1274),
.A2(n_1287),
.B1(n_1390),
.B2(n_1379),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1387),
.B(n_1275),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1419),
.A2(n_1421),
.B1(n_1287),
.B2(n_1387),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1379),
.A2(n_1385),
.B1(n_1322),
.B2(n_1301),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1295),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1295),
.B(n_1381),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1287),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1385),
.A2(n_1322),
.B1(n_1301),
.B2(n_1273),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1381),
.A2(n_1424),
.B1(n_1422),
.B2(n_1301),
.Y(n_1574)
);

CKINVDCx6p67_ASAP7_75t_R g1575 ( 
.A(n_1390),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1390),
.A2(n_1381),
.B1(n_1322),
.B2(n_1281),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1311),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1424),
.B(n_1422),
.Y(n_1578)
);

BUFx12f_ASAP7_75t_L g1579 ( 
.A(n_1410),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1411),
.A2(n_1363),
.B1(n_1259),
.B2(n_1257),
.Y(n_1580)
);

CKINVDCx8_ASAP7_75t_R g1581 ( 
.A(n_1281),
.Y(n_1581)
);

OR2x6_ASAP7_75t_L g1582 ( 
.A(n_1347),
.B(n_1374),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1513),
.B(n_1374),
.Y(n_1583)
);

AOI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1484),
.A2(n_1406),
.B1(n_1401),
.B2(n_1335),
.C(n_1312),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1446),
.Y(n_1585)
);

OAI221xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1484),
.A2(n_1504),
.B1(n_1437),
.B2(n_1507),
.C(n_1488),
.Y(n_1586)
);

BUFx12f_ASAP7_75t_L g1587 ( 
.A(n_1501),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1449),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1480),
.A2(n_1312),
.B1(n_1267),
.B2(n_1325),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1494),
.A2(n_1407),
.B1(n_1347),
.B2(n_1356),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1480),
.A2(n_1325),
.B1(n_1337),
.B2(n_1358),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1453),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1488),
.A2(n_1277),
.B1(n_1279),
.B2(n_1309),
.Y(n_1593)
);

AOI221xp5_ASAP7_75t_L g1594 ( 
.A1(n_1493),
.A2(n_1277),
.B1(n_1338),
.B2(n_1402),
.C(n_1482),
.Y(n_1594)
);

OA21x2_ASAP7_75t_L g1595 ( 
.A1(n_1560),
.A2(n_1402),
.B(n_1465),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1498),
.A2(n_1436),
.B1(n_1476),
.B2(n_1429),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1563),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_SL g1598 ( 
.A1(n_1508),
.A2(n_1540),
.B1(n_1539),
.B2(n_1530),
.Y(n_1598)
);

CKINVDCx6p67_ASAP7_75t_R g1599 ( 
.A(n_1478),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1476),
.A2(n_1503),
.B1(n_1495),
.B2(n_1505),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1520),
.A2(n_1558),
.B(n_1465),
.Y(n_1601)
);

BUFx4f_ASAP7_75t_SL g1602 ( 
.A(n_1464),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1503),
.A2(n_1456),
.B1(n_1445),
.B2(n_1425),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1452),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1493),
.A2(n_1456),
.B1(n_1447),
.B2(n_1460),
.C(n_1489),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1490),
.A2(n_1492),
.B1(n_1497),
.B2(n_1511),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1489),
.A2(n_1511),
.B(n_1444),
.C(n_1521),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1435),
.B(n_1515),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1546),
.A2(n_1550),
.B(n_1559),
.Y(n_1609)
);

AO31x2_ASAP7_75t_L g1610 ( 
.A1(n_1576),
.A2(n_1472),
.A3(n_1558),
.B(n_1520),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1470),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1460),
.A2(n_1451),
.B1(n_1519),
.B2(n_1463),
.C(n_1523),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1580),
.A2(n_1438),
.B(n_1574),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1497),
.A2(n_1441),
.B1(n_1434),
.B2(n_1443),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1479),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1550),
.A2(n_1559),
.B(n_1523),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1432),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1431),
.A2(n_1444),
.B1(n_1451),
.B2(n_1459),
.Y(n_1618)
);

OAI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1510),
.A2(n_1527),
.B(n_1526),
.C(n_1568),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1428),
.A2(n_1475),
.B1(n_1506),
.B2(n_1430),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1522),
.A2(n_1438),
.B(n_1566),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1463),
.A2(n_1448),
.B1(n_1430),
.B2(n_1474),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1525),
.A2(n_1524),
.B1(n_1518),
.B2(n_1535),
.Y(n_1623)
);

AOI21xp33_ASAP7_75t_L g1624 ( 
.A1(n_1458),
.A2(n_1457),
.B(n_1454),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1455),
.B(n_1473),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1510),
.A2(n_1525),
.B1(n_1427),
.B2(n_1426),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1455),
.B(n_1547),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1525),
.A2(n_1499),
.B1(n_1468),
.B2(n_1500),
.Y(n_1628)
);

AOI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1554),
.A2(n_1556),
.B1(n_1538),
.B2(n_1541),
.C(n_1564),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1549),
.B(n_1483),
.Y(n_1630)
);

AO21x1_ASAP7_75t_L g1631 ( 
.A1(n_1553),
.A2(n_1516),
.B(n_1566),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1502),
.A2(n_1509),
.B1(n_1481),
.B2(n_1473),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1512),
.A2(n_1572),
.B1(n_1528),
.B2(n_1517),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1467),
.A2(n_1487),
.B1(n_1534),
.B2(n_1462),
.Y(n_1634)
);

OAI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1491),
.A2(n_1514),
.B1(n_1466),
.B2(n_1440),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1532),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1467),
.A2(n_1487),
.B1(n_1477),
.B2(n_1545),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1538),
.A2(n_1467),
.B1(n_1575),
.B2(n_1469),
.Y(n_1638)
);

OAI221xp5_ASAP7_75t_L g1639 ( 
.A1(n_1568),
.A2(n_1461),
.B1(n_1537),
.B2(n_1562),
.C(n_1531),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1548),
.A2(n_1544),
.B1(n_1542),
.B2(n_1536),
.Y(n_1640)
);

OAI211xp5_ASAP7_75t_L g1641 ( 
.A1(n_1541),
.A2(n_1529),
.B(n_1567),
.C(n_1581),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1470),
.Y(n_1642)
);

AOI322xp5_ASAP7_75t_L g1643 ( 
.A1(n_1571),
.A2(n_1565),
.A3(n_1555),
.B1(n_1552),
.B2(n_1570),
.C1(n_1486),
.C2(n_1533),
.Y(n_1643)
);

OAI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1537),
.A2(n_1531),
.B1(n_1514),
.B2(n_1440),
.C(n_1450),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1537),
.A2(n_1531),
.B1(n_1514),
.B2(n_1450),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_SL g1646 ( 
.A1(n_1579),
.A2(n_1563),
.B1(n_1551),
.B2(n_1439),
.Y(n_1646)
);

OR2x6_ASAP7_75t_L g1647 ( 
.A(n_1561),
.B(n_1582),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1470),
.B(n_1485),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1485),
.A2(n_1563),
.B1(n_1551),
.B2(n_1442),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1485),
.A2(n_1582),
.B1(n_1543),
.B2(n_1557),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1433),
.A2(n_1561),
.B1(n_1543),
.B2(n_1557),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1433),
.Y(n_1652)
);

BUFx4f_ASAP7_75t_L g1653 ( 
.A(n_1471),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1471),
.A2(n_1577),
.B1(n_1578),
.B2(n_1569),
.Y(n_1654)
);

AO31x2_ASAP7_75t_L g1655 ( 
.A1(n_1573),
.A2(n_1465),
.A3(n_1576),
.B(n_1472),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1435),
.B(n_1474),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1507),
.B(n_775),
.C(n_772),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1484),
.A2(n_1272),
.B1(n_775),
.B2(n_1015),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1484),
.A2(n_1272),
.B1(n_775),
.B2(n_1015),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1494),
.A2(n_864),
.B1(n_921),
.B2(n_1261),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1484),
.A2(n_775),
.B1(n_595),
.B2(n_563),
.C(n_975),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1464),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1470),
.Y(n_1663)
);

BUFx12f_ASAP7_75t_L g1664 ( 
.A(n_1501),
.Y(n_1664)
);

AOI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1484),
.A2(n_775),
.B1(n_595),
.B2(n_563),
.C(n_975),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1496),
.B(n_1515),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1425),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1429),
.B(n_1297),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1507),
.B(n_775),
.Y(n_1669)
);

OR2x6_ASAP7_75t_L g1670 ( 
.A(n_1537),
.B(n_1270),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1435),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1446),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1470),
.Y(n_1673)
);

AOI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1484),
.A2(n_1272),
.B1(n_775),
.B2(n_1015),
.Y(n_1674)
);

OAI322xp33_ASAP7_75t_L g1675 ( 
.A1(n_1492),
.A2(n_775),
.A3(n_612),
.B1(n_563),
.B2(n_551),
.C1(n_411),
.C2(n_975),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1480),
.A2(n_1015),
.B1(n_1324),
.B2(n_1261),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1437),
.A2(n_775),
.B1(n_921),
.B2(n_1015),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1464),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1484),
.A2(n_1272),
.B1(n_775),
.B2(n_1015),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1507),
.A2(n_775),
.B1(n_818),
.B2(n_772),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1496),
.B(n_1515),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1484),
.A2(n_1272),
.B1(n_775),
.B2(n_1015),
.Y(n_1682)
);

AOI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1507),
.A2(n_775),
.B(n_772),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1484),
.A2(n_775),
.B1(n_595),
.B2(n_563),
.C(n_975),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1429),
.B(n_1297),
.Y(n_1685)
);

AOI221xp5_ASAP7_75t_L g1686 ( 
.A1(n_1484),
.A2(n_775),
.B1(n_595),
.B2(n_563),
.C(n_975),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1435),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_L g1688 ( 
.A(n_1507),
.B(n_775),
.C(n_772),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1429),
.B(n_775),
.Y(n_1689)
);

OAI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1494),
.A2(n_864),
.B1(n_921),
.B2(n_1261),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1496),
.B(n_1515),
.Y(n_1691)
);

NAND3xp33_ASAP7_75t_L g1692 ( 
.A(n_1507),
.B(n_775),
.C(n_772),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1496),
.B(n_1515),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1484),
.A2(n_1272),
.B1(n_775),
.B2(n_1015),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1484),
.A2(n_775),
.B1(n_595),
.B2(n_563),
.C(n_975),
.Y(n_1695)
);

NAND2x1_ASAP7_75t_L g1696 ( 
.A(n_1514),
.B(n_1531),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1484),
.A2(n_1272),
.B1(n_775),
.B2(n_1015),
.Y(n_1697)
);

INVx5_ASAP7_75t_L g1698 ( 
.A(n_1514),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1489),
.A2(n_775),
.B(n_772),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1446),
.Y(n_1700)
);

CKINVDCx14_ASAP7_75t_R g1701 ( 
.A(n_1428),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1437),
.A2(n_775),
.B1(n_921),
.B2(n_1015),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1507),
.A2(n_775),
.B1(n_818),
.B2(n_772),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1489),
.A2(n_775),
.B(n_772),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1437),
.A2(n_775),
.B1(n_921),
.B2(n_1015),
.Y(n_1705)
);

AO31x2_ASAP7_75t_L g1706 ( 
.A1(n_1465),
.A2(n_1576),
.A3(n_1472),
.B(n_1558),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_1470),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1588),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1588),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1585),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1655),
.B(n_1616),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1656),
.B(n_1655),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1655),
.B(n_1616),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1655),
.B(n_1616),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1617),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1604),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1706),
.B(n_1654),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1647),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1706),
.B(n_1654),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1706),
.B(n_1653),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1615),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1609),
.B(n_1647),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1609),
.B(n_1647),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1583),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1610),
.B(n_1652),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1609),
.B(n_1610),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1610),
.B(n_1671),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1610),
.B(n_1687),
.Y(n_1728)
);

NOR2xp67_ASAP7_75t_L g1729 ( 
.A(n_1644),
.B(n_1698),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1683),
.A2(n_1697),
.B1(n_1658),
.B2(n_1694),
.C(n_1659),
.Y(n_1730)
);

NOR4xp25_ASAP7_75t_SL g1731 ( 
.A(n_1669),
.B(n_1586),
.C(n_1605),
.D(n_1607),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1696),
.Y(n_1732)
);

AND2x4_ASAP7_75t_SL g1733 ( 
.A(n_1670),
.B(n_1645),
.Y(n_1733)
);

OAI321xp33_ASAP7_75t_L g1734 ( 
.A1(n_1658),
.A2(n_1674),
.A3(n_1659),
.B1(n_1697),
.B2(n_1682),
.C(n_1694),
.Y(n_1734)
);

INVx3_ASAP7_75t_L g1735 ( 
.A(n_1583),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1674),
.A2(n_1682),
.B1(n_1679),
.B2(n_1680),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1651),
.B(n_1629),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1613),
.B(n_1601),
.Y(n_1738)
);

INVx4_ASAP7_75t_R g1739 ( 
.A(n_1662),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1595),
.B(n_1670),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1670),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1689),
.B(n_1643),
.Y(n_1742)
);

OR2x2_ASAP7_75t_SL g1743 ( 
.A(n_1657),
.B(n_1688),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1592),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1698),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1632),
.B(n_1626),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1698),
.Y(n_1747)
);

NOR2x1_ASAP7_75t_L g1748 ( 
.A(n_1699),
.B(n_1704),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1626),
.B(n_1589),
.Y(n_1749)
);

NOR2xp67_ASAP7_75t_L g1750 ( 
.A(n_1698),
.B(n_1621),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1645),
.B(n_1625),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1630),
.Y(n_1752)
);

AND2x2_ASAP7_75t_SL g1753 ( 
.A(n_1612),
.B(n_1618),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1619),
.B(n_1641),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1589),
.B(n_1607),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1591),
.B(n_1593),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1591),
.B(n_1593),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1631),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1672),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1608),
.Y(n_1760)
);

NAND2x1_ASAP7_75t_L g1761 ( 
.A(n_1618),
.B(n_1640),
.Y(n_1761)
);

INVxp67_ASAP7_75t_SL g1762 ( 
.A(n_1700),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1622),
.B(n_1637),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1650),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1639),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1603),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1622),
.B(n_1637),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1668),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1685),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1640),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1627),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1724),
.B(n_1620),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1708),
.Y(n_1773)
);

AOI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1736),
.A2(n_1675),
.B1(n_1692),
.B2(n_1679),
.C(n_1684),
.Y(n_1774)
);

AOI33xp33_ASAP7_75t_L g1775 ( 
.A1(n_1731),
.A2(n_1600),
.A3(n_1703),
.B1(n_1686),
.B2(n_1665),
.B3(n_1661),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1760),
.B(n_1689),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1708),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1724),
.B(n_1642),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1744),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_L g1780 ( 
.A(n_1748),
.B(n_1695),
.C(n_1669),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1708),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1736),
.A2(n_1676),
.B1(n_1690),
.B2(n_1660),
.Y(n_1782)
);

OAI21x1_ASAP7_75t_L g1783 ( 
.A1(n_1738),
.A2(n_1584),
.B(n_1638),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1744),
.Y(n_1784)
);

INVx3_ASAP7_75t_L g1785 ( 
.A(n_1724),
.Y(n_1785)
);

CKINVDCx12_ASAP7_75t_R g1786 ( 
.A(n_1754),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1724),
.B(n_1666),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1724),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1709),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1735),
.B(n_1598),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1709),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1718),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1709),
.Y(n_1793)
);

OAI211xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1748),
.A2(n_1600),
.B(n_1606),
.C(n_1628),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1735),
.B(n_1623),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1735),
.Y(n_1796)
);

OAI211xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1730),
.A2(n_1606),
.B(n_1628),
.C(n_1614),
.Y(n_1797)
);

NAND3xp33_ASAP7_75t_SL g1798 ( 
.A(n_1731),
.B(n_1705),
.C(n_1677),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_SL g1799 ( 
.A(n_1730),
.B(n_1758),
.C(n_1754),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1732),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1743),
.A2(n_1702),
.B1(n_1596),
.B2(n_1634),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_SL g1802 ( 
.A1(n_1753),
.A2(n_1633),
.B1(n_1701),
.B2(n_1602),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1716),
.Y(n_1803)
);

OAI222xp33_ASAP7_75t_L g1804 ( 
.A1(n_1754),
.A2(n_1596),
.B1(n_1634),
.B2(n_1614),
.C1(n_1649),
.C2(n_1646),
.Y(n_1804)
);

OAI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1734),
.A2(n_1624),
.B1(n_1599),
.B2(n_1635),
.Y(n_1805)
);

AOI21xp33_ASAP7_75t_L g1806 ( 
.A1(n_1753),
.A2(n_1667),
.B(n_1681),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1753),
.B(n_1678),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1721),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1721),
.Y(n_1809)
);

OA332x1_ASAP7_75t_L g1810 ( 
.A1(n_1743),
.A2(n_1602),
.A3(n_1587),
.B1(n_1664),
.B2(n_1691),
.B3(n_1693),
.C1(n_1636),
.C2(n_1594),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1734),
.A2(n_1611),
.B1(n_1673),
.B2(n_1663),
.C(n_1590),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1765),
.A2(n_1597),
.B1(n_1587),
.B2(n_1664),
.Y(n_1812)
);

NOR3xp33_ASAP7_75t_L g1813 ( 
.A(n_1758),
.B(n_1597),
.C(n_1611),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1712),
.B(n_1648),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1715),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1753),
.A2(n_1663),
.B(n_1673),
.Y(n_1816)
);

OAI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1758),
.A2(n_1707),
.B1(n_1765),
.B2(n_1766),
.C(n_1742),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1760),
.B(n_1707),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1735),
.B(n_1707),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1710),
.Y(n_1820)
);

AO21x2_ASAP7_75t_L g1821 ( 
.A1(n_1738),
.A2(n_1707),
.B(n_1726),
.Y(n_1821)
);

OR2x6_ASAP7_75t_L g1822 ( 
.A(n_1729),
.B(n_1750),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1768),
.B(n_1769),
.Y(n_1823)
);

AOI222xp33_ASAP7_75t_L g1824 ( 
.A1(n_1755),
.A2(n_1766),
.B1(n_1742),
.B2(n_1737),
.C1(n_1765),
.C2(n_1746),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1777),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1773),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1800),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1777),
.Y(n_1828)
);

INVx1_ASAP7_75t_SL g1829 ( 
.A(n_1792),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1814),
.B(n_1712),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1821),
.B(n_1732),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1812),
.B(n_1729),
.Y(n_1832)
);

NOR3xp33_ASAP7_75t_L g1833 ( 
.A(n_1780),
.B(n_1765),
.C(n_1743),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1792),
.B(n_1722),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1823),
.B(n_1762),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1785),
.B(n_1722),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1773),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1779),
.B(n_1784),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1781),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1808),
.B(n_1762),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1814),
.B(n_1712),
.Y(n_1841)
);

OAI21x1_ASAP7_75t_SL g1842 ( 
.A1(n_1816),
.A2(n_1732),
.B(n_1745),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1809),
.B(n_1727),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1785),
.B(n_1722),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1785),
.B(n_1723),
.Y(n_1845)
);

NOR2xp33_ASAP7_75t_L g1846 ( 
.A(n_1776),
.B(n_1715),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1820),
.B(n_1768),
.Y(n_1847)
);

CKINVDCx8_ASAP7_75t_R g1848 ( 
.A(n_1815),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1781),
.B(n_1727),
.Y(n_1849)
);

INVx1_ASAP7_75t_SL g1850 ( 
.A(n_1800),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1822),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1803),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1788),
.B(n_1723),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1821),
.B(n_1723),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1803),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1821),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1815),
.B(n_1710),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1789),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1789),
.B(n_1727),
.Y(n_1859)
);

AND2x4_ASAP7_75t_SL g1860 ( 
.A(n_1772),
.B(n_1751),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1791),
.B(n_1728),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1788),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1822),
.B(n_1740),
.Y(n_1863)
);

NOR2x1_ASAP7_75t_L g1864 ( 
.A(n_1822),
.B(n_1750),
.Y(n_1864)
);

OR2x6_ASAP7_75t_L g1865 ( 
.A(n_1822),
.B(n_1741),
.Y(n_1865)
);

NAND2x1p5_ASAP7_75t_L g1866 ( 
.A(n_1783),
.B(n_1747),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1791),
.B(n_1728),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1819),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1793),
.B(n_1768),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1818),
.Y(n_1870)
);

NAND2x1p5_ASAP7_75t_L g1871 ( 
.A(n_1783),
.B(n_1747),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1838),
.Y(n_1872)
);

AOI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1833),
.A2(n_1774),
.B(n_1801),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1838),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1840),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1840),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1870),
.B(n_1847),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1830),
.B(n_1841),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1847),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1826),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1835),
.B(n_1833),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1835),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1843),
.B(n_1759),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1843),
.B(n_1759),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1830),
.B(n_1728),
.Y(n_1885)
);

NOR2x1_ASAP7_75t_SL g1886 ( 
.A(n_1865),
.B(n_1720),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1826),
.Y(n_1887)
);

NAND2xp33_ASAP7_75t_L g1888 ( 
.A(n_1864),
.B(n_1782),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1837),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1868),
.B(n_1752),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1863),
.B(n_1819),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1841),
.B(n_1768),
.Y(n_1892)
);

OAI21xp33_ASAP7_75t_L g1893 ( 
.A1(n_1866),
.A2(n_1799),
.B(n_1782),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1863),
.B(n_1787),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1837),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1868),
.B(n_1752),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1839),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1851),
.B(n_1769),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1863),
.B(n_1787),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1839),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1832),
.A2(n_1798),
.B1(n_1755),
.B2(n_1794),
.Y(n_1901)
);

NAND2x1_ASAP7_75t_L g1902 ( 
.A(n_1864),
.B(n_1739),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1851),
.B(n_1769),
.Y(n_1903)
);

NAND2x1p5_ASAP7_75t_L g1904 ( 
.A(n_1829),
.B(n_1718),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1846),
.B(n_1786),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1827),
.Y(n_1906)
);

AND2x6_ASAP7_75t_SL g1907 ( 
.A(n_1857),
.B(n_1772),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1849),
.B(n_1725),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1849),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1859),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1869),
.B(n_1769),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1863),
.B(n_1787),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1859),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1886),
.B(n_1894),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1881),
.B(n_1824),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1894),
.B(n_1865),
.Y(n_1916)
);

INVx3_ASAP7_75t_SL g1917 ( 
.A(n_1906),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1893),
.B(n_1834),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1873),
.B(n_1848),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1901),
.B(n_1872),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1880),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1880),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1887),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1906),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1874),
.B(n_1834),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1899),
.B(n_1865),
.Y(n_1926)
);

NAND2xp33_ASAP7_75t_SL g1927 ( 
.A(n_1902),
.B(n_1807),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1899),
.B(n_1912),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1912),
.B(n_1865),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1891),
.B(n_1865),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1878),
.B(n_1861),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1889),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1895),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1891),
.B(n_1882),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1897),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1900),
.B(n_1854),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1904),
.B(n_1854),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1904),
.Y(n_1938)
);

AND2x4_ASAP7_75t_SL g1939 ( 
.A(n_1905),
.B(n_1772),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1875),
.B(n_1795),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1908),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1909),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1910),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1888),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1913),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1876),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1890),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1878),
.B(n_1861),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1896),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1883),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1884),
.Y(n_1951)
);

NAND4xp25_ASAP7_75t_L g1952 ( 
.A(n_1905),
.B(n_1775),
.C(n_1802),
.D(n_1817),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1879),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1877),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1885),
.B(n_1867),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1892),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1898),
.B(n_1854),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1908),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1944),
.B(n_1888),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1939),
.B(n_1836),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1939),
.B(n_1836),
.Y(n_1961)
);

NAND2x1p5_ASAP7_75t_L g1962 ( 
.A(n_1914),
.B(n_1829),
.Y(n_1962)
);

OR4x1_ASAP7_75t_L g1963 ( 
.A(n_1921),
.B(n_1827),
.C(n_1862),
.D(n_1770),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1915),
.A2(n_1805),
.B1(n_1848),
.B2(n_1764),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1932),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1927),
.A2(n_1786),
.B1(n_1755),
.B2(n_1797),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1936),
.Y(n_1967)
);

OAI211xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1919),
.A2(n_1806),
.B(n_1903),
.C(n_1811),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1932),
.Y(n_1969)
);

OAI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1920),
.A2(n_1952),
.B(n_1918),
.Y(n_1970)
);

O2A1O1Ixp5_ASAP7_75t_R g1971 ( 
.A1(n_1940),
.A2(n_1911),
.B(n_1907),
.C(n_1869),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1950),
.B(n_1844),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1939),
.B(n_1844),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1950),
.B(n_1845),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1951),
.B(n_1885),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1951),
.B(n_1845),
.Y(n_1976)
);

AOI322xp5_ASAP7_75t_L g1977 ( 
.A1(n_1954),
.A2(n_1737),
.A3(n_1761),
.B1(n_1749),
.B2(n_1856),
.C1(n_1746),
.C2(n_1854),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1925),
.B(n_1866),
.Y(n_1978)
);

OAI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1917),
.A2(n_1764),
.B1(n_1761),
.B2(n_1737),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_SL g1980 ( 
.A1(n_1934),
.A2(n_1764),
.B1(n_1749),
.B2(n_1790),
.Y(n_1980)
);

NAND2x1p5_ASAP7_75t_L g1981 ( 
.A(n_1914),
.B(n_1850),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1934),
.A2(n_1756),
.B1(n_1757),
.B2(n_1749),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1930),
.A2(n_1756),
.B1(n_1757),
.B2(n_1795),
.Y(n_1983)
);

OAI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1946),
.A2(n_1871),
.B(n_1866),
.Y(n_1984)
);

INVxp33_ASAP7_75t_L g1985 ( 
.A(n_1924),
.Y(n_1985)
);

OAI22x1_ASAP7_75t_L g1986 ( 
.A1(n_1917),
.A2(n_1850),
.B1(n_1831),
.B2(n_1871),
.Y(n_1986)
);

XOR2x2_ASAP7_75t_L g1987 ( 
.A(n_1917),
.B(n_1761),
.Y(n_1987)
);

OAI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1946),
.A2(n_1871),
.B(n_1804),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1930),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1928),
.B(n_1853),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1947),
.B(n_1949),
.Y(n_1991)
);

AOI211xp5_ASAP7_75t_L g1992 ( 
.A1(n_1916),
.A2(n_1756),
.B(n_1757),
.C(n_1813),
.Y(n_1992)
);

INVxp67_ASAP7_75t_L g1993 ( 
.A(n_1921),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1947),
.B(n_1853),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1949),
.B(n_1790),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1981),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1965),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1969),
.Y(n_1998)
);

INVxp67_ASAP7_75t_L g1999 ( 
.A(n_1959),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1970),
.B(n_1942),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1993),
.Y(n_2001)
);

O2A1O1Ixp33_ASAP7_75t_L g2002 ( 
.A1(n_1988),
.A2(n_1922),
.B(n_1938),
.C(n_1943),
.Y(n_2002)
);

INVx1_ASAP7_75t_SL g2003 ( 
.A(n_1989),
.Y(n_2003)
);

OAI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1966),
.A2(n_1971),
.B1(n_1980),
.B2(n_1964),
.Y(n_2004)
);

OAI221xp5_ASAP7_75t_L g2005 ( 
.A1(n_1980),
.A2(n_1943),
.B1(n_1945),
.B2(n_1942),
.C(n_1938),
.Y(n_2005)
);

NOR3xp33_ASAP7_75t_L g2006 ( 
.A(n_1979),
.B(n_1922),
.C(n_1945),
.Y(n_2006)
);

BUFx2_ASAP7_75t_L g2007 ( 
.A(n_1981),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1993),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1982),
.A2(n_1928),
.B1(n_1916),
.B2(n_1926),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1983),
.B(n_1928),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1991),
.Y(n_2011)
);

AOI22xp5_ASAP7_75t_L g2012 ( 
.A1(n_1968),
.A2(n_1929),
.B1(n_1926),
.B2(n_1928),
.Y(n_2012)
);

INVxp67_ASAP7_75t_L g2013 ( 
.A(n_1987),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1960),
.B(n_1929),
.Y(n_2014)
);

XNOR2x1_ASAP7_75t_L g2015 ( 
.A(n_1987),
.B(n_1771),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1962),
.Y(n_2016)
);

OAI322xp33_ASAP7_75t_L g2017 ( 
.A1(n_1979),
.A2(n_1995),
.A3(n_1962),
.B1(n_1975),
.B2(n_1974),
.C1(n_1972),
.C2(n_1976),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1985),
.Y(n_2018)
);

INVxp67_ASAP7_75t_L g2019 ( 
.A(n_1967),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1992),
.A2(n_1860),
.B1(n_1937),
.B2(n_1931),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1967),
.Y(n_2021)
);

OAI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_1977),
.A2(n_1953),
.B1(n_1937),
.B2(n_1941),
.C(n_1958),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2021),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_2007),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_2013),
.B(n_1985),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2021),
.Y(n_2026)
);

XNOR2xp5_ASAP7_75t_L g2027 ( 
.A(n_2004),
.B(n_1860),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_2014),
.B(n_1961),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_2003),
.B(n_1973),
.Y(n_2029)
);

NOR3xp33_ASAP7_75t_L g2030 ( 
.A(n_2018),
.B(n_1968),
.C(n_1984),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_2013),
.B(n_1990),
.Y(n_2031)
);

INVxp67_ASAP7_75t_L g2032 ( 
.A(n_2000),
.Y(n_2032)
);

OAI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_2005),
.A2(n_1986),
.B1(n_1963),
.B2(n_1978),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1999),
.B(n_1953),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2001),
.Y(n_2035)
);

NOR3xp33_ASAP7_75t_SL g2036 ( 
.A(n_2017),
.B(n_1994),
.C(n_1956),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1999),
.B(n_1933),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2011),
.B(n_2008),
.Y(n_2038)
);

INVxp67_ASAP7_75t_SL g2039 ( 
.A(n_1996),
.Y(n_2039)
);

NAND4xp25_ASAP7_75t_L g2040 ( 
.A(n_2002),
.B(n_1958),
.C(n_1957),
.D(n_1941),
.Y(n_2040)
);

OAI22xp33_ASAP7_75t_L g2041 ( 
.A1(n_2012),
.A2(n_1931),
.B1(n_1948),
.B2(n_1958),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1997),
.Y(n_2042)
);

XNOR2xp5_ASAP7_75t_L g2043 ( 
.A(n_2027),
.B(n_2015),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2023),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_SL g2045 ( 
.A(n_2039),
.B(n_2016),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_2036),
.A2(n_2006),
.B1(n_2022),
.B2(n_2009),
.C(n_2020),
.Y(n_2046)
);

NAND4xp75_ASAP7_75t_L g2047 ( 
.A(n_2025),
.B(n_2016),
.C(n_2010),
.D(n_1998),
.Y(n_2047)
);

AOI211xp5_ASAP7_75t_L g2048 ( 
.A1(n_2033),
.A2(n_2006),
.B(n_2019),
.C(n_1936),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2032),
.B(n_2026),
.Y(n_2049)
);

AOI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_2033),
.A2(n_2019),
.B(n_1933),
.Y(n_2050)
);

NOR2x1_ASAP7_75t_L g2051 ( 
.A(n_2024),
.B(n_1935),
.Y(n_2051)
);

INVxp67_ASAP7_75t_L g2052 ( 
.A(n_2029),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2035),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2024),
.B(n_1935),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2042),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2051),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2052),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_2046),
.A2(n_2030),
.B1(n_2028),
.B2(n_2041),
.Y(n_2058)
);

O2A1O1Ixp33_ASAP7_75t_L g2059 ( 
.A1(n_2048),
.A2(n_2038),
.B(n_2041),
.C(n_2034),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2045),
.B(n_2031),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_SL g2061 ( 
.A(n_2047),
.B(n_2040),
.C(n_2037),
.Y(n_2061)
);

AND4x2_ASAP7_75t_L g2062 ( 
.A(n_2050),
.B(n_2037),
.C(n_1739),
.D(n_1810),
.Y(n_2062)
);

A2O1A1Ixp33_ASAP7_75t_L g2063 ( 
.A1(n_2049),
.A2(n_1936),
.B(n_1923),
.C(n_1957),
.Y(n_2063)
);

NOR3xp33_ASAP7_75t_L g2064 ( 
.A(n_2049),
.B(n_1956),
.C(n_1923),
.Y(n_2064)
);

OAI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_2054),
.A2(n_1948),
.B1(n_1923),
.B2(n_1955),
.Y(n_2065)
);

OAI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_2043),
.A2(n_1955),
.B1(n_1771),
.B2(n_1741),
.C(n_1745),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_2060),
.B(n_2053),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2056),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_2057),
.B(n_2061),
.Y(n_2069)
);

NAND2xp33_ASAP7_75t_R g2070 ( 
.A(n_2062),
.B(n_2044),
.Y(n_2070)
);

O2A1O1Ixp33_ASAP7_75t_L g2071 ( 
.A1(n_2059),
.A2(n_2055),
.B(n_1842),
.C(n_1936),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2064),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_2068),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_2071),
.A2(n_2058),
.B(n_2069),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2067),
.Y(n_2075)
);

NOR2x1_ASAP7_75t_L g2076 ( 
.A(n_2072),
.B(n_2065),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_2070),
.A2(n_2066),
.B1(n_2063),
.B2(n_1831),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2069),
.B(n_1860),
.Y(n_2078)
);

NOR3xp33_ASAP7_75t_L g2079 ( 
.A(n_2067),
.B(n_1747),
.C(n_1770),
.Y(n_2079)
);

NAND3xp33_ASAP7_75t_SL g2080 ( 
.A(n_2074),
.B(n_1763),
.C(n_1767),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_2073),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_2076),
.A2(n_1831),
.B1(n_1862),
.B2(n_1867),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2075),
.Y(n_2083)
);

OAI221xp5_ASAP7_75t_L g2084 ( 
.A1(n_2077),
.A2(n_1745),
.B1(n_1747),
.B2(n_1741),
.C(n_1771),
.Y(n_2084)
);

AND3x2_ASAP7_75t_L g2085 ( 
.A(n_2078),
.B(n_1831),
.C(n_1718),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2081),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2083),
.B(n_2079),
.Y(n_2087)
);

CKINVDCx20_ASAP7_75t_R g2088 ( 
.A(n_2080),
.Y(n_2088)
);

AOI211xp5_ASAP7_75t_L g2089 ( 
.A1(n_2082),
.A2(n_1767),
.B(n_1763),
.C(n_1746),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2086),
.Y(n_2090)
);

OAI21x1_ASAP7_75t_L g2091 ( 
.A1(n_2090),
.A2(n_2087),
.B(n_2088),
.Y(n_2091)
);

AOI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_2091),
.A2(n_2084),
.B1(n_2089),
.B2(n_2085),
.Y(n_2092)
);

INVxp67_ASAP7_75t_SL g2093 ( 
.A(n_2091),
.Y(n_2093)
);

XNOR2xp5_ASAP7_75t_L g2094 ( 
.A(n_2092),
.B(n_1763),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_2093),
.A2(n_1788),
.B1(n_1796),
.B2(n_1778),
.Y(n_2095)
);

AOI21xp33_ASAP7_75t_L g2096 ( 
.A1(n_2094),
.A2(n_2095),
.B(n_1842),
.Y(n_2096)
);

AOI222xp33_ASAP7_75t_L g2097 ( 
.A1(n_2094),
.A2(n_1767),
.B1(n_1771),
.B2(n_1733),
.C1(n_1858),
.C2(n_1810),
.Y(n_2097)
);

AOI322xp5_ASAP7_75t_L g2098 ( 
.A1(n_2096),
.A2(n_1711),
.A3(n_1714),
.B1(n_1713),
.B2(n_1726),
.C1(n_1719),
.C2(n_1717),
.Y(n_2098)
);

AOI221xp5_ASAP7_75t_L g2099 ( 
.A1(n_2098),
.A2(n_2097),
.B1(n_1858),
.B2(n_1828),
.C(n_1825),
.Y(n_2099)
);

AOI211xp5_ASAP7_75t_L g2100 ( 
.A1(n_2099),
.A2(n_1858),
.B(n_1855),
.C(n_1852),
.Y(n_2100)
);


endmodule