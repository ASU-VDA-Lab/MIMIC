module fake_jpeg_5392_n_321 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_18),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_16),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_65),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

AND2x4_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_18),
.Y(n_63)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_44),
.B(n_27),
.C(n_34),
.D(n_54),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_21),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_73),
.Y(n_86)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_35),
.B1(n_21),
.B2(n_27),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_51),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_21),
.B1(n_27),
.B2(n_34),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_69),
.Y(n_87)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_22),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_74),
.Y(n_99)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_56),
.B(n_69),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_52),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_42),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_54),
.B1(n_39),
.B2(n_41),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_90),
.B1(n_50),
.B2(n_45),
.Y(n_114)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_88),
.B1(n_96),
.B2(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_38),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_41),
.B(n_38),
.C(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_16),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_17),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_100),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_73),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_105),
.C(n_109),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_77),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_22),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_110),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_75),
.B(n_62),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_113),
.Y(n_127)
);

CKINVDCx12_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_114),
.A2(n_50),
.B1(n_47),
.B2(n_34),
.Y(n_140)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_122),
.Y(n_142)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_70),
.B1(n_45),
.B2(n_83),
.Y(n_135)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_66),
.B(n_26),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_79),
.B(n_99),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_99),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_87),
.B1(n_81),
.B2(n_98),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_126),
.B1(n_137),
.B2(n_140),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_128),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_86),
.B1(n_80),
.B2(n_77),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_80),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_86),
.C(n_84),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_138),
.C(n_139),
.Y(n_152)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_79),
.CI(n_96),
.CON(n_130),
.SN(n_130)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_136),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_113),
.B(n_116),
.Y(n_153)
);

AO21x2_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_121),
.B(n_107),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_15),
.B1(n_19),
.B2(n_23),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_41),
.B1(n_50),
.B2(n_45),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_47),
.C(n_36),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_47),
.C(n_36),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_89),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_146),
.C(n_94),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_36),
.C(n_46),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_71),
.B1(n_51),
.B2(n_25),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_26),
.B1(n_17),
.B2(n_22),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_148),
.B(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_117),
.B1(n_115),
.B2(n_100),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_153),
.B(n_170),
.Y(n_181)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_155),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_103),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_157),
.B(n_166),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_158),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_120),
.B(n_92),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_127),
.B1(n_143),
.B2(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_163),
.B1(n_130),
.B2(n_93),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_126),
.C(n_125),
.Y(n_190)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_164),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_65),
.B1(n_94),
.B2(n_33),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_57),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_171),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_94),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_133),
.A2(n_15),
.B(n_14),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_175),
.B1(n_17),
.B2(n_26),
.Y(n_183)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_189),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_128),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_185),
.C(n_190),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_180),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_145),
.Y(n_185)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_159),
.B(n_170),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_195),
.B1(n_177),
.B2(n_188),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_14),
.B(n_28),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_199),
.A2(n_173),
.B(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_14),
.Y(n_200)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_158),
.B1(n_152),
.B2(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_206),
.B(n_207),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_152),
.C(n_161),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_221),
.C(n_187),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_168),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_181),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_201),
.B1(n_176),
.B2(n_179),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_223),
.B1(n_19),
.B2(n_23),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_93),
.B1(n_151),
.B2(n_15),
.Y(n_217)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_194),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_193),
.B(n_197),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_192),
.C(n_181),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_57),
.C(n_29),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_186),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_227),
.C(n_244),
.Y(n_247)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_233),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_216),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_177),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_203),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_199),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_186),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_208),
.A2(n_182),
.B1(n_200),
.B2(n_28),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_11),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_57),
.C(n_76),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_240),
.C(n_241),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_239),
.B(n_243),
.CI(n_219),
.CON(n_249),
.SN(n_249)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_28),
.C(n_25),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_76),
.C(n_72),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_76),
.C(n_48),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_33),
.C(n_30),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_13),
.C(n_12),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_33),
.Y(n_244)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

BUFx12_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_262),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_214),
.B1(n_223),
.B2(n_205),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_248),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_210),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_253),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_2),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_204),
.B1(n_203),
.B2(n_217),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_260),
.B1(n_0),
.B2(n_1),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_225),
.B(n_13),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_225),
.B(n_12),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_258),
.B(n_11),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_241),
.Y(n_273)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_30),
.C(n_1),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_0),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_3),
.Y(n_289)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_255),
.A2(n_229),
.B1(n_243),
.B2(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_278),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_238),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_275),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_254),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_259),
.A2(n_0),
.B(n_2),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_277),
.B(n_263),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_2),
.Y(n_277)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_252),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_249),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_287),
.Y(n_297)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_246),
.B(n_256),
.Y(n_281)
);

OAI21x1_ASAP7_75t_SL g293 ( 
.A1(n_281),
.A2(n_282),
.B(n_275),
.Y(n_293)
);

NOR2xp67_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_247),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_254),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_290),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_256),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_274),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_288),
.B(n_283),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_300),
.B1(n_299),
.B2(n_301),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_266),
.C(n_264),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_295),
.C(n_296),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_269),
.C(n_268),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_3),
.C(n_4),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_4),
.C(n_5),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_302),
.C(n_5),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_283),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_303),
.B(n_10),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_305),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_6),
.C(n_7),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_10),
.B(n_8),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_8),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_310),
.B(n_298),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_8),
.B(n_9),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_311),
.B(n_304),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_312),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_315),
.B(n_9),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_9),
.C(n_10),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_9),
.Y(n_321)
);


endmodule