module fake_jpeg_17920_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx10_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_20),
.A2(n_26),
.B(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_28),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_9),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_15),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_10),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_31),
.B(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_21),
.B(n_17),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_19),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_19),
.B1(n_10),
.B2(n_16),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_6),
.B1(n_9),
.B2(n_31),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_20),
.B1(n_19),
.B2(n_9),
.Y(n_43)
);

AO21x1_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_51),
.B(n_37),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_48),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_22),
.C(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_30),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_50),
.B1(n_46),
.B2(n_47),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_22),
.B1(n_23),
.B2(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_52),
.B(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_58),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_56),
.B1(n_60),
.B2(n_58),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_33),
.B(n_36),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_44),
.C(n_43),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_41),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_45),
.Y(n_62)
);

BUFx24_ASAP7_75t_SL g61 ( 
.A(n_57),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_63),
.C(n_64),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_50),
.B(n_43),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_55),
.C(n_60),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_56),
.B(n_39),
.Y(n_74)
);

AOI31xp67_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_34),
.A3(n_39),
.B(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_34),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_75),
.C(n_34),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_68),
.Y(n_79)
);


endmodule