module real_aes_11753_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_884;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_860;
wire n_748;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_733;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_653;
wire n_155;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
NAND2xp5_ASAP7_75t_L g622 ( .A(n_0), .B(n_200), .Y(n_622) );
INVx1_ASAP7_75t_L g244 ( .A(n_1), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_2), .B(n_194), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_3), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_4), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_5), .B(n_575), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_6), .B(n_150), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_7), .Y(n_618) );
NOR2xp67_ASAP7_75t_L g106 ( .A(n_8), .B(n_91), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_9), .B(n_168), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_10), .B(n_154), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_11), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_12), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_13), .B(n_168), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_14), .B(n_171), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_15), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_16), .B(n_192), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_17), .B(n_168), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_18), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_19), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_20), .B(n_154), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_21), .B(n_150), .Y(n_586) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_22), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_23), .B(n_171), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_24), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_25), .B(n_612), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_26), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_27), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_28), .B(n_171), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_29), .A2(n_104), .B1(n_114), .B2(n_913), .Y(n_103) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_30), .Y(n_152) );
OAI21xp33_ASAP7_75t_L g342 ( .A1(n_31), .A2(n_157), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_32), .B(n_154), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_33), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_34), .B(n_556), .Y(n_555) );
NAND2xp33_ASAP7_75t_SL g545 ( .A(n_35), .B(n_232), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_36), .B(n_154), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_37), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_38), .B(n_175), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_39), .B(n_195), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g108 ( .A(n_40), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g124 ( .A(n_40), .Y(n_124) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_41), .A2(n_72), .B(n_164), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_42), .Y(n_212) );
XOR2xp5_ASAP7_75t_L g135 ( .A(n_43), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_44), .B(n_154), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_45), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_46), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_47), .B(n_175), .Y(n_588) );
AND2x6_ASAP7_75t_L g177 ( .A(n_48), .B(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_49), .B(n_539), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_50), .A2(n_87), .B1(n_194), .B2(n_231), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_51), .B(n_539), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_52), .B(n_192), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_53), .B(n_202), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_54), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_55), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_56), .Y(n_273) );
INVx1_ASAP7_75t_L g178 ( .A(n_57), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_58), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_59), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_60), .B(n_231), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_61), .B(n_231), .Y(n_230) );
NAND2xp33_ASAP7_75t_L g543 ( .A(n_62), .B(n_232), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_63), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_64), .B(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_65), .B(n_175), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_66), .B(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g111 ( .A(n_67), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g254 ( .A(n_68), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_69), .B(n_171), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_70), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_71), .B(n_598), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_73), .B(n_154), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g890 ( .A1(n_74), .A2(n_891), .B(n_899), .Y(n_890) );
INVxp33_ASAP7_75t_SL g901 ( .A(n_74), .Y(n_901) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_75), .B(n_168), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_76), .B(n_192), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_77), .B(n_127), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_77), .Y(n_885) );
INVx1_ASAP7_75t_L g247 ( .A(n_78), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_79), .B(n_175), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_80), .Y(n_173) );
BUFx10_ASAP7_75t_L g131 ( .A(n_81), .Y(n_131) );
INVx1_ASAP7_75t_L g160 ( .A(n_82), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_83), .B(n_168), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_84), .B(n_154), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_85), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_86), .B(n_229), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_88), .B(n_202), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_89), .B(n_168), .Y(n_583) );
INVx1_ASAP7_75t_L g256 ( .A(n_90), .Y(n_256) );
INVx2_ASAP7_75t_L g164 ( .A(n_92), .Y(n_164) );
AOI22x1_ASAP7_75t_SL g893 ( .A1(n_93), .A2(n_95), .B1(n_894), .B2(n_895), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_93), .Y(n_894) );
INVx1_ASAP7_75t_L g113 ( .A(n_94), .Y(n_113) );
OR2x2_ASAP7_75t_L g121 ( .A(n_94), .B(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g528 ( .A(n_94), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_94), .B(n_123), .Y(n_912) );
INVx1_ASAP7_75t_L g895 ( .A(n_95), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_96), .B(n_252), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_97), .B(n_556), .Y(n_643) );
INVx1_ASAP7_75t_L g112 ( .A(n_98), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_99), .B(n_150), .Y(n_610) );
NOR2xp67_ASAP7_75t_L g339 ( .A(n_100), .B(n_340), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_101), .Y(n_573) );
NAND2xp33_ASAP7_75t_L g207 ( .A(n_102), .B(n_202), .Y(n_207) );
INVx3_ASAP7_75t_L g913 ( .A(n_104), .Y(n_913) );
BUFx10_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
AND2x4_ASAP7_75t_L g123 ( .A(n_106), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g110 ( .A(n_111), .B(n_113), .Y(n_110) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_886), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_125), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_117), .A2(n_900), .B(n_904), .Y(n_899) );
NOR2x1p5_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
BUFx12f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_121), .Y(n_898) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x6_ASAP7_75t_L g129 ( .A(n_123), .B(n_130), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_132), .B1(n_133), .B2(n_884), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_127), .B(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g911 ( .A(n_130), .B(n_912), .Y(n_911) );
INVx2_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
BUFx12f_ASAP7_75t_L g889 ( .A(n_131), .Y(n_889) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
XNOR2x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_137), .Y(n_133) );
INVx1_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
OAI22x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_526), .B1(n_529), .B2(n_883), .Y(n_137) );
AND3x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_410), .C(n_483), .Y(n_138) );
NOR2xp67_ASAP7_75t_L g139 ( .A(n_140), .B(n_318), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_299), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_237), .B(n_258), .C(n_284), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_180), .Y(n_142) );
INVx1_ASAP7_75t_L g260 ( .A(n_143), .Y(n_260) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g265 ( .A(n_145), .Y(n_265) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx3_ASAP7_75t_L g303 ( .A(n_146), .Y(n_303) );
INVx1_ASAP7_75t_L g328 ( .A(n_146), .Y(n_328) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_165), .B(n_174), .Y(n_146) );
AO21x1_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_156), .B(n_159), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B1(n_153), .B2(n_155), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g605 ( .A1(n_150), .A2(n_197), .B(n_606), .C(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g598 ( .A(n_151), .Y(n_598) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_152), .Y(n_154) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
INVx2_ASAP7_75t_L g195 ( .A(n_152), .Y(n_195) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_152), .Y(n_232) );
INVx2_ASAP7_75t_L g245 ( .A(n_153), .Y(n_245) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_154), .A2(n_195), .B1(n_617), .B2(n_618), .Y(n_616) );
AOI21x1_ASAP7_75t_L g165 ( .A1(n_156), .A2(n_166), .B(n_169), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_156), .A2(n_250), .B(n_255), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
BUFx2_ASAP7_75t_L g248 ( .A(n_157), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_157), .B(n_279), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_157), .A2(n_339), .B1(n_342), .B2(n_344), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_157), .A2(n_609), .B(n_610), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_157), .A2(n_620), .B(n_621), .Y(n_619) );
BUFx12f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx5_ASAP7_75t_L g197 ( .A(n_158), .Y(n_197) );
INVx5_ASAP7_75t_L g210 ( .A(n_158), .Y(n_210) );
INVxp67_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx3_ASAP7_75t_L g175 ( .A(n_161), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_161), .B(n_256), .Y(n_255) );
AOI21xp33_ASAP7_75t_L g257 ( .A1(n_161), .A2(n_177), .B(n_255), .Y(n_257) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_162), .Y(n_200) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g203 ( .A(n_163), .Y(n_203) );
OR2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx5_ASAP7_75t_L g192 ( .A(n_168), .Y(n_192) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_173), .Y(n_170) );
INVxp67_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_171), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g274 ( .A(n_172), .Y(n_274) );
INVx2_ASAP7_75t_L g556 ( .A(n_172), .Y(n_556) );
INVx2_ASAP7_75t_L g570 ( .A(n_172), .Y(n_570) );
INVx2_ASAP7_75t_L g575 ( .A(n_172), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_179), .Y(n_174) );
INVx8_ASAP7_75t_L g198 ( .A(n_176), .Y(n_198) );
INVx2_ASAP7_75t_SL g297 ( .A(n_176), .Y(n_297) );
INVx8_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g220 ( .A(n_177), .Y(n_220) );
INVx1_ASAP7_75t_L g277 ( .A(n_177), .Y(n_277) );
OAI21x1_ASAP7_75t_L g581 ( .A1(n_177), .A2(n_582), .B(n_585), .Y(n_581) );
OAI21x1_ASAP7_75t_SL g604 ( .A1(n_177), .A2(n_605), .B(n_608), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g615 ( .A1(n_177), .A2(n_296), .B(n_616), .C(n_619), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_180), .A2(n_496), .B1(n_498), .B2(n_500), .Y(n_495) );
AND2x4_ASAP7_75t_L g180 ( .A(n_181), .B(n_204), .Y(n_180) );
AND2x4_ASAP7_75t_L g369 ( .A(n_181), .B(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x4_ASAP7_75t_L g261 ( .A(n_182), .B(n_221), .Y(n_261) );
INVx2_ASAP7_75t_L g385 ( .A(n_182), .Y(n_385) );
AND2x2_ASAP7_75t_L g404 ( .A(n_182), .B(n_317), .Y(n_404) );
AND2x2_ASAP7_75t_L g420 ( .A(n_182), .B(n_205), .Y(n_420) );
AND2x2_ASAP7_75t_L g516 ( .A(n_182), .B(n_328), .Y(n_516) );
BUFx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g307 ( .A(n_183), .Y(n_307) );
OAI21x1_ASAP7_75t_SL g183 ( .A1(n_184), .A2(n_199), .B(n_201), .Y(n_183) );
OAI21x1_ASAP7_75t_SL g184 ( .A1(n_185), .A2(n_190), .B(n_198), .Y(n_184) );
AOI21x1_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_189), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .B(n_196), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_192), .A2(n_194), .B1(n_212), .B2(n_213), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_192), .A2(n_251), .B1(n_253), .B2(n_254), .Y(n_250) );
OAI22xp33_ASAP7_75t_L g272 ( .A1(n_194), .A2(n_273), .B1(n_274), .B2(n_275), .Y(n_272) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g229 ( .A(n_195), .Y(n_229) );
INVx1_ASAP7_75t_L g281 ( .A(n_195), .Y(n_281) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_197), .A2(n_234), .B(n_235), .Y(n_233) );
OAI21xp33_ASAP7_75t_L g271 ( .A1(n_197), .A2(n_272), .B(n_276), .Y(n_271) );
O2A1O1Ixp5_ASAP7_75t_L g572 ( .A1(n_197), .A2(n_573), .B(n_574), .C(n_576), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_197), .A2(n_583), .B(n_584), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_197), .A2(n_645), .B(n_646), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_198), .A2(n_227), .B(n_233), .Y(n_226) );
AO31x2_ASAP7_75t_L g336 ( .A1(n_198), .A2(n_337), .A3(n_338), .B(n_345), .Y(n_336) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_198), .A2(n_554), .B(n_558), .Y(n_553) );
OAI21x1_ASAP7_75t_L g640 ( .A1(n_198), .A2(n_641), .B(n_644), .Y(n_640) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_199), .A2(n_289), .B(n_298), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_199), .A2(n_590), .B(n_599), .Y(n_589) );
OAI21x1_ASAP7_75t_L g634 ( .A1(n_199), .A2(n_590), .B(n_599), .Y(n_634) );
BUFx4f_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g225 ( .A(n_200), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_200), .B(n_277), .Y(n_276) );
OAI21x1_ASAP7_75t_L g603 ( .A1(n_200), .A2(n_604), .B(n_611), .Y(n_603) );
NOR2x1p5_ASAP7_75t_SL g219 ( .A(n_202), .B(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g337 ( .A(n_202), .Y(n_337) );
OAI21x1_ASAP7_75t_L g552 ( .A1(n_202), .A2(n_553), .B(n_561), .Y(n_552) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_202), .A2(n_567), .B(n_577), .Y(n_566) );
OA21x2_ASAP7_75t_L g614 ( .A1(n_202), .A2(n_615), .B(n_622), .Y(n_614) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_202), .A2(n_640), .B(n_647), .Y(n_639) );
BUFx5_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g347 ( .A(n_203), .Y(n_347) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_203), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_204), .B(n_327), .Y(n_455) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_221), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_205), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g332 ( .A(n_205), .Y(n_332) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g306 ( .A(n_206), .Y(n_306) );
HB1xp67_ASAP7_75t_SL g330 ( .A(n_206), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_206), .B(n_328), .Y(n_359) );
AND2x2_ASAP7_75t_L g374 ( .A(n_206), .B(n_307), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_206), .B(n_317), .Y(n_375) );
INVx1_ASAP7_75t_L g403 ( .A(n_206), .Y(n_403) );
AND2x2_ASAP7_75t_L g426 ( .A(n_206), .B(n_265), .Y(n_426) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_211), .B(n_214), .C(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_209), .A2(n_228), .B(n_230), .Y(n_227) );
CKINVDCx6p67_ASAP7_75t_R g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_SL g218 ( .A(n_210), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_210), .A2(n_291), .B(n_292), .Y(n_290) );
INVx2_ASAP7_75t_SL g296 ( .A(n_210), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g541 ( .A1(n_210), .A2(n_281), .B(n_542), .C(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_210), .A2(n_555), .B(n_557), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_210), .A2(n_592), .B(n_593), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_217), .C(n_218), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_218), .A2(n_569), .B(n_571), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_218), .A2(n_586), .B(n_587), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_218), .A2(n_642), .B(n_643), .Y(n_641) );
BUFx2_ASAP7_75t_L g263 ( .A(n_221), .Y(n_263) );
AND2x4_ASAP7_75t_L g384 ( .A(n_221), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g419 ( .A(n_221), .Y(n_419) );
INVx3_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x4_ASAP7_75t_L g370 ( .A(n_222), .B(n_303), .Y(n_370) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g317 ( .A(n_223), .Y(n_317) );
OAI21x1_ASAP7_75t_SL g223 ( .A1(n_224), .A2(n_226), .B(n_236), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g252 ( .A(n_232), .Y(n_252) );
INVx2_ASAP7_75t_L g341 ( .A(n_232), .Y(n_341) );
INVx2_ASAP7_75t_L g343 ( .A(n_232), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_237), .B(n_335), .Y(n_501) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g421 ( .A(n_238), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_238), .B(n_409), .Y(n_497) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_239), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g467 ( .A(n_239), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_239), .B(n_468), .Y(n_494) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g309 ( .A(n_240), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g433 ( .A(n_240), .B(n_302), .Y(n_433) );
AND2x2_ASAP7_75t_L g442 ( .A(n_240), .B(n_366), .Y(n_442) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g269 ( .A(n_241), .Y(n_269) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_249), .B(n_257), .Y(n_241) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_246), .B(n_248), .Y(n_242) );
NOR2x1_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI21xp33_ASAP7_75t_SL g258 ( .A1(n_259), .A2(n_262), .B(n_266), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g323 ( .A1(n_261), .A2(n_324), .B(n_329), .C(n_331), .Y(n_323) );
AND2x2_ASAP7_75t_L g425 ( .A(n_261), .B(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_261), .B(n_330), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_261), .B(n_479), .Y(n_478) );
OAI222xp33_ASAP7_75t_L g520 ( .A1(n_262), .A2(n_321), .B1(n_438), .B2(n_521), .C1(n_522), .C2(n_525), .Y(n_520) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x4_ASAP7_75t_L g304 ( .A(n_263), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g331 ( .A(n_263), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g463 ( .A(n_263), .Y(n_463) );
INVx2_ASAP7_75t_L g313 ( .A(n_265), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_266), .A2(n_449), .B(n_451), .C(n_454), .Y(n_448) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_267), .A2(n_300), .B1(n_308), .B2(n_311), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_267), .A2(n_459), .B1(n_460), .B2(n_461), .Y(n_458) );
AND2x2_ASAP7_75t_L g504 ( .A(n_267), .B(n_335), .Y(n_504) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g439 ( .A(n_268), .B(n_409), .Y(n_439) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
OR2x2_ASAP7_75t_L g349 ( .A(n_269), .B(n_270), .Y(n_349) );
INVx2_ASAP7_75t_L g355 ( .A(n_269), .Y(n_355) );
INVx2_ASAP7_75t_SL g310 ( .A(n_270), .Y(n_310) );
AND2x2_ASAP7_75t_L g354 ( .A(n_270), .B(n_355), .Y(n_354) );
AND2x4_ASAP7_75t_L g394 ( .A(n_270), .B(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_270), .Y(n_407) );
INVx1_ASAP7_75t_L g423 ( .A(n_270), .Y(n_423) );
OA21x2_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_278), .B(n_283), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_274), .A2(n_280), .B1(n_281), .B2(n_282), .Y(n_279) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g308 ( .A(n_286), .B(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g353 ( .A(n_286), .Y(n_353) );
OR2x2_ASAP7_75t_L g444 ( .A(n_286), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_286), .B(n_392), .Y(n_519) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g335 ( .A(n_287), .B(n_336), .Y(n_335) );
AND2x4_ASAP7_75t_L g428 ( .A(n_287), .B(n_380), .Y(n_428) );
BUFx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g366 ( .A(n_288), .Y(n_366) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_293), .B(n_297), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B(n_296), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_296), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_296), .A2(n_559), .B(n_560), .Y(n_558) );
AOI21x1_ASAP7_75t_L g594 ( .A1(n_296), .A2(n_595), .B(n_596), .Y(n_594) );
OAI21x1_ASAP7_75t_L g540 ( .A1(n_297), .A2(n_541), .B(n_544), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_297), .A2(n_568), .B(n_572), .Y(n_567) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_297), .A2(n_591), .B(n_594), .Y(n_590) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
AND2x2_ASAP7_75t_L g322 ( .A(n_301), .B(n_305), .Y(n_322) );
OR2x2_ASAP7_75t_L g417 ( .A(n_301), .B(n_373), .Y(n_417) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_301), .Y(n_491) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_304), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g511 ( .A(n_304), .B(n_512), .Y(n_511) );
AND2x4_ASAP7_75t_L g314 ( .A(n_305), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g432 ( .A(n_305), .B(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g437 ( .A(n_305), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_305), .B(n_370), .Y(n_499) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g326 ( .A(n_307), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_307), .B(n_317), .Y(n_398) );
INVx2_ASAP7_75t_L g388 ( .A(n_309), .Y(n_388) );
AND2x4_ASAP7_75t_SL g427 ( .A(n_309), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g474 ( .A(n_309), .B(n_353), .Y(n_474) );
AND2x2_ASAP7_75t_L g378 ( .A(n_310), .B(n_366), .Y(n_378) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
OR2x2_ASAP7_75t_L g382 ( .A(n_313), .B(n_375), .Y(n_382) );
INVx2_ASAP7_75t_L g391 ( .A(n_313), .Y(n_391) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g357 ( .A(n_316), .B(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g472 ( .A(n_316), .B(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g477 ( .A(n_316), .B(n_402), .Y(n_477) );
AND2x2_ASAP7_75t_L g482 ( .A(n_316), .B(n_374), .Y(n_482) );
AND2x2_ASAP7_75t_L g503 ( .A(n_316), .B(n_426), .Y(n_503) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND3xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_356), .C(n_389), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_350), .Y(n_319) );
AOI21xp33_ASAP7_75t_SL g320 ( .A1(n_321), .A2(n_323), .B(n_333), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
BUFx2_ASAP7_75t_L g471 ( .A(n_326), .Y(n_471) );
INVx1_ASAP7_75t_L g372 ( .A(n_327), .Y(n_372) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g402 ( .A(n_328), .B(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_332), .B(n_404), .Y(n_431) );
AND2x4_ASAP7_75t_SL g515 ( .A(n_332), .B(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_334), .A2(n_390), .B1(n_392), .B2(n_396), .C(n_399), .Y(n_389) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_348), .Y(n_334) );
INVx2_ASAP7_75t_L g387 ( .A(n_335), .Y(n_387) );
INVx1_ASAP7_75t_L g450 ( .A(n_335), .Y(n_450) );
AND2x2_ASAP7_75t_L g481 ( .A(n_335), .B(n_354), .Y(n_481) );
INVx1_ASAP7_75t_L g364 ( .A(n_336), .Y(n_364) );
INVx2_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
INVx2_ASAP7_75t_SL g395 ( .A(n_336), .Y(n_395) );
AND2x2_ASAP7_75t_L g409 ( .A(n_336), .B(n_366), .Y(n_409) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx2_ASAP7_75t_SL g539 ( .A(n_347), .Y(n_539) );
INVx1_ASAP7_75t_L g612 ( .A(n_347), .Y(n_612) );
AND2x2_ASAP7_75t_L g429 ( .A(n_348), .B(n_362), .Y(n_429) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g453 ( .A(n_349), .Y(n_453) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g525 ( .A(n_352), .Y(n_525) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AND2x2_ASAP7_75t_L g512 ( .A(n_353), .B(n_422), .Y(n_512) );
AND2x4_ASAP7_75t_L g379 ( .A(n_355), .B(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_355), .Y(n_393) );
AOI211xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_360), .B(n_367), .C(n_381), .Y(n_356) );
INVx1_ASAP7_75t_L g412 ( .A(n_357), .Y(n_412) );
AND2x2_ASAP7_75t_L g396 ( .A(n_358), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g464 ( .A(n_359), .Y(n_464) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_363), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g457 ( .A(n_363), .Y(n_457) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g422 ( .A(n_364), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g489 ( .A(n_366), .Y(n_489) );
AOI31xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .A3(n_375), .B(n_376), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_369), .A2(n_441), .B1(n_443), .B2(n_446), .Y(n_440) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x4_ASAP7_75t_L g466 ( .A(n_378), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_378), .B(n_494), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_386), .Y(n_381) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_382), .A2(n_400), .B(n_405), .Y(n_399) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g390 ( .A(n_384), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g414 ( .A(n_386), .Y(n_414) );
OR2x6_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVxp67_ASAP7_75t_L g434 ( .A(n_387), .Y(n_434) );
OR2x6_ASAP7_75t_L g507 ( .A(n_391), .B(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g524 ( .A(n_393), .Y(n_524) );
AND2x2_ASAP7_75t_L g441 ( .A(n_394), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g445 ( .A(n_394), .Y(n_445) );
AND2x2_ASAP7_75t_L g523 ( .A(n_394), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g468 ( .A(n_395), .Y(n_468) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_404), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g473 ( .A(n_402), .Y(n_473) );
AND2x2_ASAP7_75t_L g460 ( .A(n_404), .B(n_426), .Y(n_460) );
OR2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_435), .C(n_456), .Y(n_410) );
OAI211xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_413), .B(n_415), .C(n_424), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B(n_421), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_418), .A2(n_486), .B1(n_490), .B2(n_492), .Y(n_485) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx2_ASAP7_75t_L g508 ( .A(n_420), .Y(n_508) );
AOI222xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_427), .B1(n_429), .B2(n_430), .C1(n_432), .C2(n_434), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_426), .A2(n_470), .B(n_472), .Y(n_469) );
INVx2_ASAP7_75t_L g479 ( .A(n_426), .Y(n_479) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI211xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B(n_440), .C(n_448), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_437), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g506 ( .A(n_441), .Y(n_506) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_444), .B(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g487 ( .A(n_445), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_452), .A2(n_479), .B1(n_506), .B2(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g459 ( .A(n_453), .Y(n_459) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_458), .B(n_465), .C(n_480), .Y(n_456) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_469), .B1(n_474), .B2(n_475), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_466), .A2(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_509), .C(n_520), .Y(n_483) );
NAND3xp33_ASAP7_75t_SL g484 ( .A(n_485), .B(n_495), .C(n_502), .Y(n_484) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVxp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AOI21xp33_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_504), .B(n_505), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_517), .Y(n_509) );
NOR2xp67_ASAP7_75t_L g510 ( .A(n_511), .B(n_513), .Y(n_510) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g521 ( .A(n_516), .Y(n_521) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
BUFx8_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
BUFx8_ASAP7_75t_L g883 ( .A(n_528), .Y(n_883) );
XOR2x1_ASAP7_75t_L g892 ( .A(n_529), .B(n_893), .Y(n_892) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_762), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_692), .C(n_733), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_532), .B(n_675), .Y(n_531) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_578), .B1(n_623), .B2(n_626), .C(n_659), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_548), .Y(n_534) );
INVx1_ASAP7_75t_L g674 ( .A(n_535), .Y(n_674) );
INVx1_ASAP7_75t_L g688 ( .A(n_535), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_535), .B(n_662), .Y(n_761) );
INVx1_ASAP7_75t_L g813 ( .A(n_535), .Y(n_813) );
AND2x2_ASAP7_75t_L g862 ( .A(n_535), .B(n_752), .Y(n_862) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g664 ( .A(n_536), .B(n_625), .Y(n_664) );
AND2x2_ASAP7_75t_L g855 ( .A(n_536), .B(n_803), .Y(n_855) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_537), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_537), .B(n_625), .Y(n_739) );
INVx2_ASAP7_75t_L g768 ( .A(n_537), .Y(n_768) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g653 ( .A(n_538), .B(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_538), .Y(n_832) );
OAI21x1_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B(n_547), .Y(n_538) );
OAI21x1_ASAP7_75t_L g580 ( .A1(n_539), .A2(n_581), .B(n_588), .Y(n_580) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_549), .B(n_653), .Y(n_699) );
INVx1_ASAP7_75t_L g723 ( .A(n_549), .Y(n_723) );
INVxp67_ASAP7_75t_SL g772 ( .A(n_549), .Y(n_772) );
NAND2x1_ASAP7_75t_L g814 ( .A(n_549), .B(n_751), .Y(n_814) );
AND2x2_ASAP7_75t_L g859 ( .A(n_549), .B(n_801), .Y(n_859) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_563), .Y(n_549) );
INVx3_ASAP7_75t_L g760 ( .A(n_550), .Y(n_760) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g685 ( .A(n_551), .Y(n_685) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g625 ( .A(n_552), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_563), .B(n_703), .Y(n_781) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_564), .B(n_685), .Y(n_769) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g672 ( .A(n_565), .Y(n_672) );
AND2x2_ASAP7_75t_L g729 ( .A(n_565), .B(n_638), .Y(n_729) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g663 ( .A(n_566), .Y(n_663) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_600), .Y(n_578) );
INVx2_ASAP7_75t_L g665 ( .A(n_579), .Y(n_665) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_579), .Y(n_716) );
AND2x2_ASAP7_75t_L g741 ( .A(n_579), .B(n_681), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_579), .B(n_756), .Y(n_835) );
AND2x2_ASAP7_75t_L g838 ( .A(n_579), .B(n_790), .Y(n_838) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_589), .Y(n_579) );
INVx2_ASAP7_75t_L g631 ( .A(n_580), .Y(n_631) );
BUFx2_ASAP7_75t_L g678 ( .A(n_589), .Y(n_678) );
AND2x2_ASAP7_75t_L g697 ( .A(n_589), .B(n_631), .Y(n_697) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx2_ASAP7_75t_L g666 ( .A(n_600), .Y(n_666) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_601), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_613), .Y(n_601) );
INVx1_ASAP7_75t_L g630 ( .A(n_602), .Y(n_630) );
INVx2_ASAP7_75t_SL g658 ( .A(n_602), .Y(n_658) );
AND2x2_ASAP7_75t_L g719 ( .A(n_602), .B(n_631), .Y(n_719) );
AND2x2_ASAP7_75t_L g790 ( .A(n_602), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g819 ( .A(n_602), .Y(n_819) );
INVxp67_ASAP7_75t_SL g842 ( .A(n_602), .Y(n_842) );
INVx3_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g706 ( .A(n_603), .B(n_614), .Y(n_706) );
AND2x2_ASAP7_75t_L g632 ( .A(n_613), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g681 ( .A(n_613), .B(n_658), .Y(n_681) );
AND2x2_ASAP7_75t_L g713 ( .A(n_613), .B(n_685), .Y(n_713) );
INVx1_ASAP7_75t_L g791 ( .A(n_613), .Y(n_791) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g669 ( .A(n_614), .B(n_633), .Y(n_669) );
INVx2_ASAP7_75t_L g732 ( .A(n_614), .Y(n_732) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g753 ( .A(n_624), .B(n_663), .Y(n_753) );
INVx2_ASAP7_75t_L g877 ( .A(n_624), .Y(n_877) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_635), .B1(n_648), .B2(n_652), .C(n_655), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g874 ( .A1(n_627), .A2(n_872), .B1(n_875), .B2(n_878), .C(n_880), .Y(n_874) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x4_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
NOR2xp67_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_630), .Y(n_807) );
AND2x2_ASAP7_75t_L g657 ( .A(n_631), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g709 ( .A(n_631), .Y(n_709) );
INVx1_ASAP7_75t_L g798 ( .A(n_631), .Y(n_798) );
INVx1_ASAP7_75t_L g817 ( .A(n_631), .Y(n_817) );
AND2x2_ASAP7_75t_L g656 ( .A(n_632), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g721 ( .A(n_632), .Y(n_721) );
INVx2_ASAP7_75t_SL g651 ( .A(n_633), .Y(n_651) );
AND2x4_ASAP7_75t_L g797 ( .A(n_633), .B(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVxp67_ASAP7_75t_R g749 ( .A(n_634), .Y(n_749) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g880 ( .A1(n_636), .A2(n_723), .B(n_840), .C(n_881), .Y(n_880) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g831 ( .A(n_637), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g654 ( .A(n_638), .Y(n_654) );
AND2x2_ASAP7_75t_L g687 ( .A(n_638), .B(n_672), .Y(n_687) );
INVx1_ASAP7_75t_L g703 ( .A(n_638), .Y(n_703) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_SL g757 ( .A(n_648), .Y(n_757) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_L g784 ( .A(n_651), .B(n_719), .Y(n_784) );
NAND4xp25_ASAP7_75t_SL g810 ( .A(n_652), .B(n_788), .C(n_811), .D(n_814), .Y(n_810) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_653), .B(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_653), .B(n_671), .Y(n_867) );
INVx1_ASAP7_75t_L g803 ( .A(n_654), .Y(n_803) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g668 ( .A(n_657), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g731 ( .A(n_657), .B(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g745 ( .A(n_657), .B(n_746), .Y(n_745) );
OAI32xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_665), .A3(n_666), .B1(n_667), .B2(n_670), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OA21x2_ASAP7_75t_L g700 ( .A1(n_661), .A2(n_701), .B(n_704), .Y(n_700) );
AND2x4_ASAP7_75t_SL g661 ( .A(n_662), .B(n_664), .Y(n_661) );
AND2x2_ASAP7_75t_L g812 ( .A(n_662), .B(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g776 ( .A(n_664), .B(n_702), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_666), .A2(n_676), .B1(n_682), .B2(n_689), .Y(n_675) );
INVx1_ASAP7_75t_L g860 ( .A(n_666), .Y(n_860) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
O2A1O1Ixp5_ASAP7_75t_SL g846 ( .A1(n_668), .A2(n_847), .B(n_849), .C(n_853), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g702 ( .A(n_672), .B(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_672), .Y(n_737) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g780 ( .A(n_674), .B(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g746 ( .A(n_678), .Y(n_746) );
AND2x2_ASAP7_75t_L g818 ( .A(n_678), .B(n_819), .Y(n_818) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OR2x6_ASAP7_75t_L g695 ( .A(n_680), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g773 ( .A(n_681), .B(n_749), .Y(n_773) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_686), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g689 ( .A(n_684), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g701 ( .A(n_684), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g728 ( .A(n_684), .B(n_729), .Y(n_728) );
BUFx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_686), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g821 ( .A(n_686), .Y(n_821) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
AND2x2_ASAP7_75t_L g690 ( .A(n_687), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g715 ( .A(n_687), .Y(n_715) );
AND2x2_ASAP7_75t_L g726 ( .A(n_691), .B(n_702), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_710), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_698), .B(n_700), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g834 ( .A(n_702), .Y(n_834) );
BUFx2_ASAP7_75t_L g751 ( .A(n_703), .Y(n_751) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_706), .B(n_708), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_706), .A2(n_858), .B1(n_860), .B2(n_861), .Y(n_857) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI221xp5_ASAP7_75t_SL g710 ( .A1(n_711), .A2(n_716), .B1(n_717), .B2(n_722), .C(n_724), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_714), .B(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g788 ( .A(n_715), .B(n_760), .Y(n_788) );
INVx1_ASAP7_75t_L g873 ( .A(n_715), .Y(n_873) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI22xp33_ASAP7_75t_SL g866 ( .A1(n_718), .A2(n_848), .B1(n_867), .B2(n_868), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
AND2x2_ASAP7_75t_L g748 ( .A(n_719), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g755 ( .A(n_719), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g879 ( .A(n_719), .Y(n_879) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI21xp5_ASAP7_75t_SL g724 ( .A1(n_725), .A2(n_727), .B(n_730), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g785 ( .A(n_726), .Y(n_785) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g844 ( .A(n_729), .B(n_813), .Y(n_844) );
INVx1_ASAP7_75t_L g852 ( .A(n_729), .Y(n_852) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx4_ASAP7_75t_L g756 ( .A(n_732), .Y(n_756) );
NAND2x1_ASAP7_75t_L g796 ( .A(n_732), .B(n_797), .Y(n_796) );
OAI211xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_740), .B(n_742), .C(n_754), .Y(n_733) );
O2A1O1Ixp33_ASAP7_75t_L g799 ( .A1(n_734), .A2(n_800), .B(n_804), .C(n_806), .Y(n_799) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g794 ( .A(n_739), .Y(n_794) );
AOI21xp33_ASAP7_75t_L g853 ( .A1(n_740), .A2(n_823), .B(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_747), .Y(n_743) );
INVx1_ASAP7_75t_L g778 ( .A(n_746), .Y(n_778) );
AND2x2_ASAP7_75t_L g789 ( .A(n_746), .B(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_L g868 ( .A(n_748), .Y(n_868) );
AND2x2_ASAP7_75t_L g841 ( .A(n_749), .B(n_842), .Y(n_841) );
AND2x4_ASAP7_75t_L g750 ( .A(n_751), .B(n_752), .Y(n_750) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OR2x2_ASAP7_75t_L g823 ( .A(n_753), .B(n_767), .Y(n_823) );
INVx1_ASAP7_75t_L g829 ( .A(n_753), .Y(n_829) );
OAI21xp33_ASAP7_75t_SL g754 ( .A1(n_755), .A2(n_757), .B(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g779 ( .A(n_756), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_756), .B(n_797), .Y(n_824) );
OR2x2_ASAP7_75t_L g878 ( .A(n_756), .B(n_879), .Y(n_878) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NOR2x1_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
OR2x2_ASAP7_75t_L g848 ( .A(n_760), .B(n_802), .Y(n_848) );
NOR2x1_ASAP7_75t_L g851 ( .A(n_760), .B(n_852), .Y(n_851) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_845), .Y(n_762) );
NAND4xp25_ASAP7_75t_L g763 ( .A(n_764), .B(n_786), .C(n_809), .D(n_825), .Y(n_763) );
O2A1O1Ixp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_770), .B(n_773), .C(n_774), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OR2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_769), .Y(n_766) );
OR2x2_ASAP7_75t_L g833 ( .A(n_767), .B(n_834), .Y(n_833) );
AND2x4_ASAP7_75t_L g881 ( .A(n_767), .B(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OR2x2_ASAP7_75t_L g802 ( .A(n_768), .B(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g805 ( .A(n_769), .Y(n_805) );
INVx1_ASAP7_75t_L g882 ( .A(n_769), .Y(n_882) );
INVxp67_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
OAI322xp33_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_777), .A3(n_779), .B1(n_780), .B2(n_782), .C1(n_783), .C2(n_785), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g870 ( .A(n_779), .B(n_784), .Y(n_870) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_789), .B1(n_792), .B2(n_795), .C(n_799), .Y(n_786) );
INVxp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g822 ( .A(n_789), .Y(n_822) );
AND2x2_ASAP7_75t_L g816 ( .A(n_791), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g808 ( .A(n_797), .Y(n_808) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OR2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_815), .B(n_820), .Y(n_809) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_L g815 ( .A(n_816), .B(n_818), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_816), .B(n_818), .Y(n_827) );
AND2x4_ASAP7_75t_L g840 ( .A(n_816), .B(n_841), .Y(n_840) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_817), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B1(n_823), .B2(n_824), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_836), .Y(n_825) );
OAI22xp33_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_828), .B1(n_833), .B2(n_835), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
AOI21xp33_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_839), .B(n_843), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NAND3xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_856), .C(n_869), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND2xp67_ASAP7_75t_SL g876 ( .A(n_855), .B(n_877), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g856 ( .A1(n_857), .A2(n_863), .B(n_866), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_871), .B(n_874), .Y(n_869) );
INVxp67_ASAP7_75t_SL g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
BUFx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AOI21xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_890), .B(n_905), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_889), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_896), .Y(n_891) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_892), .Y(n_904) );
INVx6_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
INVx5_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
BUFx6f_ASAP7_75t_L g903 ( .A(n_898), .Y(n_903) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
INVx4_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
INVx3_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx4_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
BUFx6f_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
BUFx12f_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
endmodule