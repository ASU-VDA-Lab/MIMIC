module fake_jpeg_21802_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_31),
.Y(n_48)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_31),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_51),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_20),
.B(n_1),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_28),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_66),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_28),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_65),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_46),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_35),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_20),
.B1(n_30),
.B2(n_43),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_78),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_44),
.B1(n_43),
.B2(n_30),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_44),
.B1(n_43),
.B2(n_58),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_76),
.Y(n_116)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_77),
.A2(n_83),
.B1(n_101),
.B2(n_102),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_44),
.B1(n_30),
.B2(n_20),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_22),
.B1(n_34),
.B2(n_29),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_85),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_44),
.B1(n_22),
.B2(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_82),
.A2(n_87),
.B1(n_96),
.B2(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_40),
.B1(n_38),
.B2(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_84),
.Y(n_115)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_50),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_86),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_22),
.B1(n_29),
.B2(n_23),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_88),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_66),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_90),
.Y(n_140)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_18),
.B1(n_16),
.B2(n_35),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_56),
.A2(n_47),
.B1(n_27),
.B2(n_26),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_40),
.B1(n_38),
.B2(n_47),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_16),
.B1(n_27),
.B2(n_26),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_18),
.Y(n_104)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_64),
.A2(n_46),
.B1(n_38),
.B2(n_21),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_64),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_50),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g108 ( 
.A(n_61),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_46),
.B1(n_19),
.B2(n_42),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_61),
.A2(n_42),
.B1(n_46),
.B2(n_45),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_65),
.A2(n_42),
.A3(n_45),
.B1(n_39),
.B2(n_36),
.Y(n_111)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_129),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_117),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_65),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_72),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_65),
.B(n_67),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_93),
.B(n_49),
.Y(n_162)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_135),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_95),
.Y(n_145)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_73),
.C(n_95),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_150),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_160),
.B(n_166),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_74),
.B1(n_75),
.B2(n_69),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_152),
.B1(n_155),
.B2(n_158),
.Y(n_175)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_123),
.B(n_119),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_69),
.C(n_79),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_143),
.A2(n_74),
.B1(n_79),
.B2(n_70),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_120),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_159),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_154),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_70),
.B1(n_100),
.B2(n_111),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_49),
.C(n_107),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_142),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_70),
.B1(n_100),
.B2(n_103),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_89),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_113),
.B(n_86),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_76),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_145),
.B(n_153),
.Y(n_184)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_163),
.B(n_121),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_110),
.Y(n_164)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_108),
.B1(n_85),
.B2(n_55),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_131),
.B1(n_119),
.B2(n_127),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_0),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_126),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_172),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_0),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_131),
.Y(n_178)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_39),
.Y(n_173)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_184),
.B(n_206),
.Y(n_208)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_181),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_45),
.Y(n_223)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_187),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g188 ( 
.A(n_149),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_190),
.Y(n_220)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_191),
.B(n_194),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_193),
.A2(n_195),
.B1(n_197),
.B2(n_141),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_135),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_127),
.B1(n_123),
.B2(n_140),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_152),
.B1(n_146),
.B2(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_201),
.Y(n_215)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_161),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_202),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_150),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_160),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_126),
.Y(n_204)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_144),
.A2(n_115),
.B(n_137),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_209),
.B(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_162),
.C(n_159),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_214),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_177),
.B(n_147),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_236),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_163),
.C(n_118),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_223),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_146),
.B1(n_171),
.B2(n_166),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_221),
.B1(n_226),
.B2(n_235),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_183),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_219),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_189),
.A2(n_171),
.B1(n_166),
.B2(n_157),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_45),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_225),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_112),
.C(n_138),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_176),
.A2(n_115),
.B(n_84),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_233),
.B(n_174),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_182),
.B(n_36),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_236),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_0),
.B(n_1),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_197),
.A2(n_98),
.B1(n_91),
.B2(n_81),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_36),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_240),
.B(n_241),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_187),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_234),
.B(n_179),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_195),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_250),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_199),
.B1(n_175),
.B2(n_200),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_256),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_191),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_207),
.B(n_201),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_259),
.B1(n_212),
.B2(n_233),
.Y(n_273)
);

A2O1A1O1Ixp25_ASAP7_75t_L g255 ( 
.A1(n_208),
.A2(n_214),
.B(n_213),
.C(n_206),
.D(n_229),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_255),
.B(n_208),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_211),
.A2(n_175),
.B1(n_178),
.B2(n_196),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_215),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_260),
.B1(n_32),
.B2(n_17),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_258),
.A2(n_248),
.B1(n_246),
.B2(n_257),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_178),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_237),
.A2(n_220),
.B1(n_235),
.B2(n_218),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_261),
.A2(n_278),
.B1(n_277),
.B2(n_268),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_262),
.B(n_9),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_243),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_230),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_224),
.C(n_223),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_274),
.C(n_275),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_242),
.A2(n_251),
.B1(n_256),
.B2(n_241),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_221),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_88),
.C(n_36),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_39),
.C(n_60),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_39),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_279),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_117),
.B1(n_32),
.B2(n_17),
.Y(n_278)
);

XOR2x2_ASAP7_75t_SL g279 ( 
.A(n_240),
.B(n_245),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_60),
.C(n_25),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_1),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_285),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_239),
.Y(n_285)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_266),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_32),
.B1(n_17),
.B2(n_25),
.Y(n_289)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_293),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_32),
.B1(n_9),
.B2(n_10),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_291),
.B(n_296),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_297),
.C(n_13),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_8),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_8),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_5),
.B(n_12),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_279),
.A2(n_6),
.B1(n_13),
.B2(n_4),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_11),
.Y(n_297)
);

O2A1O1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_263),
.B1(n_271),
.B2(n_269),
.Y(n_300)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_281),
.B(n_276),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_306),
.C(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_295),
.B(n_299),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g307 ( 
.A1(n_294),
.A2(n_12),
.B(n_13),
.C(n_15),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_307),
.B(n_15),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_12),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_311),
.B(n_292),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_301),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_314),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_282),
.C(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_322),
.C(n_317),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_319),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_282),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_317),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_313),
.A3(n_307),
.B1(n_308),
.B2(n_312),
.C1(n_3),
.C2(n_2),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_284),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_323),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_284),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_303),
.B1(n_323),
.B2(n_310),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_328),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_326),
.B(n_329),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_308),
.C(n_2),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_328),
.Y(n_335)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_2),
.B(n_3),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_333),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_SL g334 ( 
.A1(n_330),
.A2(n_331),
.B(n_324),
.C(n_325),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_334),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_332),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_335),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_336),
.B(n_337),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_327),
.Y(n_342)
);


endmodule