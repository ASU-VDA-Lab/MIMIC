module fake_jpeg_19072_n_121 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx4f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_58),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_0),
.Y(n_61)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_69),
.B(n_71),
.C(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_41),
.B1(n_36),
.B2(n_37),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_38),
.B1(n_46),
.B2(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_82),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_75),
.B(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_43),
.B(n_51),
.C(n_52),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_81),
.B1(n_84),
.B2(n_74),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_3),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_98),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_94),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_53),
.B1(n_47),
.B2(n_42),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_35),
.B1(n_9),
.B2(n_11),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_2),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_34),
.C(n_49),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_95),
.B(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_3),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_96),
.B1(n_88),
.B2(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_104),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_106),
.Y(n_110)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_5),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.C(n_108),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_102),
.C(n_100),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_103),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_101),
.B(n_99),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_101),
.Y(n_121)
);


endmodule