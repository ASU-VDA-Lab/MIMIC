module fake_jpeg_800_n_156 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_156);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_0),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_0),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_46),
.B1(n_52),
.B2(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_59),
.A2(n_53),
.B1(n_54),
.B2(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_50),
.B1(n_49),
.B2(n_47),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_68),
.Y(n_78)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_46),
.B1(n_40),
.B2(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_52),
.C(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_70),
.B(n_51),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_49),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_71),
.C(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_82),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_86),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_38),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_65),
.B1(n_64),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_96),
.B1(n_100),
.B2(n_11),
.Y(n_120)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_66),
.B(n_50),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_95),
.B(n_9),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_48),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_93),
.B1(n_103),
.B2(n_85),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_48),
.B1(n_16),
.B2(n_18),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_1),
.B(n_2),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_102),
.A2(n_85),
.B1(n_73),
.B2(n_10),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_8),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_112),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_25),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_118),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_92),
.B1(n_103),
.B2(n_97),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_28),
.B1(n_34),
.B2(n_20),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_11),
.B(n_12),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_9),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_101),
.B(n_10),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_119),
.B(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_132),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_12),
.B(n_13),
.C(n_21),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_134),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_13),
.B1(n_24),
.B2(n_27),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_141),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_125),
.A2(n_108),
.B(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_137),
.B1(n_112),
.B2(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_147),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_124),
.C(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_143),
.A2(n_138),
.B1(n_139),
.B2(n_127),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_147),
.C(n_126),
.Y(n_150)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_144),
.B(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_148),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_128),
.Y(n_154)
);

AO21x1_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_145),
.B(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_105),
.Y(n_156)
);


endmodule