module fake_jpeg_822_n_450 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_450);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_450;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVxp33_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_55),
.B(n_61),
.Y(n_116)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_56),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_57),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_27),
.A2(n_7),
.B1(n_16),
.B2(n_14),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_59),
.A2(n_39),
.B1(n_34),
.B2(n_54),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_7),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_62),
.Y(n_152)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_64),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_18),
.B(n_6),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_66),
.B(n_67),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_11),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_68),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g167 ( 
.A(n_69),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_70),
.B(n_73),
.Y(n_129)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_42),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_5),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_82),
.Y(n_131)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_12),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_81),
.B(n_89),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_23),
.B(n_12),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_83),
.Y(n_169)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_85),
.B(n_29),
.Y(n_189)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_86),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_12),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_92),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_24),
.B(n_17),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_90),
.Y(n_183)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_91),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_45),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_95),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_47),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_99),
.B(n_104),
.Y(n_181)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_101),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_37),
.B(n_14),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_106),
.Y(n_146)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_51),
.Y(n_124)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_108),
.Y(n_148)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_111),
.Y(n_151)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_29),
.B1(n_50),
.B2(n_51),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_113),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_50),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_43),
.B1(n_54),
.B2(n_22),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_118),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_69),
.A2(n_51),
.B1(n_50),
.B2(n_22),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_124),
.B(n_134),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_57),
.A2(n_43),
.B1(n_39),
.B2(n_44),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_38),
.B1(n_53),
.B2(n_36),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_126),
.A2(n_137),
.B1(n_143),
.B2(n_145),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_67),
.B(n_44),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_41),
.B(n_40),
.C(n_53),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_136),
.B(n_181),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_84),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_140),
.A2(n_157),
.B1(n_162),
.B2(n_177),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_142),
.B(n_159),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_58),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_60),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_1),
.B1(n_4),
.B2(n_62),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_150),
.A2(n_182),
.B1(n_140),
.B2(n_170),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_75),
.A2(n_1),
.B1(n_80),
.B2(n_79),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_64),
.B(n_1),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_78),
.A2(n_102),
.B1(n_88),
.B2(n_65),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_63),
.B(n_113),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_142),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_93),
.A2(n_56),
.B1(n_71),
.B2(n_104),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_166),
.A2(n_128),
.B(n_141),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_74),
.B(n_100),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_168),
.B(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_86),
.B(n_106),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_109),
.B(n_72),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_174),
.B(n_175),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_91),
.B(n_96),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_98),
.B(n_101),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_176),
.B(n_178),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_110),
.A2(n_71),
.B1(n_83),
.B2(n_97),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_66),
.B(n_81),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_66),
.B(n_81),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_186),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_99),
.A2(n_29),
.B1(n_28),
.B2(n_37),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_66),
.B(n_81),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_66),
.B(n_81),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_127),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx4_ASAP7_75t_SL g284 ( 
.A(n_191),
.Y(n_284)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_192),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_193),
.B(n_227),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_124),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_194),
.B(n_199),
.Y(n_254)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_134),
.B(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_201),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_203),
.B(n_212),
.Y(n_272)
);

BUFx12_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx13_ASAP7_75t_L g296 ( 
.A(n_204),
.Y(n_296)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_206),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_130),
.B(n_165),
.C(n_146),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_207),
.B(n_220),
.C(n_237),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_SL g299 ( 
.A1(n_208),
.A2(n_225),
.B(n_234),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_121),
.A2(n_188),
.B1(n_131),
.B2(n_116),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_210),
.A2(n_173),
.B1(n_199),
.B2(n_217),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_245),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_139),
.B(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_215),
.B(n_218),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_130),
.B(n_136),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_181),
.B(n_183),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_223),
.B(n_228),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_123),
.A2(n_120),
.B1(n_167),
.B2(n_185),
.Y(n_225)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_158),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_151),
.B(n_153),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_153),
.B(n_154),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_229),
.B(n_230),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_135),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_231),
.Y(n_265)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_152),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_235),
.Y(n_259)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_233),
.B(n_251),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_177),
.A2(n_157),
.B1(n_120),
.B2(n_164),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_152),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_236),
.B(n_238),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_155),
.B(n_166),
.C(n_164),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_155),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_119),
.B(n_160),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_241),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_141),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_252),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_119),
.B(n_160),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_132),
.B(n_185),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_244),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_147),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_243),
.B(n_250),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_132),
.B(n_138),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_133),
.A2(n_135),
.B1(n_167),
.B2(n_138),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_163),
.B(n_147),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_194),
.Y(n_286)
);

AO21x2_ASAP7_75t_L g282 ( 
.A1(n_248),
.A2(n_249),
.B(n_247),
.Y(n_282)
);

BUFx12_ASAP7_75t_L g249 ( 
.A(n_128),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_163),
.B(n_133),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_167),
.A2(n_173),
.B1(n_169),
.B2(n_190),
.Y(n_251)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_173),
.A2(n_99),
.B1(n_29),
.B2(n_140),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_253),
.A2(n_211),
.B1(n_249),
.B2(n_224),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_255),
.B(n_260),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_196),
.A2(n_193),
.B1(n_226),
.B2(n_220),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_260),
.A2(n_295),
.B1(n_293),
.B2(n_274),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_209),
.A2(n_248),
.B(n_222),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_267),
.A2(n_293),
.B(n_255),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_294),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_282),
.A2(n_297),
.B(n_270),
.C(n_298),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_216),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_213),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_289),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g288 ( 
.A1(n_226),
.A2(n_211),
.B1(n_202),
.B2(n_251),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_299),
.B1(n_257),
.B2(n_267),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_213),
.B(n_200),
.Y(n_289)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_207),
.B(n_221),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_291),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_191),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_205),
.B(n_233),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_292),
.B(n_284),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_237),
.A2(n_227),
.B1(n_239),
.B2(n_244),
.Y(n_293)
);

AND2x2_ASAP7_75t_SL g294 ( 
.A(n_241),
.B(n_242),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_197),
.A2(n_206),
.B1(n_231),
.B2(n_198),
.Y(n_295)
);

O2A1O1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_245),
.A2(n_204),
.B(n_235),
.C(n_238),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_271),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_300),
.B(n_304),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_238),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_301),
.B(n_328),
.C(n_319),
.Y(n_361)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_303),
.B(n_312),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_307),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_262),
.B(n_252),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_308),
.B(n_315),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_270),
.A2(n_204),
.B(n_235),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_254),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_321),
.B1(n_326),
.B2(n_301),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_254),
.B(n_283),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_314),
.B(n_320),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_268),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_316),
.Y(n_343)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_256),
.Y(n_317)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_317),
.Y(n_358)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_261),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_324),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_333),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_283),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_288),
.A2(n_282),
.B1(n_257),
.B2(n_275),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_322),
.A2(n_282),
.B1(n_280),
.B2(n_298),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_256),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_323),
.B(n_325),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_285),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_268),
.B(n_278),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_272),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_329),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_294),
.C(n_277),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_330),
.B(n_331),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_258),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_285),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_332),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_279),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_334),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_336),
.A2(n_342),
.B1(n_346),
.B2(n_351),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_330),
.A2(n_298),
.B1(n_297),
.B2(n_259),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_337),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_333),
.A2(n_273),
.B(n_265),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_339),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_306),
.A2(n_284),
.B1(n_269),
.B2(n_273),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_313),
.A2(n_295),
.B1(n_261),
.B2(n_266),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_322),
.A2(n_266),
.B1(n_276),
.B2(n_258),
.Y(n_346)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_316),
.A2(n_296),
.B(n_263),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_359),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_326),
.A2(n_263),
.B1(n_269),
.B2(n_296),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_361),
.B(n_310),
.C(n_321),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_345),
.B(n_325),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_368),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_361),
.B(n_328),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_350),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_367),
.C(n_371),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_312),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_315),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_357),
.B(n_331),
.Y(n_369)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_341),
.Y(n_370)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_323),
.C(n_314),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_320),
.Y(n_372)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_372),
.Y(n_391)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_373),
.Y(n_400)
);

XOR2x1_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_306),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_379),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_306),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_356),
.C(n_303),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_305),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_378),
.Y(n_393)
);

XNOR2x2_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_311),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_340),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_380),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_355),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_382),
.Y(n_395)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_327),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_360),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_367),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_348),
.C(n_358),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_389),
.C(n_379),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_343),
.B(n_338),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_392),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_356),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_375),
.B(n_354),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_336),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_376),
.A2(n_354),
.B1(n_343),
.B2(n_353),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_399),
.A2(n_364),
.B1(n_370),
.B2(n_373),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_401),
.A2(n_391),
.B1(n_397),
.B2(n_392),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_405),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_386),
.B(n_377),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_412),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_396),
.A2(n_376),
.B1(n_359),
.B2(n_374),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_409),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_395),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_408),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_395),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_366),
.C(n_371),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_410),
.B(n_413),
.C(n_384),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_388),
.A2(n_374),
.B1(n_372),
.B2(n_353),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_411),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_400),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_414),
.A2(n_390),
.B1(n_355),
.B2(n_344),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_417),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_402),
.C(n_389),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_401),
.A2(n_391),
.B1(n_365),
.B2(n_364),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_385),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_407),
.A2(n_365),
.B(n_399),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_422),
.A2(n_347),
.B(n_335),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_424),
.A2(n_393),
.B(n_407),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_431),
.B(n_423),
.Y(n_434)
);

AO22x2_ASAP7_75t_SL g426 ( 
.A1(n_420),
.A2(n_417),
.B1(n_422),
.B2(n_413),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_426),
.B(n_419),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_412),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_427),
.B(n_429),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_421),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_L g431 ( 
.A1(n_421),
.A2(n_387),
.B(n_405),
.C(n_410),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_432),
.B(n_423),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_434),
.A2(n_435),
.B(n_308),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_436),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_437),
.B(n_433),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_428),
.A2(n_415),
.B(n_347),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_438),
.A2(n_429),
.B(n_436),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_439),
.B(n_441),
.Y(n_445)
);

NAND4xp25_ASAP7_75t_L g443 ( 
.A(n_440),
.B(n_426),
.C(n_414),
.D(n_418),
.Y(n_443)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_443),
.Y(n_446)
);

AOI322xp5_ASAP7_75t_L g444 ( 
.A1(n_442),
.A2(n_358),
.A3(n_348),
.B1(n_344),
.B2(n_346),
.C1(n_347),
.C2(n_418),
.Y(n_444)
);

INVxp33_ASAP7_75t_L g447 ( 
.A(n_444),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_446),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_448),
.B(n_447),
.C(n_445),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_398),
.Y(n_450)
);


endmodule