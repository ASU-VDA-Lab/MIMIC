module fake_jpeg_10619_n_142 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_21),
.B1(n_15),
.B2(n_26),
.Y(n_49)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx5_ASAP7_75t_SL g41 ( 
.A(n_34),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_16),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_14),
.Y(n_42)
);

OA21x2_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_46),
.B(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_15),
.B1(n_21),
.B2(n_26),
.Y(n_60)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_56),
.B1(n_57),
.B2(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_41),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_10),
.C(n_11),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_9),
.Y(n_85)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_36),
.B1(n_37),
.B2(n_30),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_64),
.B1(n_70),
.B2(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_63),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_66),
.B1(n_31),
.B2(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_17),
.Y(n_87)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_36),
.B1(n_37),
.B2(n_24),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_20),
.B(n_43),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_31),
.B1(n_34),
.B2(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_19),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_31),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_46),
.Y(n_79)
);

NAND2x1_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_65),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_87),
.B1(n_56),
.B2(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_86),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_11),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_1),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_79),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_87),
.B1(n_83),
.B2(n_77),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_100),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_38),
.B(n_32),
.C(n_53),
.D(n_61),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_61),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_82),
.C(n_80),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_77),
.C(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_106),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_93),
.B(n_92),
.C(n_99),
.D(n_89),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_111),
.C(n_93),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_78),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_112),
.C(n_98),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_88),
.B(n_98),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_118),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_116),
.C(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_88),
.C(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_96),
.B1(n_105),
.B2(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_103),
.C(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_125),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_107),
.C(n_95),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_95),
.C(n_76),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_85),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_129),
.B(n_130),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_122),
.B(n_67),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_85),
.B(n_4),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_131),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_54),
.B1(n_17),
.B2(n_23),
.Y(n_135)
);

AOI322xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_17),
.A3(n_22),
.B1(n_23),
.B2(n_6),
.C1(n_2),
.C2(n_32),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_137),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_22),
.B(n_23),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_138),
.A2(n_136),
.B(n_23),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_22),
.B1(n_38),
.B2(n_139),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_22),
.Y(n_142)
);


endmodule