module fake_jpeg_14333_n_40 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_40);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_15),
.A2(n_12),
.B1(n_11),
.B2(n_8),
.Y(n_21)
);

OAI32xp33_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_13),
.A3(n_14),
.B1(n_3),
.B2(n_4),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_0),
.Y(n_26)
);

XOR2x2_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_26),
.Y(n_30)
);

AND2x6_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_31),
.B1(n_22),
.B2(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_25),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_5),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_35),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_22),
.B1(n_14),
.B2(n_5),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_34),
.B(n_32),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_2),
.B(n_3),
.Y(n_39)
);


endmodule