module real_jpeg_17142_n_22 (n_17, n_8, n_0, n_21, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_16, n_15, n_13, n_22);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;

output n_22;

wire n_43;
wire n_57;
wire n_37;
wire n_54;
wire n_65;
wire n_33;
wire n_38;
wire n_50;
wire n_35;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_31;
wire n_58;
wire n_52;
wire n_67;
wire n_63;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_28;
wire n_60;
wire n_44;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_71;
wire n_47;
wire n_45;
wire n_25;
wire n_61;
wire n_51;
wire n_42;
wire n_53;
wire n_39;
wire n_40;
wire n_36;
wire n_70;
wire n_41;
wire n_27;
wire n_26;
wire n_32;
wire n_48;
wire n_30;
wire n_56;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_1),
.A2(n_15),
.B1(n_39),
.B2(n_43),
.Y(n_42)
);

OAI211xp5_ASAP7_75t_L g63 ( 
.A1(n_1),
.A2(n_16),
.B(n_64),
.C(n_66),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

OAI222xp33_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_5),
.B1(n_8),
.B2(n_27),
.C1(n_28),
.C2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

AOI221xp5_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.C(n_50),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_8),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_8),
.A2(n_10),
.B(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

OAI31xp33_ASAP7_75t_L g29 ( 
.A1(n_10),
.A2(n_19),
.A3(n_30),
.B(n_31),
.Y(n_29)
);

AOI222xp33_ASAP7_75t_L g37 ( 
.A1(n_11),
.A2(n_13),
.B1(n_15),
.B2(n_38),
.C1(n_39),
.C2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_11),
.B(n_14),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_13),
.B(n_46),
.Y(n_49)
);

AOI221xp5_ASAP7_75t_SL g67 ( 
.A1(n_13),
.A2(n_64),
.B1(n_68),
.B2(n_69),
.C(n_71),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_14),
.B(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_15),
.Y(n_65)
);

OAI221xp5_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.C(n_37),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

AOI31xp33_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_26),
.A3(n_32),
.B(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_17),
.A2(n_26),
.B(n_32),
.Y(n_35)
);

AOI31xp33_ASAP7_75t_L g56 ( 
.A1(n_17),
.A2(n_20),
.A3(n_57),
.B(n_61),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_17),
.A2(n_57),
.B(n_61),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_24),
.A3(n_41),
.B1(n_44),
.B2(n_55),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_18),
.A2(n_37),
.B(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

OAI321xp33_ASAP7_75t_SL g57 ( 
.A1(n_27),
.A2(n_28),
.A3(n_31),
.B1(n_33),
.B2(n_58),
.C(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_28),
.B(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_39),
.B1(n_43),
.B2(n_65),
.Y(n_68)
);

AOI222xp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.C1(n_48),
.C2(n_65),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_48),
.B(n_70),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND4xp25_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.C(n_53),
.D(n_54),
.Y(n_50)
);

NOR4xp25_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.C(n_53),
.D(n_54),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.A3(n_63),
.B1(n_67),
.B2(n_72),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);


endmodule