module fake_jpeg_228_n_61 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_31;
wire n_25;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx5_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_20),
.A2(n_29),
.B1(n_32),
.B2(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_15),
.B(n_1),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_31),
.C(n_23),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_28),
.B1(n_18),
.B2(n_9),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_11),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_8),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_13),
.A2(n_9),
.B1(n_19),
.B2(n_18),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_13),
.B1(n_19),
.B2(n_16),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);

OAI221xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_22),
.C(n_36),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_33),
.C(n_39),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_34),
.B(n_41),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_44),
.C(n_33),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.C(n_22),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_44),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_37),
.B(n_29),
.Y(n_57)
);

AOI31xp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_57),
.A3(n_38),
.B(n_40),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_53),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_59),
.C(n_40),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_42),
.B(n_21),
.Y(n_61)
);


endmodule