module real_jpeg_4340_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_493;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_0),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_0),
.B(n_180),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_0),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_0),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_0),
.B(n_282),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_0),
.B(n_324),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_0),
.B(n_303),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_0),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_1),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_1),
.B(n_93),
.Y(n_160)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_1),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_1),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_1),
.B(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_1),
.B(n_341),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_1),
.B(n_405),
.Y(n_404)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_2),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_2),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_2),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_3),
.Y(n_528)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_4),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g231 ( 
.A(n_4),
.Y(n_231)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_4),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_5),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_5),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_5),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_5),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_5),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_5),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_5),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_6),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_6),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_6),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_6),
.B(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_6),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_6),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_6),
.B(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_7),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_7),
.Y(n_226)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_8),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_9),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_9),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_9),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_9),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_9),
.B(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_10),
.Y(n_202)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_10),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_10),
.Y(n_309)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_12),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_12),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_12),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_13),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_13),
.B(n_42),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_13),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_13),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_13),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_13),
.B(n_279),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_13),
.B(n_375),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_13),
.B(n_98),
.Y(n_401)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_15),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_48),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_15),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_15),
.B(n_32),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_15),
.B(n_216),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_15),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_15),
.B(n_324),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_15),
.B(n_171),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_16),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_16),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_16),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_16),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_16),
.B(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_16),
.B(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_16),
.B(n_174),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_17),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_17),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_17),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_17),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_17),
.B(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_17),
.B(n_382),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_17),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_18),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_18),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_18),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_18),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_18),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_18),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_18),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_18),
.B(n_254),
.Y(n_253)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_523),
.B(n_525),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_38),
.B(n_76),
.C(n_522),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_24),
.B(n_43),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.C(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_26),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_26),
.A2(n_29),
.B1(n_37),
.B2(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_27),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_47),
.B1(n_53),
.B2(n_54),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_47),
.C(n_55),
.Y(n_73)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_33),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_34),
.B(n_75),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_72),
.C(n_74),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_44),
.B(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_59),
.C(n_62),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_45),
.B(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_55),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_47),
.A2(n_54),
.B1(n_68),
.B2(n_111),
.Y(n_115)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_49),
.B(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_51),
.Y(n_145)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_52),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_52),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_63),
.C(n_68),
.Y(n_62)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_59),
.B(n_62),
.Y(n_118)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_63),
.A2(n_64),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_68),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_68),
.A2(n_106),
.B1(n_107),
.B2(n_111),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_70),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_70),
.Y(n_214)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_70),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_70),
.Y(n_405)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_71),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_71),
.Y(n_347)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_71),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_74),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_122),
.B(n_521),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_119),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_78),
.B(n_119),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_116),
.C(n_117),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_79),
.A2(n_80),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_104),
.C(n_112),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_81),
.A2(n_82),
.B1(n_497),
.B2(n_499),
.Y(n_496)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_91),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_87),
.C(n_91),
.Y(n_116)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_86),
.Y(n_263)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_86),
.Y(n_395)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.C(n_99),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_92),
.B(n_487),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_487)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_104),
.A2(n_112),
.B1(n_113),
.B2(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_104),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.C(n_111),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_105),
.B(n_493),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_106),
.A2(n_107),
.B1(n_188),
.B2(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_107),
.B(n_185),
.C(n_188),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_116),
.B(n_117),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_515),
.B(n_520),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_480),
.B(n_512),
.Y(n_123)
);

OAI21x1_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_291),
.B(n_479),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_239),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_126),
.B(n_239),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_182),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_127),
.B(n_183),
.C(n_217),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_158),
.C(n_165),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_128),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.C(n_146),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_129),
.B(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_133),
.C(n_134),
.Y(n_164)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_136),
.A2(n_137),
.B1(n_146),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_144),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_138),
.B(n_144),
.Y(n_454)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_141),
.B(n_454),
.Y(n_453)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_146),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_147),
.B(n_149),
.C(n_154),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_149),
.Y(n_157)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_153),
.B(n_188),
.C(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_153),
.A2(n_154),
.B1(n_188),
.B2(n_192),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_156),
.Y(n_254)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_156),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_158),
.B(n_165),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_161),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_162),
.C(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_161),
.A2(n_163),
.B1(n_228),
.B2(n_232),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_163),
.B(n_222),
.C(n_232),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_164),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_176),
.C(n_179),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_166),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.C(n_173),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_167),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_170),
.B(n_173),
.Y(n_251)
);

BUFx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_172),
.Y(n_266)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_176),
.B(n_179),
.Y(n_271)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_181),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_217),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_193),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_184),
.B(n_194),
.C(n_206),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_206),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.C(n_203),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_203),
.Y(n_238)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_198),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_198),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_202),
.Y(n_279)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_215),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_208),
.B(n_211),
.C(n_215),
.Y(n_495)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_233),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_219),
.B(n_221),
.C(n_233),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.C(n_237),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_237),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.C(n_246),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_241),
.B(n_244),
.Y(n_474)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_246),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_269),
.C(n_272),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_248),
.B(n_467),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.C(n_259),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_249),
.A2(n_250),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_252),
.A2(n_253),
.B(n_255),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_252),
.B(n_259),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.C(n_267),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_422)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_267),
.B(n_422),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_268),
.B(n_363),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_272),
.Y(n_468)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_284),
.C(n_288),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_274),
.B(n_456),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_275),
.B(n_434),
.Y(n_433)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_278),
.A2(n_280),
.B1(n_281),
.B2(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_278),
.Y(n_435)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_284),
.B(n_288),
.Y(n_456)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g403 ( 
.A(n_286),
.Y(n_403)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_289),
.Y(n_393)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_472),
.B(n_478),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_459),
.B(n_471),
.Y(n_292)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_441),
.B(n_458),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_415),
.B(n_440),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_386),
.B(n_414),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_355),
.B(n_385),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_336),
.B(n_354),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_316),
.B(n_335),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_310),
.B(n_315),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_308),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_308),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_306),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_306),
.Y(n_317)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_305),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

INVx4_ASAP7_75t_SL g363 ( 
.A(n_309),
.Y(n_363)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_318),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_325),
.B2(n_326),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_328),
.C(n_331),
.Y(n_353)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_323),
.Y(n_343)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_331),
.B2(n_332),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_353),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_353),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_344),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_343),
.C(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_342),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_344),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_348),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_371),
.C(n_372),
.Y(n_370)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_352),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_358),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_369),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_359),
.B(n_370),
.C(n_373),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_362),
.C(n_364),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_365),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_368),
.Y(n_396)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_373),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_378),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_381),
.C(n_383),
.Y(n_412)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_379),
.A2(n_381),
.B1(n_383),
.B2(n_384),
.Y(n_378)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_379),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_381),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_413),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_387),
.B(n_413),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_398),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_397),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_389),
.B(n_397),
.C(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_396),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_394),
.Y(n_390)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_391),
.Y(n_429)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_394),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_429),
.C(n_430),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_406),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_408),
.C(n_411),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_404),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

MAJx2_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_402),
.C(n_404),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_408),
.B1(n_411),
.B2(n_412),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_409),
.B(n_410),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_438),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_438),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_427),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_419),
.C(n_427),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_423),
.B2(n_424),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_450),
.C(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_425),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_431),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_432),
.C(n_437),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_436),
.B2(n_437),
.Y(n_431)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_432),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_433),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_457),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_457),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_448),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_447),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_447),
.C(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_445),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_449),
.B(n_453),
.C(n_455),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_469),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_460),
.B(n_469),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_461),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_463),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_476),
.C(n_477),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_475),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_473),
.B(n_475),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_508),
.Y(n_480)
);

OAI21xp33_ASAP7_75t_L g512 ( 
.A1(n_481),
.A2(n_513),
.B(n_514),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_501),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_482),
.B(n_501),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_484),
.B1(n_490),
.B2(n_500),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_483),
.B(n_491),
.C(n_496),
.Y(n_519)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.C(n_488),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_503),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_486),
.A2(n_488),
.B1(n_489),
.B2(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_486),
.Y(n_504)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_490),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_496),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_494),
.C(n_495),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_506),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_495),
.Y(n_506)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_497),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_505),
.C(n_507),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_505),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_507),
.B(n_510),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_509),
.B(n_511),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_509),
.B(n_511),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_519),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_519),
.Y(n_520)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_517),
.Y(n_518)
);

INVx8_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_524),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_528),
.Y(n_525)
);

BUFx12f_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);


endmodule