module fake_aes_7014_n_27 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_1), .Y(n_11) );
NOR2x1p5_ASAP7_75t_L g12 ( .A(n_3), .B(n_9), .Y(n_12) );
BUFx3_ASAP7_75t_L g13 ( .A(n_0), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_11), .B(n_10), .Y(n_15) );
OAI22xp5_ASAP7_75t_L g16 ( .A1(n_14), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_14), .B(n_3), .Y(n_17) );
OAI22xp5_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_16), .B(n_13), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_19), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_21), .B1(n_20), .B2(n_18), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
BUFx2_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
OAI22x1_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_12), .B1(n_6), .B2(n_8), .Y(n_26) );
AOI22xp5_ASAP7_75t_SL g27 ( .A1(n_26), .A2(n_13), .B1(n_5), .B2(n_8), .Y(n_27) );
endmodule