module real_jpeg_17178_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_258;
wire n_205;
wire n_61;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_216;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

AND2x4_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_58),
.Y(n_57)
);

AND2x4_ASAP7_75t_SL g69 ( 
.A(n_0),
.B(n_70),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_0),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_0),
.B(n_52),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_0),
.Y(n_136)
);

NAND2x1p5_ASAP7_75t_L g177 ( 
.A(n_0),
.B(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_2),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_3),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_3),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_3),
.B(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_4),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_5),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_5),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_5),
.B(n_36),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_5),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_5),
.B(n_178),
.Y(n_241)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_7),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_7),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_7),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_7),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_7),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_7),
.B(n_216),
.Y(n_215)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_8),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_8),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_9),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g222 ( 
.A(n_10),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_11),
.Y(n_178)
);

BUFx8_ASAP7_75t_L g216 ( 
.A(n_11),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_230),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_228),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_193),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_155),
.B(n_192),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_122),
.B(n_154),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_92),
.B(n_121),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_21),
.B(n_74),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_23),
.B(n_39),
.C(n_53),
.Y(n_123)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_25),
.B(n_31),
.C(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_31),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_31),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_34),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_34),
.A2(n_151),
.B1(n_165),
.B2(n_171),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_37),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.C(n_49),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_40),
.A2(n_41),
.B1(n_49),
.B2(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_40),
.A2(n_41),
.B1(n_166),
.B2(n_170),
.Y(n_248)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_41),
.B(n_205),
.Y(n_204)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_41),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_45),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_44),
.A2(n_45),
.B1(n_144),
.B2(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_45),
.A2(n_104),
.B(n_113),
.C(n_145),
.Y(n_161)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_49),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_49),
.A2(n_77),
.B1(n_128),
.B2(n_140),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_86),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_50),
.B(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_65),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_55),
.A2(n_110),
.B(n_114),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_55),
.A2(n_66),
.B(n_73),
.Y(n_141)
);

NOR2x1_ASAP7_75t_R g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_56),
.A2(n_57),
.B1(n_84),
.B2(n_85),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_69),
.B(n_71),
.Y(n_68)
);

NAND2x1p5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_69),
.Y(n_71)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

O2A1O1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_95),
.B(n_98),
.C(n_104),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_95),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_66),
.A2(n_72),
.B1(n_95),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_80),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_69),
.B(n_99),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_69),
.A2(n_90),
.B1(n_99),
.B2(n_102),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_71),
.B(n_128),
.C(n_135),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.C(n_88),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_77),
.B(n_140),
.C(n_200),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_88),
.B1(n_89),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_80),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_84),
.A2(n_85),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_85),
.B(n_215),
.C(n_219),
.Y(n_260)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_108),
.B(n_120),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.Y(n_93)
);

NOR2xp67_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_105),
.Y(n_120)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_95),
.B(n_112),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_95),
.B(n_113),
.C(n_177),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_95),
.A2(n_118),
.B1(n_204),
.B2(n_208),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_95),
.B(n_206),
.Y(n_246)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_99),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_99),
.A2(n_102),
.B1(n_166),
.B2(n_170),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_99),
.B(n_151),
.C(n_166),
.Y(n_225)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_116),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_115),
.B(n_119),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_112),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_113),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_118),
.B(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_124),
.Y(n_154)
);

XOR2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_142),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_141),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_126),
.B(n_141),
.C(n_142),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_134),
.B1(n_135),
.B2(n_140),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_148),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_149),
.C(n_153),
.Y(n_158)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_191),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_191),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_172),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_159),
.C(n_172),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_164),
.C(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_190),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_180),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_180),
.C(n_190),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_187),
.B(n_189),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_187),
.Y(n_189)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_195),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_211),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_196),
.B(n_212),
.C(n_227),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_209),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_202),
.B2(n_203),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_202),
.C(n_209),
.Y(n_234)
);

XNOR2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_227),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_223),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_225),
.C(n_226),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_264),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_263),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_263),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_249),
.B2(n_250),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2x2_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_247),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_261),
.B2(n_262),
.Y(n_252)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_254),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);


endmodule