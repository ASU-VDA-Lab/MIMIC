module real_jpeg_3032_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_1),
.A2(n_26),
.B1(n_38),
.B2(n_41),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_1),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_1),
.A2(n_26),
.B1(n_69),
.B2(n_71),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_37),
.B1(n_58),
.B2(n_59),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_37),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_37),
.B1(n_69),
.B2(n_71),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_2),
.B(n_59),
.C(n_67),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_65),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_2),
.B(n_38),
.C(n_53),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_2),
.B(n_23),
.C(n_45),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_2),
.B(n_51),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_29),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_2),
.B(n_179),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_5),
.A2(n_38),
.B1(n_41),
.B2(n_70),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_70),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_33),
.B1(n_38),
.B2(n_41),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_9),
.A2(n_33),
.B1(n_69),
.B2(n_71),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_9),
.A2(n_33),
.B1(n_58),
.B2(n_59),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_308),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_270),
.B(n_305),
.Y(n_14)
);

A2O1A1O1Ixp25_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_131),
.B(n_250),
.C(n_251),
.D(n_269),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_109),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_17),
.B(n_109),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_76),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_18),
.B(n_77),
.C(n_103),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_50),
.C(n_62),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_19),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_34),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_20),
.B(n_34),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_30),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_21),
.A2(n_28),
.B(n_84),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_22),
.A2(n_23),
.B1(n_44),
.B2(n_45),
.Y(n_47)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_23),
.B(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_27),
.B(n_32),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_27),
.A2(n_28),
.B(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_27),
.B(n_83),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_27),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_28),
.B(n_208),
.Y(n_222)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_29),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_30),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_31),
.B(n_207),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_48),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_35),
.B(n_193),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_36),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_36),
.B(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_41),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_38),
.B(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_42),
.B(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_42),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_48),
.A2(n_87),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_48),
.B(n_180),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_50),
.A2(n_62),
.B1(n_63),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_50),
.A2(n_113),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B(n_61),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_51),
.B(n_61),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_51),
.B(n_124),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_51),
.A2(n_147),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_53),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_55),
.B(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_56),
.B(n_99),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_56),
.A2(n_284),
.B(n_285),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_59),
.B(n_175),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_72),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_65),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_74)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_72),
.A2(n_262),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_102),
.B2(n_103),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_89),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_79),
.B(n_90),
.C(n_97),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_85),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_81),
.B(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_84),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

AOI21x1_ASAP7_75t_SL g144 ( 
.A1(n_86),
.A2(n_107),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_86),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_88),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_88),
.B(n_178),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_96),
.B2(n_97),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_94),
.B(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_94),
.A2(n_142),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_98),
.B(n_122),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_98),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_101),
.B(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_104),
.A2(n_105),
.B1(n_173),
.B2(n_174),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_104),
.A2(n_105),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_105),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_105),
.B(n_106),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_105),
.A2(n_258),
.B(n_260),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_106),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_130),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_110),
.A2(n_111),
.B1(n_130),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_114),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_125),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_117),
.B(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_117),
.A2(n_142),
.B(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_120),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_130),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_241),
.B(n_247),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_165),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_151),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_134),
.B(n_151),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_135),
.B(n_138),
.C(n_150),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_150),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_146),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_141),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_143),
.A2(n_144),
.B1(n_283),
.B2(n_286),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_143),
.A2(n_144),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_144),
.B(n_278),
.C(n_283),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_144),
.B(n_302),
.C(n_304),
.Y(n_314)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_147),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.C(n_158),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_152),
.A2(n_153),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_158),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.C(n_161),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_164),
.B(n_222),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_185),
.B(n_240),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_182),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_167),
.B(n_182),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.C(n_176),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_169),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_176),
.B1(n_177),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI21x1_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_196),
.B(n_239),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_191),
.Y(n_239)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_188),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.C(n_195),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_194),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_234),
.B(n_238),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_216),
.B(n_233),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_204),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_209),
.B1(n_210),
.B2(n_215),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_213),
.C(n_215),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_223),
.B(n_232),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_220),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_228),
.B(n_231),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_230),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_236),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_246),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_253),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_256),
.C(n_264),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_263),
.B2(n_264),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B(n_268),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_266),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_268),
.A2(n_276),
.B1(n_277),
.B2(n_287),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_268),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_274),
.C(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_288),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_273),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_279),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_291),
.C(n_295),
.Y(n_315)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_283),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_290),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_299),
.B1(n_300),
.B2(n_304),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_297),
.Y(n_304)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_315),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_310),
.B(n_315),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_312),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);


endmodule