module real_aes_8100_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_252;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g537 ( .A1(n_0), .A2(n_184), .B(n_538), .C(n_541), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_1), .B(n_526), .Y(n_542) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_91), .C(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g429 ( .A(n_2), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_3), .A2(n_748), .B1(n_751), .B2(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_3), .Y(n_752) );
INVx1_ASAP7_75t_L g202 ( .A(n_4), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_5), .B(n_173), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_6), .A2(n_441), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_7), .A2(n_149), .B(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_8), .A2(n_36), .B1(n_129), .B2(n_138), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_9), .B(n_149), .Y(n_213) );
AND2x6_ASAP7_75t_L g147 ( .A(n_10), .B(n_148), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_11), .A2(n_147), .B(n_444), .C(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_12), .B(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_12), .B(n_37), .Y(n_430) );
INVx1_ASAP7_75t_L g145 ( .A(n_13), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_14), .B(n_136), .Y(n_156) );
INVx1_ASAP7_75t_L g194 ( .A(n_15), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_16), .B(n_173), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_17), .B(n_150), .Y(n_218) );
AO32x2_ASAP7_75t_L g181 ( .A1(n_18), .A2(n_146), .A3(n_149), .B1(n_182), .B2(n_186), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_19), .B(n_138), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_20), .B(n_150), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_21), .A2(n_52), .B1(n_129), .B2(n_138), .Y(n_185) );
AOI22xp33_ASAP7_75t_SL g135 ( .A1(n_22), .A2(n_82), .B1(n_136), .B2(n_138), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_23), .B(n_138), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g443 ( .A1(n_24), .A2(n_146), .B(n_444), .C(n_446), .Y(n_443) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_25), .A2(n_146), .B(n_444), .C(n_491), .Y(n_490) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_26), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_27), .B(n_141), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_28), .A2(n_441), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_29), .B(n_141), .Y(n_179) );
INVx2_ASAP7_75t_L g131 ( .A(n_30), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_31), .A2(n_465), .B(n_474), .C(n_476), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_32), .B(n_138), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_33), .B(n_141), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g113 ( .A1(n_34), .A2(n_73), .B1(n_114), .B2(n_115), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_34), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_35), .B(n_158), .Y(n_492) );
INVx1_ASAP7_75t_L g106 ( .A(n_37), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_38), .B(n_440), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_39), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_40), .B(n_173), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_41), .B(n_441), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_42), .A2(n_465), .B(n_474), .C(n_511), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_43), .A2(n_119), .B1(n_423), .B2(n_424), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g423 ( .A(n_43), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_43), .A2(n_79), .B1(n_423), .B2(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_44), .B(n_138), .Y(n_208) );
INVx1_ASAP7_75t_L g539 ( .A(n_45), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_46), .A2(n_90), .B1(n_129), .B2(n_132), .Y(n_128) );
INVx1_ASAP7_75t_L g512 ( .A(n_47), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_48), .B(n_138), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_49), .B(n_138), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_50), .B(n_441), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_51), .B(n_200), .Y(n_212) );
AOI22xp33_ASAP7_75t_SL g222 ( .A1(n_53), .A2(n_58), .B1(n_136), .B2(n_138), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_54), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_55), .B(n_138), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_56), .B(n_138), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_57), .Y(n_756) );
INVx1_ASAP7_75t_L g148 ( .A(n_59), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_60), .B(n_441), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_61), .B(n_526), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_62), .A2(n_197), .B(n_200), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_63), .B(n_138), .Y(n_203) );
INVx1_ASAP7_75t_L g144 ( .A(n_64), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_65), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_66), .B(n_173), .Y(n_478) );
AO32x2_ASAP7_75t_L g126 ( .A1(n_67), .A2(n_127), .A3(n_140), .B1(n_146), .B2(n_149), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_68), .B(n_139), .Y(n_502) );
INVx1_ASAP7_75t_L g236 ( .A(n_69), .Y(n_236) );
INVx1_ASAP7_75t_L g171 ( .A(n_70), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_71), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_72), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g460 ( .A1(n_74), .A2(n_444), .B(n_461), .C(n_465), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_75), .B(n_136), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_76), .Y(n_521) );
INVx1_ASAP7_75t_L g110 ( .A(n_77), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_78), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_79), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_80), .A2(n_103), .B1(n_111), .B2(n_759), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_81), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_83), .B(n_129), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_84), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_85), .B(n_136), .Y(n_176) );
INVx2_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_87), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_88), .B(n_133), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_89), .B(n_136), .Y(n_209) );
OR2x2_ASAP7_75t_L g427 ( .A(n_91), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g727 ( .A(n_91), .Y(n_727) );
OR2x2_ASAP7_75t_L g746 ( .A(n_91), .B(n_740), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_92), .A2(n_101), .B1(n_136), .B2(n_137), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_93), .B(n_441), .Y(n_472) );
INVx1_ASAP7_75t_L g477 ( .A(n_94), .Y(n_477) );
INVxp67_ASAP7_75t_L g524 ( .A(n_95), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_96), .B(n_136), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_97), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g462 ( .A(n_98), .Y(n_462) );
INVx1_ASAP7_75t_L g498 ( .A(n_99), .Y(n_498) );
AND2x2_ASAP7_75t_L g514 ( .A(n_100), .B(n_141), .Y(n_514) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx6p67_ASAP7_75t_R g760 ( .A(n_104), .Y(n_760) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO221x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_741), .B1(n_744), .B2(n_753), .C(n_755), .Y(n_111) );
OAI222xp33_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_116), .B1(n_728), .B2(n_729), .C1(n_735), .C2(n_736), .Y(n_112) );
INVx1_ASAP7_75t_L g728 ( .A(n_113), .Y(n_728) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_425), .B1(n_431), .B2(n_724), .Y(n_117) );
INVx1_ASAP7_75t_L g731 ( .A(n_118), .Y(n_731) );
INVx2_ASAP7_75t_L g424 ( .A(n_119), .Y(n_424) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
XOR2x2_ASAP7_75t_L g748 ( .A(n_120), .B(n_749), .Y(n_748) );
AND3x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_343), .C(n_391), .Y(n_120) );
NOR4xp25_ASAP7_75t_L g121 ( .A(n_122), .B(n_271), .C(n_316), .D(n_330), .Y(n_121) );
OAI311xp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_187), .A3(n_214), .B1(n_224), .C1(n_239), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_151), .Y(n_123) );
OAI21xp33_ASAP7_75t_L g224 ( .A1(n_124), .A2(n_225), .B(n_227), .Y(n_224) );
AND2x2_ASAP7_75t_L g332 ( .A(n_124), .B(n_259), .Y(n_332) );
AND2x2_ASAP7_75t_L g389 ( .A(n_124), .B(n_275), .Y(n_389) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g282 ( .A(n_125), .B(n_180), .Y(n_282) );
AND2x2_ASAP7_75t_L g339 ( .A(n_125), .B(n_287), .Y(n_339) );
INVx1_ASAP7_75t_L g380 ( .A(n_125), .Y(n_380) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_126), .Y(n_248) );
AND2x2_ASAP7_75t_L g289 ( .A(n_126), .B(n_180), .Y(n_289) );
AND2x2_ASAP7_75t_L g293 ( .A(n_126), .B(n_181), .Y(n_293) );
INVx1_ASAP7_75t_L g305 ( .A(n_126), .Y(n_305) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_133), .B1(n_135), .B2(n_139), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx3_ASAP7_75t_L g132 ( .A(n_130), .Y(n_132) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
AND2x6_ASAP7_75t_L g444 ( .A(n_130), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g137 ( .A(n_131), .Y(n_137) );
INVx1_ASAP7_75t_L g201 ( .A(n_131), .Y(n_201) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_132), .Y(n_479) );
INVx2_ASAP7_75t_L g541 ( .A(n_132), .Y(n_541) );
INVx2_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_133), .A2(n_183), .B1(n_184), .B2(n_185), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_133), .A2(n_184), .B1(n_221), .B2(n_222), .Y(n_220) );
INVx4_ASAP7_75t_L g540 ( .A(n_133), .Y(n_540) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx3_ASAP7_75t_L g139 ( .A(n_134), .Y(n_139) );
INVx1_ASAP7_75t_L g158 ( .A(n_134), .Y(n_158) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
AND2x2_ASAP7_75t_L g442 ( .A(n_134), .B(n_201), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_134), .Y(n_445) );
INVx2_ASAP7_75t_L g195 ( .A(n_136), .Y(n_195) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_138), .Y(n_464) );
INVx5_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
INVx1_ASAP7_75t_L g451 ( .A(n_140), .Y(n_451) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OA21x2_ASAP7_75t_L g152 ( .A1(n_141), .A2(n_153), .B(n_163), .Y(n_152) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_141), .A2(n_168), .B(n_179), .Y(n_167) );
INVx1_ASAP7_75t_L g454 ( .A(n_141), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_141), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_141), .A2(n_509), .B(n_510), .Y(n_508) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_L g150 ( .A(n_142), .B(n_143), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
NAND3xp33_ASAP7_75t_L g219 ( .A(n_146), .B(n_220), .C(n_223), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_146), .A2(n_232), .B(n_235), .Y(n_231) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_147), .A2(n_154), .B(n_159), .Y(n_153) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_147), .A2(n_169), .B(n_174), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_147), .A2(n_193), .B(n_198), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_147), .A2(n_207), .B(n_210), .Y(n_206) );
AND2x4_ASAP7_75t_L g441 ( .A(n_147), .B(n_442), .Y(n_441) );
INVx4_ASAP7_75t_SL g466 ( .A(n_147), .Y(n_466) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_147), .B(n_442), .Y(n_499) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_149), .A2(n_206), .B(n_213), .Y(n_205) );
INVx4_ASAP7_75t_L g223 ( .A(n_149), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_149), .A2(n_489), .B(n_490), .Y(n_488) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_149), .Y(n_518) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_164), .Y(n_151) );
AND2x2_ASAP7_75t_L g226 ( .A(n_152), .B(n_180), .Y(n_226) );
INVx2_ASAP7_75t_L g260 ( .A(n_152), .Y(n_260) );
AND2x2_ASAP7_75t_L g275 ( .A(n_152), .B(n_181), .Y(n_275) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_152), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_152), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g295 ( .A(n_152), .B(n_258), .Y(n_295) );
INVx1_ASAP7_75t_L g307 ( .A(n_152), .Y(n_307) );
INVx1_ASAP7_75t_L g348 ( .A(n_152), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_152), .B(n_248), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_157), .Y(n_154) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_162), .Y(n_159) );
O2A1O1Ixp5_ASAP7_75t_L g235 ( .A1(n_162), .A2(n_199), .B(n_236), .C(n_237), .Y(n_235) );
NOR2xp67_ASAP7_75t_L g164 ( .A(n_165), .B(n_180), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g225 ( .A(n_166), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_166), .Y(n_253) );
AND2x2_ASAP7_75t_SL g306 ( .A(n_166), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g310 ( .A(n_166), .B(n_180), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_166), .B(n_305), .Y(n_368) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g258 ( .A(n_167), .Y(n_258) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_167), .Y(n_274) );
OR2x2_ASAP7_75t_L g347 ( .A(n_167), .B(n_348), .Y(n_347) );
O2A1O1Ixp5_ASAP7_75t_SL g169 ( .A1(n_170), .A2(n_171), .B(n_172), .C(n_173), .Y(n_169) );
INVx2_ASAP7_75t_L g184 ( .A(n_173), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_173), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_173), .A2(n_233), .B(n_234), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_173), .B(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .Y(n_174) );
INVx1_ASAP7_75t_L g197 ( .A(n_177), .Y(n_197) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g448 ( .A(n_178), .Y(n_448) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx2_ASAP7_75t_L g254 ( .A(n_181), .Y(n_254) );
AND2x2_ASAP7_75t_L g259 ( .A(n_181), .B(n_260), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_184), .A2(n_199), .B(n_202), .C(n_203), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_184), .A2(n_211), .B(n_212), .Y(n_210) );
INVx2_ASAP7_75t_L g191 ( .A(n_186), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_186), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_187), .B(n_242), .Y(n_405) );
INVx1_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g375 ( .A(n_188), .B(n_216), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_205), .Y(n_188) );
AND2x2_ASAP7_75t_L g251 ( .A(n_189), .B(n_242), .Y(n_251) );
INVx2_ASAP7_75t_L g263 ( .A(n_189), .Y(n_263) );
AND2x2_ASAP7_75t_L g297 ( .A(n_189), .B(n_245), .Y(n_297) );
AND2x2_ASAP7_75t_L g364 ( .A(n_189), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_190), .B(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g244 ( .A(n_190), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g284 ( .A(n_190), .B(n_205), .Y(n_284) );
AND2x2_ASAP7_75t_L g301 ( .A(n_190), .B(n_302), .Y(n_301) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_204), .Y(n_190) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_191), .A2(n_231), .B(n_238), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .C(n_197), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_195), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_195), .A2(n_502), .B(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_197), .A2(n_462), .B(n_463), .C(n_464), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_199), .A2(n_447), .B(n_449), .Y(n_446) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g227 ( .A(n_205), .B(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g245 ( .A(n_205), .Y(n_245) );
AND2x2_ASAP7_75t_L g250 ( .A(n_205), .B(n_230), .Y(n_250) );
AND2x2_ASAP7_75t_L g323 ( .A(n_205), .B(n_302), .Y(n_323) );
AND2x2_ASAP7_75t_L g388 ( .A(n_205), .B(n_378), .Y(n_388) );
OAI311xp33_ASAP7_75t_L g271 ( .A1(n_214), .A2(n_272), .A3(n_276), .B1(n_278), .C1(n_298), .Y(n_271) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g283 ( .A(n_215), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g342 ( .A(n_215), .B(n_250), .Y(n_342) );
AND2x2_ASAP7_75t_L g416 ( .A(n_215), .B(n_297), .Y(n_416) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_216), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g351 ( .A(n_216), .Y(n_351) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g242 ( .A(n_217), .Y(n_242) );
NOR2x1_ASAP7_75t_L g314 ( .A(n_217), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g371 ( .A(n_217), .B(n_245), .Y(n_371) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
INVx1_ASAP7_75t_L g268 ( .A(n_218), .Y(n_268) );
AO21x1_ASAP7_75t_L g267 ( .A1(n_220), .A2(n_223), .B(n_268), .Y(n_267) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_223), .A2(n_459), .B(n_468), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_223), .B(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_223), .B(n_481), .Y(n_480) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_223), .A2(n_497), .B(n_504), .Y(n_496) );
INVx3_ASAP7_75t_L g526 ( .A(n_223), .Y(n_526) );
AND2x2_ASAP7_75t_L g246 ( .A(n_226), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g299 ( .A(n_226), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g379 ( .A(n_226), .B(n_380), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_227), .A2(n_259), .B1(n_279), .B2(n_283), .C(n_285), .Y(n_278) );
INVx1_ASAP7_75t_L g403 ( .A(n_228), .Y(n_403) );
OR2x2_ASAP7_75t_L g369 ( .A(n_229), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g264 ( .A(n_230), .B(n_245), .Y(n_264) );
OR2x2_ASAP7_75t_L g266 ( .A(n_230), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g291 ( .A(n_230), .Y(n_291) );
INVx2_ASAP7_75t_L g302 ( .A(n_230), .Y(n_302) );
AND2x2_ASAP7_75t_L g329 ( .A(n_230), .B(n_267), .Y(n_329) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_230), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_246), .B1(n_249), .B2(n_252), .C(n_255), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
AND2x2_ASAP7_75t_L g340 ( .A(n_242), .B(n_250), .Y(n_340) );
AND2x2_ASAP7_75t_L g390 ( .A(n_242), .B(n_244), .Y(n_390) );
INVx2_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g277 ( .A(n_244), .B(n_248), .Y(n_277) );
AND2x2_ASAP7_75t_L g356 ( .A(n_244), .B(n_329), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_245), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g315 ( .A(n_245), .Y(n_315) );
OAI21xp33_ASAP7_75t_L g325 ( .A1(n_246), .A2(n_326), .B(n_328), .Y(n_325) );
OR2x2_ASAP7_75t_L g269 ( .A(n_247), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g335 ( .A(n_247), .B(n_295), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_247), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g312 ( .A(n_248), .B(n_281), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_248), .B(n_395), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_249), .B(n_275), .Y(n_385) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g308 ( .A(n_250), .B(n_263), .Y(n_308) );
INVx1_ASAP7_75t_L g324 ( .A(n_251), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_261), .B1(n_265), .B2(n_269), .Y(n_255) );
INVx2_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g287 ( .A(n_258), .Y(n_287) );
INVx1_ASAP7_75t_L g300 ( .A(n_258), .Y(n_300) );
INVx1_ASAP7_75t_L g270 ( .A(n_259), .Y(n_270) );
AND2x2_ASAP7_75t_L g341 ( .A(n_259), .B(n_287), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_259), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
OR2x2_ASAP7_75t_L g265 ( .A(n_262), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_262), .B(n_378), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_262), .B(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g412 ( .A(n_264), .B(n_364), .Y(n_412) );
INVx1_ASAP7_75t_SL g378 ( .A(n_266), .Y(n_378) );
AND2x2_ASAP7_75t_L g318 ( .A(n_267), .B(n_302), .Y(n_318) );
INVx1_ASAP7_75t_L g365 ( .A(n_267), .Y(n_365) );
OAI222xp33_ASAP7_75t_L g406 ( .A1(n_272), .A2(n_362), .B1(n_407), .B2(n_408), .C1(n_411), .C2(n_413), .Y(n_406) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g327 ( .A(n_274), .Y(n_327) );
AND2x2_ASAP7_75t_L g338 ( .A(n_275), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_275), .B(n_380), .Y(n_407) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_277), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g382 ( .A(n_279), .Y(n_382) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_SL g320 ( .A(n_282), .Y(n_320) );
AND2x2_ASAP7_75t_L g399 ( .A(n_282), .B(n_360), .Y(n_399) );
AND2x2_ASAP7_75t_L g422 ( .A(n_282), .B(n_306), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_284), .B(n_318), .Y(n_317) );
OAI32xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .A3(n_290), .B1(n_292), .B2(n_296), .Y(n_285) );
BUFx2_ASAP7_75t_L g360 ( .A(n_287), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_288), .B(n_306), .Y(n_387) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g326 ( .A(n_289), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g394 ( .A(n_289), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g383 ( .A(n_290), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AND2x2_ASAP7_75t_L g354 ( .A(n_293), .B(n_327), .Y(n_354) );
INVx2_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OAI221xp5_ASAP7_75t_SL g316 ( .A1(n_295), .A2(n_317), .B1(n_319), .B2(n_321), .C(n_325), .Y(n_316) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g328 ( .A(n_297), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g334 ( .A(n_297), .B(n_318), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B1(n_303), .B2(n_308), .C(n_309), .Y(n_298) );
INVx1_ASAP7_75t_L g417 ( .A(n_299), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_300), .B(n_394), .Y(n_393) );
NAND2x1p5_ASAP7_75t_L g313 ( .A(n_301), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_306), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g372 ( .A(n_306), .Y(n_372) );
BUFx3_ASAP7_75t_L g395 ( .A(n_307), .Y(n_395) );
INVx1_ASAP7_75t_SL g336 ( .A(n_308), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_308), .B(n_350), .Y(n_349) );
AOI21xp33_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_311), .B(n_313), .Y(n_309) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_310), .A2(n_411), .B1(n_415), .B2(n_417), .C(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g357 ( .A(n_315), .B(n_318), .Y(n_357) );
INVx1_ASAP7_75t_L g421 ( .A(n_315), .Y(n_421) );
INVx2_ASAP7_75t_L g410 ( .A(n_318), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_318), .B(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g363 ( .A(n_323), .B(n_364), .Y(n_363) );
OAI221xp5_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_333), .B1(n_335), .B2(n_336), .C(n_337), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_340), .B1(n_341), .B2(n_342), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_339), .A2(n_401), .B1(n_402), .B2(n_404), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_342), .A2(n_419), .B(n_422), .Y(n_418) );
NOR4xp25_ASAP7_75t_SL g343 ( .A(n_344), .B(n_352), .C(n_361), .D(n_381), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B1(n_358), .B2(n_359), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_366), .B1(n_369), .B2(n_372), .C(n_373), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g384 ( .A(n_364), .Y(n_384) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI21xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_376), .B(n_379), .Y(n_373) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI211xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_385), .C(n_386), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_389), .B2(n_390), .Y(n_386) );
CKINVDCx14_ASAP7_75t_R g396 ( .A(n_390), .Y(n_396) );
NOR3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_406), .C(n_414), .Y(n_391) );
OAI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B1(n_397), .B2(n_398), .C(n_400), .Y(n_392) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
CKINVDCx16_ASAP7_75t_R g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g732 ( .A(n_426), .Y(n_732) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g726 ( .A(n_428), .B(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g740 ( .A(n_428), .Y(n_740) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g733 ( .A(n_432), .Y(n_733) );
AND3x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_628), .C(n_685), .Y(n_432) );
NOR3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_573), .C(n_609), .Y(n_433) );
OAI211xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_482), .B(n_528), .C(n_560), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_455), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g531 ( .A(n_437), .B(n_532), .Y(n_531) );
INVx5_ASAP7_75t_L g559 ( .A(n_437), .Y(n_559) );
AND2x2_ASAP7_75t_L g632 ( .A(n_437), .B(n_548), .Y(n_632) );
AND2x2_ASAP7_75t_L g670 ( .A(n_437), .B(n_576), .Y(n_670) );
AND2x2_ASAP7_75t_L g690 ( .A(n_437), .B(n_533), .Y(n_690) );
OR2x6_ASAP7_75t_L g437 ( .A(n_438), .B(n_452), .Y(n_437) );
AOI21xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_443), .B(n_451), .Y(n_438) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx5_ASAP7_75t_L g475 ( .A(n_444), .Y(n_475) );
INVx2_ASAP7_75t_L g450 ( .A(n_448), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_450), .A2(n_477), .B(n_478), .C(n_479), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_450), .A2(n_479), .B(n_512), .C(n_513), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_455), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_470), .Y(n_455) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_456), .Y(n_571) );
AND2x2_ASAP7_75t_L g585 ( .A(n_456), .B(n_532), .Y(n_585) );
INVx1_ASAP7_75t_L g608 ( .A(n_456), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_456), .B(n_559), .Y(n_647) );
OR2x2_ASAP7_75t_L g684 ( .A(n_456), .B(n_530), .Y(n_684) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_457), .Y(n_620) );
AND2x2_ASAP7_75t_L g627 ( .A(n_457), .B(n_533), .Y(n_627) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g548 ( .A(n_458), .B(n_533), .Y(n_548) );
BUFx2_ASAP7_75t_L g576 ( .A(n_458), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_466), .A2(n_475), .B(n_521), .C(n_522), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_466), .A2(n_475), .B(n_536), .C(n_537), .Y(n_535) );
INVx5_ASAP7_75t_L g530 ( .A(n_470), .Y(n_530) );
BUFx2_ASAP7_75t_L g552 ( .A(n_470), .Y(n_552) );
AND2x2_ASAP7_75t_L g709 ( .A(n_470), .B(n_563), .Y(n_709) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_515), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g609 ( .A1(n_484), .A2(n_610), .B1(n_617), .B2(n_618), .C(n_621), .Y(n_609) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
AND2x2_ASAP7_75t_L g516 ( .A(n_485), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_485), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g544 ( .A(n_486), .B(n_495), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_486), .B(n_496), .Y(n_554) );
OR2x2_ASAP7_75t_L g565 ( .A(n_486), .B(n_517), .Y(n_565) );
AND2x2_ASAP7_75t_L g568 ( .A(n_486), .B(n_556), .Y(n_568) );
AND2x2_ASAP7_75t_L g584 ( .A(n_486), .B(n_506), .Y(n_584) );
OR2x2_ASAP7_75t_L g600 ( .A(n_486), .B(n_496), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_486), .B(n_517), .Y(n_662) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_487), .B(n_506), .Y(n_654) );
AND2x2_ASAP7_75t_L g657 ( .A(n_487), .B(n_496), .Y(n_657) );
OR2x2_ASAP7_75t_L g578 ( .A(n_494), .B(n_565), .Y(n_578) );
INVx2_ASAP7_75t_L g604 ( .A(n_494), .Y(n_604) );
OR2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_506), .Y(n_494) );
AND2x2_ASAP7_75t_L g527 ( .A(n_495), .B(n_507), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_495), .B(n_517), .Y(n_583) );
OR2x2_ASAP7_75t_L g594 ( .A(n_495), .B(n_507), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_495), .B(n_556), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g686 ( .A1(n_495), .A2(n_687), .B1(n_689), .B2(n_691), .C(n_694), .Y(n_686) );
INVx5_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_496), .B(n_517), .Y(n_625) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_500), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_506), .B(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_506), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g572 ( .A(n_506), .B(n_544), .Y(n_572) );
OR2x2_ASAP7_75t_L g616 ( .A(n_506), .B(n_517), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_506), .B(n_568), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_506), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g681 ( .A(n_506), .B(n_682), .Y(n_681) );
INVx5_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_SL g545 ( .A(n_507), .B(n_516), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_507), .A2(n_550), .B(n_553), .C(n_557), .Y(n_549) );
OR2x2_ASAP7_75t_L g587 ( .A(n_507), .B(n_583), .Y(n_587) );
OR2x2_ASAP7_75t_L g623 ( .A(n_507), .B(n_565), .Y(n_623) );
OAI311xp33_ASAP7_75t_L g629 ( .A1(n_507), .A2(n_568), .A3(n_630), .B1(n_633), .C1(n_640), .Y(n_629) );
AND2x2_ASAP7_75t_L g680 ( .A(n_507), .B(n_517), .Y(n_680) );
AND2x2_ASAP7_75t_L g688 ( .A(n_507), .B(n_543), .Y(n_688) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_507), .Y(n_706) );
AND2x2_ASAP7_75t_L g723 ( .A(n_507), .B(n_544), .Y(n_723) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_527), .Y(n_515) );
AND2x2_ASAP7_75t_L g551 ( .A(n_516), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g707 ( .A(n_516), .Y(n_707) );
AND2x2_ASAP7_75t_L g543 ( .A(n_517), .B(n_544), .Y(n_543) );
INVx3_ASAP7_75t_L g556 ( .A(n_517), .Y(n_556) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_517), .Y(n_599) );
INVxp67_ASAP7_75t_L g638 ( .A(n_517), .Y(n_638) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_525), .Y(n_517) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_526), .A2(n_534), .B(n_542), .Y(n_533) );
AND2x2_ASAP7_75t_L g716 ( .A(n_527), .B(n_564), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_543), .B1(n_545), .B2(n_546), .C(n_549), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_530), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g569 ( .A(n_530), .B(n_559), .Y(n_569) );
AND2x2_ASAP7_75t_L g577 ( .A(n_530), .B(n_532), .Y(n_577) );
OR2x2_ASAP7_75t_L g589 ( .A(n_530), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g607 ( .A(n_530), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g631 ( .A(n_530), .B(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_530), .Y(n_651) );
AND2x2_ASAP7_75t_L g703 ( .A(n_530), .B(n_627), .Y(n_703) );
OAI31xp33_ASAP7_75t_L g711 ( .A1(n_530), .A2(n_580), .A3(n_679), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_531), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g675 ( .A(n_531), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_531), .B(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g563 ( .A(n_532), .B(n_559), .Y(n_563) );
INVx1_ASAP7_75t_L g650 ( .A(n_532), .Y(n_650) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g700 ( .A(n_533), .B(n_559), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_SL g710 ( .A(n_543), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_544), .B(n_615), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_545), .A2(n_657), .B1(n_695), .B2(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g558 ( .A(n_548), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g617 ( .A(n_548), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_548), .B(n_569), .Y(n_722) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g692 ( .A(n_551), .B(n_693), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_552), .A2(n_611), .B(n_613), .Y(n_610) );
OR2x2_ASAP7_75t_L g618 ( .A(n_552), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g639 ( .A(n_552), .B(n_627), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_552), .B(n_650), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_552), .B(n_690), .Y(n_689) );
OAI221xp5_ASAP7_75t_SL g666 ( .A1(n_553), .A2(n_667), .B1(n_672), .B2(n_675), .C(n_676), .Y(n_666) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
OR2x2_ASAP7_75t_L g643 ( .A(n_554), .B(n_616), .Y(n_643) );
INVx1_ASAP7_75t_L g682 ( .A(n_554), .Y(n_682) );
INVx2_ASAP7_75t_L g658 ( .A(n_555), .Y(n_658) );
INVx1_ASAP7_75t_L g592 ( .A(n_556), .Y(n_592) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g597 ( .A(n_559), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_559), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g626 ( .A(n_559), .B(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g714 ( .A(n_559), .B(n_684), .Y(n_714) );
AOI222xp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B1(n_566), .B2(n_569), .C1(n_570), .C2(n_572), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g570 ( .A(n_563), .B(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_563), .A2(n_613), .B1(n_641), .B2(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_563), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
OAI21xp33_ASAP7_75t_SL g601 ( .A1(n_572), .A2(n_602), .B(n_605), .Y(n_601) );
OAI211xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_578), .B(n_579), .C(n_601), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_577), .A2(n_580), .B1(n_585), .B2(n_586), .C(n_588), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_577), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g671 ( .A(n_577), .Y(n_671) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
AND2x2_ASAP7_75t_L g673 ( .A(n_582), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g590 ( .A(n_585), .Y(n_590) );
AND2x2_ASAP7_75t_L g596 ( .A(n_585), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B1(n_595), .B2(n_598), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_592), .B(n_604), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_593), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g693 ( .A(n_597), .Y(n_693) );
AND2x2_ASAP7_75t_L g712 ( .A(n_597), .B(n_627), .Y(n_712) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_604), .B(n_661), .Y(n_720) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_607), .B(n_675), .Y(n_718) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g641 ( .A(n_619), .Y(n_641) );
BUFx2_ASAP7_75t_L g665 ( .A(n_620), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g621 ( .A1(n_622), .A2(n_624), .B(n_626), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_644), .C(n_666), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_639), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_648), .B(n_652), .C(n_655), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_645), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NOR2xp67_ASAP7_75t_SL g649 ( .A(n_650), .B(n_651), .Y(n_649) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_SL g674 ( .A(n_654), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_659), .B(n_663), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
AND2x2_ASAP7_75t_L g679 ( .A(n_657), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B1(n_681), .B2(n_683), .Y(n_676) );
INVx2_ASAP7_75t_SL g697 ( .A(n_684), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_701), .C(n_713), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_697), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B1(n_708), .B2(n_710), .C(n_711), .Y(n_701) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_702), .A2(n_714), .B(n_715), .C(n_717), .Y(n_713) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B1(n_721), .B2(n_723), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g734 ( .A(n_725), .Y(n_734) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_727), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_730) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
BUFx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_SL g754 ( .A(n_742), .Y(n_754) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g758 ( .A(n_746), .Y(n_758) );
INVx1_ASAP7_75t_L g751 ( .A(n_748), .Y(n_751) );
BUFx3_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
endmodule