module fake_jpeg_18841_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_16),
.B(n_6),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_14),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_46),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_0),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_49),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_20),
.B1(n_28),
.B2(n_19),
.Y(n_61)
);

CKINVDCx9p33_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_51),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_29),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_60),
.C(n_21),
.Y(n_87)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_67),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_35),
.C(n_23),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_48),
.B1(n_20),
.B2(n_18),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_28),
.B1(n_34),
.B2(n_33),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_26),
.B1(n_25),
.B2(n_24),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_46),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_92),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_72),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_73),
.B(n_84),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_36),
.B1(n_18),
.B2(n_34),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_78),
.B1(n_81),
.B2(n_88),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_75),
.A2(n_105),
.B1(n_104),
.B2(n_106),
.Y(n_117)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_98),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_83),
.B(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_52),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_94),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_33),
.B1(n_25),
.B2(n_26),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_24),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_67),
.C(n_57),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_11),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_41),
.C(n_40),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_97),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_51),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_97),
.B1(n_86),
.B2(n_82),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_44),
.Y(n_97)
);

FAx1_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_44),
.CI(n_32),
.CON(n_98),
.SN(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_50),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_99),
.A2(n_101),
.B1(n_32),
.B2(n_23),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_103),
.Y(n_116)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_10),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_35),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_22),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_58),
.A2(n_23),
.B1(n_22),
.B2(n_35),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_107),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_64),
.B1(n_23),
.B2(n_22),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_117),
.B1(n_133),
.B2(n_81),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_127),
.B1(n_129),
.B2(n_105),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_132),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_0),
.B(n_1),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_73),
.C(n_89),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_22),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_132),
.B(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_137),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_136),
.A2(n_139),
.B1(n_145),
.B2(n_116),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_75),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_78),
.B1(n_69),
.B2(n_97),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_109),
.B(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_143),
.B(n_149),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_124),
.B1(n_108),
.B2(n_107),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_118),
.B1(n_110),
.B2(n_133),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_82),
.B1(n_101),
.B2(n_93),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_107),
.B(n_71),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_99),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_76),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_100),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_154),
.B(n_110),
.Y(n_161)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_134),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_156),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_113),
.B(n_102),
.Y(n_156)
);

OA21x2_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_113),
.B(n_110),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_5),
.B(n_11),
.C(n_130),
.D(n_2),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_156),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_166),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_121),
.B1(n_123),
.B2(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_169),
.B1(n_176),
.B2(n_180),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_144),
.B1(n_141),
.B2(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_123),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_172),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_128),
.B(n_116),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_147),
.B(n_154),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_116),
.B1(n_114),
.B2(n_121),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_157),
.B1(n_151),
.B2(n_135),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_114),
.Y(n_178)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_126),
.B1(n_122),
.B2(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_181),
.Y(n_185)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_191),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_142),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_197),
.C(n_201),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_190),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_174),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_157),
.B1(n_151),
.B2(n_138),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_181),
.B1(n_175),
.B2(n_179),
.Y(n_204)
);

AOI221xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_138),
.B1(n_151),
.B2(n_122),
.C(n_5),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_130),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_199),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_173),
.C(n_164),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_212),
.B1(n_203),
.B2(n_192),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_182),
.A2(n_179),
.B(n_171),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_205),
.A2(n_191),
.B(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_182),
.B1(n_183),
.B2(n_185),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_186),
.C(n_197),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_216),
.C(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_217),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_169),
.B1(n_172),
.B2(n_165),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_165),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_189),
.C(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_208),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_220),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_228),
.B(n_205),
.Y(n_236)
);

NOR3xp33_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_163),
.C(n_193),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_233),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_225),
.B1(n_162),
.B2(n_159),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_163),
.B1(n_167),
.B2(n_170),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_230),
.C(n_231),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_213),
.C(n_216),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_164),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_232),
.Y(n_245)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_235),
.C(n_245),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_207),
.C(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_241),
.Y(n_247)
);

XNOR2x1_ASAP7_75t_SL g238 ( 
.A(n_220),
.B(n_207),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_242),
.B(n_228),
.C(n_226),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_240),
.B(n_165),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

AOI21x1_ASAP7_75t_SL g242 ( 
.A1(n_232),
.A2(n_215),
.B(n_212),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_159),
.B(n_167),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_235),
.C(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_229),
.B1(n_219),
.B2(n_178),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_233),
.C(n_166),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_256),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_238),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_2),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_240),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_244),
.B(n_242),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_255),
.A2(n_249),
.B(n_246),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_262),
.C(n_263),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_258),
.A2(n_165),
.B(n_11),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_254),
.C(n_3),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_267),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_265),
.B(n_3),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_3),
.C(n_4),
.Y(n_271)
);


endmodule