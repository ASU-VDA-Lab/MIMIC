module fake_jpeg_18091_n_260 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_260);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_260;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx6_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_49),
.Y(n_69)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_54),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_56),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_36),
.Y(n_76)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_17),
.B1(n_26),
.B2(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_17),
.B1(n_26),
.B2(n_29),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_17),
.B1(n_29),
.B2(n_31),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_49),
.B1(n_28),
.B2(n_31),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_38),
.B1(n_32),
.B2(n_28),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_18),
.B1(n_32),
.B2(n_25),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_43),
.B1(n_54),
.B2(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_35),
.B(n_37),
.C(n_27),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_19),
.B(n_23),
.C(n_24),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_25),
.B1(n_22),
.B2(n_37),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_30),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_80),
.Y(n_127)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_44),
.C(n_41),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_116),
.B(n_57),
.C(n_44),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_85),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_22),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_88),
.A2(n_100),
.B1(n_108),
.B2(n_112),
.Y(n_140)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_19),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_91),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_23),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_101),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_27),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_65),
.B(n_14),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_104),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_107),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_46),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_111),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_57),
.B(n_34),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_41),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_114),
.B1(n_73),
.B2(n_63),
.Y(n_131)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_115),
.A2(n_76),
.B1(n_73),
.B2(n_78),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_59),
.B(n_44),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_118),
.B1(n_125),
.B2(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_83),
.B1(n_97),
.B2(n_106),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_116),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_73),
.B1(n_78),
.B2(n_61),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_84),
.A2(n_94),
.B1(n_115),
.B2(n_99),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_152),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_146),
.B1(n_131),
.B2(n_117),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_153),
.C(n_154),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_99),
.B1(n_114),
.B2(n_82),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_132),
.B(n_92),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_147),
.B(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_105),
.Y(n_148)
);

NOR2x1_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_80),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_149),
.A2(n_137),
.B(n_138),
.C(n_88),
.Y(n_177)
);

BUFx8_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g165 ( 
.A(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_101),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_89),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_120),
.C(n_124),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_95),
.C(n_93),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_158),
.Y(n_162)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_103),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_119),
.B(n_107),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_108),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_87),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_161),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_176),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_127),
.B1(n_126),
.B2(n_140),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_173),
.B1(n_180),
.B2(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_126),
.B1(n_125),
.B2(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_137),
.C(n_132),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_179),
.C(n_181),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

OAI321xp33_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_143),
.A3(n_135),
.B1(n_136),
.B2(n_51),
.C(n_68),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_137),
.C(n_138),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_145),
.A2(n_110),
.B1(n_81),
.B2(n_104),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_134),
.C(n_123),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_170),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_189),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_186),
.B(n_194),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_136),
.B1(n_156),
.B2(n_149),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_146),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_191),
.C(n_195),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_155),
.C(n_159),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_175),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_196),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_147),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_135),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_134),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_199),
.C(n_168),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_123),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_163),
.B(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_203),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_178),
.A3(n_177),
.B1(n_162),
.B2(n_173),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_207),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_178),
.C(n_180),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_211),
.Y(n_222)
);

OAI322xp33_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_177),
.A3(n_165),
.B1(n_30),
.B2(n_3),
.C1(n_5),
.C2(n_6),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_209),
.B(n_10),
.Y(n_226)
);

OAI321xp33_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_177),
.A3(n_122),
.B1(n_150),
.B2(n_30),
.C(n_86),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_10),
.B1(n_15),
.B2(n_2),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_193),
.C(n_196),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_177),
.A3(n_150),
.B1(n_122),
.B2(n_98),
.C1(n_68),
.C2(n_6),
.Y(n_212)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_212),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_63),
.C(n_150),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_0),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_198),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_217),
.A2(n_16),
.B1(n_5),
.B2(n_10),
.Y(n_237)
);

FAx1_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_197),
.CI(n_190),
.CON(n_218),
.SN(n_218)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_226),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_7),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_220),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_6),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_227),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_225),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_228),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_218),
.A2(n_214),
.B1(n_211),
.B2(n_201),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_11),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_11),
.C(n_3),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_221),
.C(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_218),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_231),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_230),
.B(n_236),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_217),
.B(n_223),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_242),
.B(n_244),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_236),
.B1(n_230),
.B2(n_224),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_238),
.B(n_229),
.C(n_234),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_249),
.B(n_250),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_253),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_242),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_16),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_256),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_258),
.B(n_16),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_255),
.A2(n_252),
.B(n_12),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_1),
.Y(n_260)
);


endmodule