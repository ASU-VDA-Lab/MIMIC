module fake_jpeg_15114_n_18 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_18);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_18;

wire n_13;
wire n_16;
wire n_10;
wire n_9;
wire n_14;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;

INVx6_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

AOI22xp33_ASAP7_75t_L g10 ( 
.A1(n_1),
.A2(n_0),
.B1(n_5),
.B2(n_3),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_1),
.Y(n_14)
);

AOI21x1_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_15),
.B(n_13),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_2),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_10),
.Y(n_17)
);

AOI322xp5_ASAP7_75t_L g18 ( 
.A1(n_17),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_16),
.C2(n_15),
.Y(n_18)
);


endmodule