module fake_jpeg_2356_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_41),
.Y(n_43)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_31),
.B(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_40),
.Y(n_47)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_15),
.B(n_10),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_10),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_9),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_54),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_14),
.B1(n_23),
.B2(n_21),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_50),
.B1(n_21),
.B2(n_35),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_13),
.B1(n_26),
.B2(n_19),
.Y(n_50)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_8),
.Y(n_52)
);

OAI32xp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_17),
.A3(n_41),
.B1(n_25),
.B2(n_9),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_26),
.B1(n_19),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_30),
.A2(n_27),
.B1(n_14),
.B2(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_67),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_68),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_36),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_71),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_41),
.C(n_35),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_33),
.B(n_25),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_50),
.B(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_33),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_55),
.B(n_46),
.C(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_90),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_48),
.B1(n_61),
.B2(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_86),
.B1(n_45),
.B2(n_64),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_73),
.B1(n_65),
.B2(n_71),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_58),
.B(n_59),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_38),
.B1(n_53),
.B2(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_74),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_70),
.C(n_63),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_86),
.B1(n_81),
.B2(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_107),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_100),
.C(n_96),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_84),
.C(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_SL g111 ( 
.A1(n_101),
.A2(n_82),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_1),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_97),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_94),
.C(n_99),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_118),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_100),
.B(n_104),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_113),
.B(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_109),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_82),
.B(n_5),
.C(n_6),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_123),
.C(n_82),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_113),
.B1(n_105),
.B2(n_96),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_117),
.A3(n_119),
.B1(n_112),
.B2(n_109),
.C1(n_114),
.C2(n_89),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_125),
.B(n_126),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_122),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_122),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_129),
.B(n_128),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_4),
.Y(n_131)
);


endmodule