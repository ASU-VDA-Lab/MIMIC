module fake_jpeg_13212_n_295 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_295);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_245;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_51),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_55),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_54),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_0),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_39),
.Y(n_100)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_29),
.B(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_39),
.Y(n_76)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_72),
.B(n_100),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_73),
.A2(n_85),
.B(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_76),
.B(n_83),
.Y(n_143)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_62),
.C(n_58),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_79),
.B(n_40),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_69),
.B1(n_45),
.B2(n_37),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_45),
.A2(n_33),
.B1(n_26),
.B2(n_30),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_33),
.B1(n_30),
.B2(n_25),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_96),
.B1(n_64),
.B2(n_56),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_33),
.B1(n_30),
.B2(n_25),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_41),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_35),
.Y(n_137)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_24),
.B1(n_21),
.B2(n_31),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_24),
.B1(n_31),
.B2(n_42),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_50),
.A2(n_43),
.B1(n_42),
.B2(n_40),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_36),
.B1(n_3),
.B2(n_4),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_44),
.B(n_43),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_52),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_119),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_117),
.B(n_125),
.Y(n_175)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_51),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_121),
.A2(n_139),
.B1(n_110),
.B2(n_4),
.Y(n_160)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_122),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_64),
.B1(n_56),
.B2(n_53),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_123),
.A2(n_127),
.B1(n_128),
.B2(n_134),
.Y(n_177)
);

NAND2x1_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_53),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_110),
.B(n_70),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_89),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_73),
.A2(n_95),
.B1(n_77),
.B2(n_87),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_54),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_7),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_135),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_146),
.C(n_94),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_87),
.A2(n_111),
.B1(n_108),
.B2(n_98),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_35),
.Y(n_135)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_138),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_86),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_18),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_17),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_74),
.B(n_36),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_104),
.B(n_82),
.C(n_94),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_147),
.A2(n_126),
.B(n_120),
.C(n_12),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_144),
.A2(n_104),
.B(n_106),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_124),
.B(n_146),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_117),
.A2(n_111),
.B1(n_108),
.B2(n_98),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_160),
.B1(n_164),
.B2(n_167),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_133),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_155),
.Y(n_178)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_17),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_13),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_146),
.C(n_175),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_125),
.A2(n_106),
.B1(n_4),
.B2(n_6),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_115),
.B(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_112),
.B(n_6),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_112),
.A2(n_106),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_123),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_165),
.B1(n_173),
.B2(n_177),
.Y(n_203)
);

INVx6_ASAP7_75t_SL g170 ( 
.A(n_122),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_13),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_173),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_127),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_134),
.B1(n_133),
.B2(n_129),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g223 ( 
.A1(n_179),
.A2(n_183),
.B(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_177),
.C(n_164),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_114),
.A3(n_143),
.B1(n_130),
.B2(n_116),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_193),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_151),
.A2(n_140),
.B1(n_129),
.B2(n_113),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_170),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_192),
.Y(n_213)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_137),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_195),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_113),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_196),
.A2(n_176),
.B(n_162),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

HAxp5_ASAP7_75t_SL g198 ( 
.A(n_156),
.B(n_142),
.CON(n_198),
.SN(n_198)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_198),
.A2(n_176),
.B(n_149),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_162),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_116),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_167),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_154),
.A2(n_120),
.B1(n_126),
.B2(n_118),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_204),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_160),
.B1(n_174),
.B2(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_161),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_206),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_166),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_212),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_147),
.B(n_152),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_222),
.B(n_225),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_200),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_210),
.B(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_155),
.C(n_169),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_218),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_172),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_176),
.C(n_149),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_226),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_162),
.B(n_179),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_185),
.B(n_193),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_178),
.C(n_186),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_229),
.A2(n_235),
.B(n_209),
.Y(n_252)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_213),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_236),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_223),
.A2(n_202),
.B(n_191),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_211),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_237),
.B(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_189),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_242),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_216),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_243),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_208),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_250),
.C(n_236),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_191),
.B1(n_205),
.B2(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_212),
.B1(n_226),
.B2(n_184),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_249),
.B1(n_253),
.B2(n_231),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_241),
.B1(n_238),
.B2(n_227),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_224),
.C(n_218),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_252),
.A2(n_229),
.B(n_222),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_220),
.B1(n_214),
.B2(n_206),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_230),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_264),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_237),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_258),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_262),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_263),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_239),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_234),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_249),
.B(n_235),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_234),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_267),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_252),
.B(n_255),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_275),
.B(n_254),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_255),
.B1(n_251),
.B2(n_266),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_270),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_251),
.B1(n_247),
.B2(n_248),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_280),
.Y(n_282)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_278),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_267),
.C(n_257),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_281),
.B1(n_271),
.B2(n_190),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_180),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_271),
.B1(n_274),
.B2(n_273),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_285),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_280),
.A2(n_248),
.B1(n_232),
.B2(n_194),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_182),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_204),
.C(n_187),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_287),
.A2(n_282),
.B(n_188),
.Y(n_291)
);

AO21x2_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_282),
.B(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_291),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_288),
.C(n_289),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_202),
.C(n_187),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_202),
.Y(n_295)
);


endmodule