module real_jpeg_7889_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_32, n_33, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_32;
input n_33;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_17;
wire n_21;
wire n_29;
wire n_10;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_0),
.A2(n_3),
.B(n_13),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_SL g26 ( 
.A(n_0),
.B(n_3),
.C(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_19),
.B(n_20),
.Y(n_18)
);

NOR3xp33_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_19),
.C(n_20),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_28),
.B(n_29),
.Y(n_27)
);

NOR3xp33_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_28),
.C(n_29),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_SL g12 ( 
.A(n_7),
.B(n_8),
.C(n_13),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_7),
.A2(n_8),
.B(n_13),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_15),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_14),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_33),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_27),
.B(n_30),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_25),
.B(n_26),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_21),
.B(n_24),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_32),
.Y(n_19)
);


endmodule