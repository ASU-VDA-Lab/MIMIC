module fake_ibex_221_n_2958 (n_151, n_85, n_507, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_8, n_224, n_183, n_508, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_483, n_141, n_487, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_479, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_382, n_502, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_425, n_2958);

input n_151;
input n_85;
input n_507;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_508;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_141;
input n_487;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_479;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_382;
input n_502;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2958;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_523;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1960;
wire n_1723;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_2723;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2879;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_2779;
wire n_521;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_524;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1599;
wire n_712;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_2654;
wire n_2463;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_528;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1845;
wire n_1104;
wire n_1667;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_545;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_961;
wire n_634;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_2862;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_2920;
wire n_604;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_1625;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1348;
wire n_838;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_2945;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1642;
wire n_1455;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_2447;
wire n_2818;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_520;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_2608;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2861;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_2518;
wire n_2784;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1572;
wire n_1635;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_2882;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_543;
wire n_580;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_999;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2931;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_924;
wire n_2937;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2704;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_2754;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_534;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1947;
wire n_1675;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_565;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

BUFx3_ASAP7_75t_L g516 ( 
.A(n_354),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_332),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_411),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_344),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_511),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_219),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_467),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_330),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_68),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_90),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_45),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_227),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_173),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_258),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_217),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_259),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_421),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_141),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_439),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_323),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_215),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_309),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_289),
.Y(n_539)
);

BUFx8_ASAP7_75t_SL g540 ( 
.A(n_184),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_394),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_469),
.Y(n_542)
);

BUFx2_ASAP7_75t_SL g543 ( 
.A(n_353),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_161),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_138),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_222),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_364),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_159),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_193),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_48),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_407),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_388),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_205),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_468),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_201),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_25),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_159),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_503),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_63),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_172),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_192),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_197),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_307),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_498),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_133),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_157),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_395),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_393),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_435),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_370),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_487),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_56),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_249),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_190),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_461),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_197),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_63),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_314),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_259),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_389),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_437),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_134),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_491),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_40),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_161),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_86),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_218),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_432),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_29),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_429),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_10),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_77),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_458),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_390),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_371),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_20),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_338),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_305),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_490),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_131),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_16),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_195),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_53),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_324),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_369),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_333),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_492),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_408),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_392),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_228),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_315),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_463),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_50),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_235),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_418),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_480),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_441),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_325),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_489),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_182),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_273),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_176),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_317),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_241),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_267),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_415),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_292),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_217),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_430),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_287),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_309),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_396),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_423),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_482),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_454),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_252),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_453),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_166),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_227),
.B(n_470),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_177),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_20),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_170),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_501),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_202),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_240),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_331),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_313),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_92),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_6),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_64),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_130),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_499),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_83),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_304),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_361),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_422),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_238),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_145),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_213),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_253),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_505),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_310),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_101),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_452),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_2),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_433),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_78),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_36),
.Y(n_669)
);

CKINVDCx16_ASAP7_75t_R g670 ( 
.A(n_226),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_436),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_420),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_280),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_78),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_229),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_69),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_477),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_8),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_450),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_130),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_274),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_118),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_200),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_464),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_48),
.B(n_384),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_51),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_359),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_502),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_484),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_279),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_152),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_391),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_237),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_224),
.B(n_367),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_497),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_342),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_236),
.Y(n_697)
);

NOR2xp67_ASAP7_75t_L g698 ( 
.A(n_31),
.B(n_425),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_401),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_195),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_479),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_278),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_386),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_146),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_424),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_58),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_64),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_155),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_474),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_68),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_146),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_301),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_69),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_215),
.Y(n_714)
);

BUFx8_ASAP7_75t_SL g715 ( 
.A(n_350),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_300),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_428),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_132),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_488),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_362),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_385),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_223),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_39),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_507),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_45),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_443),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_462),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_465),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_335),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_31),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_96),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_294),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_483),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_506),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_145),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_481),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_281),
.Y(n_737)
);

INVxp33_ASAP7_75t_SL g738 ( 
.A(n_382),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_153),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_11),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_L g741 ( 
.A(n_185),
.B(n_136),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_366),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_273),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_86),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_214),
.Y(n_745)
);

INVxp33_ASAP7_75t_R g746 ( 
.A(n_431),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_306),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_181),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_98),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_357),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_256),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_410),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_88),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_123),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_440),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_129),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_504),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_23),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_13),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_300),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_434),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_358),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_365),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_134),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_444),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_282),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_101),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_376),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_448),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_142),
.Y(n_770)
);

CKINVDCx16_ASAP7_75t_R g771 ( 
.A(n_274),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_58),
.Y(n_772)
);

BUFx10_ASAP7_75t_L g773 ( 
.A(n_473),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_127),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_225),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_216),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_311),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_144),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_89),
.Y(n_779)
);

BUFx10_ASAP7_75t_L g780 ( 
.A(n_486),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_202),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_326),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_363),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_327),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_284),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_107),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_278),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_265),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_339),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_0),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_291),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_92),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_356),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_301),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_51),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_251),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_414),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_180),
.Y(n_798)
);

CKINVDCx14_ASAP7_75t_R g799 ( 
.A(n_514),
.Y(n_799)
);

BUFx10_ASAP7_75t_L g800 ( 
.A(n_216),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_46),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_355),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_131),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_205),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_302),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_307),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_485),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_251),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_77),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_256),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_165),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_186),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_85),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_184),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_455),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_478),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_296),
.Y(n_817)
);

CKINVDCx14_ASAP7_75t_R g818 ( 
.A(n_85),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_165),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_88),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_345),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_378),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_114),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_8),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_0),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_509),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_406),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_214),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_257),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_117),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_40),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_315),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_26),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_65),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_258),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_267),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_79),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_445),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_397),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_368),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_387),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_177),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_66),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_442),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_95),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_303),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_67),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_229),
.Y(n_848)
);

BUFx8_ASAP7_75t_SL g849 ( 
.A(n_404),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_360),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_228),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_340),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_230),
.Y(n_853)
);

INVx1_ASAP7_75t_SL g854 ( 
.A(n_3),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_281),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_400),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_475),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_167),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_210),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_438),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_493),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_377),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_24),
.Y(n_863)
);

CKINVDCx14_ASAP7_75t_R g864 ( 
.A(n_351),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_818),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_673),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_591),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_519),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_527),
.B(n_1),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_785),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_519),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_519),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_673),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_519),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_673),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_534),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_670),
.B(n_1),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_534),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_609),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_618),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_618),
.Y(n_881)
);

BUFx12f_ASAP7_75t_L g882 ( 
.A(n_591),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_578),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_618),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_618),
.Y(n_885)
);

CKINVDCx11_ASAP7_75t_R g886 ( 
.A(n_536),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_654),
.B(n_2),
.Y(n_887)
);

OAI22x1_ASAP7_75t_L g888 ( 
.A1(n_654),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_688),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_578),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_689),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_624),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_591),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_789),
.Y(n_894)
);

INVx5_ASAP7_75t_L g895 ( 
.A(n_620),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_689),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_624),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_689),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_620),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_680),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_602),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_680),
.B(n_4),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_779),
.B(n_5),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_630),
.Y(n_904)
);

INVx6_ASAP7_75t_L g905 ( 
.A(n_620),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_630),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_800),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_719),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_779),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_602),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_800),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_719),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_706),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_706),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_689),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_713),
.Y(n_916)
);

AND2x6_ASAP7_75t_L g917 ( 
.A(n_516),
.B(n_665),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_808),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_862),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_862),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_540),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_566),
.Y(n_922)
);

BUFx12f_ASAP7_75t_L g923 ( 
.A(n_733),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_808),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_566),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_809),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_764),
.B(n_771),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_733),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_733),
.Y(n_929)
);

OAI22x1_ASAP7_75t_SL g930 ( 
.A1(n_536),
.A2(n_9),
.B1(n_6),
.B2(n_7),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_566),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_809),
.Y(n_932)
);

OA21x2_ASAP7_75t_L g933 ( 
.A1(n_517),
.A2(n_318),
.B(n_316),
.Y(n_933)
);

BUFx12f_ASAP7_75t_L g934 ( 
.A(n_773),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_516),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_567),
.B(n_7),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_715),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_829),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_566),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_715),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_567),
.B(n_9),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_607),
.B(n_10),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_608),
.B(n_11),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_829),
.B(n_539),
.Y(n_944)
);

OAI22x1_ASAP7_75t_SL g945 ( 
.A1(n_549),
.A2(n_14),
.B1(n_12),
.B2(n_13),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_773),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_608),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_522),
.A2(n_320),
.B(n_319),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_725),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_665),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_539),
.B(n_12),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_695),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_540),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_849),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_695),
.Y(n_955)
);

AND2x6_ASAP7_75t_L g956 ( 
.A(n_736),
.B(n_321),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_561),
.Y(n_957)
);

BUFx12f_ASAP7_75t_L g958 ( 
.A(n_773),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_780),
.Y(n_959)
);

AND2x6_ASAP7_75t_L g960 ( 
.A(n_736),
.B(n_322),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_780),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_561),
.Y(n_962)
);

OA21x2_ASAP7_75t_L g963 ( 
.A1(n_538),
.A2(n_329),
.B(n_328),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_725),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_725),
.Y(n_965)
);

OAI22xp33_ASAP7_75t_SL g966 ( 
.A1(n_905),
.A2(n_524),
.B1(n_528),
.B2(n_521),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_937),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_865),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_873),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_937),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_940),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_954),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_921),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_873),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_921),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_953),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_953),
.Y(n_977)
);

NAND2xp33_ASAP7_75t_R g978 ( 
.A(n_869),
.B(n_738),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_886),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_886),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_882),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_923),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_865),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_R g984 ( 
.A(n_923),
.B(n_799),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_928),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_875),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_R g987 ( 
.A(n_928),
.B(n_864),
.Y(n_987)
);

CKINVDCx16_ASAP7_75t_R g988 ( 
.A(n_934),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_934),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_944),
.Y(n_990)
);

BUFx10_ASAP7_75t_L g991 ( 
.A(n_905),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_944),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_958),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_927),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_958),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_870),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_879),
.A2(n_598),
.B1(n_617),
.B2(n_571),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_877),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_867),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_929),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_875),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_887),
.Y(n_1002)
);

NAND2xp33_ASAP7_75t_SL g1003 ( 
.A(n_929),
.B(n_571),
.Y(n_1003)
);

OAI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_888),
.A2(n_560),
.B1(n_590),
.B2(n_549),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_905),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_911),
.B(n_598),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_959),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_959),
.Y(n_1008)
);

AO21x2_ASAP7_75t_L g1009 ( 
.A1(n_948),
.A2(n_551),
.B(n_541),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_914),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_944),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_926),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_932),
.Y(n_1013)
);

BUFx10_ASAP7_75t_L g1014 ( 
.A(n_887),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_893),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_893),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_893),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_893),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_895),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_887),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_902),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_895),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_895),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_868),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_868),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_899),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_868),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_899),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_899),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_899),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_946),
.B(n_858),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_946),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_902),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_946),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_935),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_868),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_911),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_883),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_871),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_935),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_902),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_903),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_955),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_961),
.B(n_529),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_907),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_890),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_950),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_889),
.B(n_589),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_890),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_901),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_951),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_901),
.B(n_780),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_913),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_952),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_951),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_952),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_913),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_924),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_871),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_951),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_924),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_866),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_900),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_894),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_909),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_936),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_930),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_941),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_942),
.Y(n_1069)
);

BUFx10_ASAP7_75t_L g1070 ( 
.A(n_910),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_917),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_945),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_876),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_956),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_947),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_876),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_947),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_943),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_878),
.Y(n_1079)
);

BUFx10_ASAP7_75t_L g1080 ( 
.A(n_916),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_918),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_938),
.B(n_564),
.Y(n_1082)
);

NAND2xp33_ASAP7_75t_R g1083 ( 
.A(n_933),
.B(n_531),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_957),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_962),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_871),
.Y(n_1086)
);

BUFx2_ASAP7_75t_L g1087 ( 
.A(n_892),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_892),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_897),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_871),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_897),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_904),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_904),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_906),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_906),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_908),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_908),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_912),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_919),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_R g1100 ( 
.A(n_917),
.B(n_619),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_956),
.A2(n_653),
.B1(n_696),
.B2(n_619),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_919),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_920),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_872),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_920),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_917),
.Y(n_1106)
);

INVxp33_ASAP7_75t_L g1107 ( 
.A(n_922),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_917),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_965),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_956),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_872),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_922),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_922),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_R g1114 ( 
.A(n_960),
.B(n_721),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_922),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_960),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_960),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_R g1118 ( 
.A(n_960),
.B(n_721),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_925),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_925),
.Y(n_1120)
);

CKINVDCx16_ASAP7_75t_R g1121 ( 
.A(n_925),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_925),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_931),
.Y(n_1123)
);

CKINVDCx16_ASAP7_75t_R g1124 ( 
.A(n_931),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_931),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_931),
.B(n_660),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_939),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_933),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_939),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_939),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_939),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_965),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_949),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_965),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_965),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_949),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1066),
.B(n_634),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_991),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1078),
.B(n_518),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1089),
.B(n_520),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1000),
.B(n_662),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1096),
.B(n_523),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1014),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_1007),
.B(n_552),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1035),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_968),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1040),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1008),
.B(n_600),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1005),
.B(n_752),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1091),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_986),
.B(n_763),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1046),
.B(n_1001),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1091),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_999),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_L g1155 ( 
.A(n_1110),
.B(n_532),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1043),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1079),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1102),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1097),
.B(n_535),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1074),
.B(n_542),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1044),
.B(n_765),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_L g1162 ( 
.A(n_1083),
.B(n_963),
.C(n_933),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1098),
.B(n_547),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_988),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1103),
.B(n_554),
.Y(n_1165)
);

INVxp33_ASAP7_75t_L g1166 ( 
.A(n_1006),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1071),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_SL g1168 ( 
.A(n_991),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1079),
.Y(n_1169)
);

AND2x6_ASAP7_75t_SL g1170 ( 
.A(n_980),
.B(n_746),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1099),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_1010),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1105),
.B(n_558),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1052),
.B(n_568),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1102),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1063),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1065),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1087),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1070),
.B(n_569),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1070),
.B(n_570),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_L g1181 ( 
.A(n_1004),
.B(n_775),
.C(n_710),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_990),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1099),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1073),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1076),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1083),
.B(n_963),
.C(n_580),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1037),
.B(n_815),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1080),
.B(n_581),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1075),
.B(n_583),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_992),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1011),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1014),
.B(n_595),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1126),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1126),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1077),
.B(n_596),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1048),
.B(n_605),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_996),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_969),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1049),
.A2(n_755),
.B1(n_757),
.B2(n_734),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_974),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1048),
.B(n_610),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1047),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_997),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1042),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_L g1205 ( 
.A(n_1004),
.B(n_743),
.C(n_686),
.Y(n_1205)
);

NAND2xp33_ASAP7_75t_L g1206 ( 
.A(n_1117),
.B(n_613),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1042),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1054),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1002),
.A2(n_526),
.B1(n_530),
.B2(n_525),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1056),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1045),
.B(n_627),
.Y(n_1211)
);

NAND3xp33_ASAP7_75t_L g1212 ( 
.A(n_1020),
.B(n_963),
.C(n_587),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1021),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1071),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1033),
.B(n_635),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1041),
.B(n_636),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1088),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1116),
.Y(n_1218)
);

INVxp33_ASAP7_75t_L g1219 ( 
.A(n_1006),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1051),
.B(n_638),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1055),
.B(n_575),
.Y(n_1221)
);

INVx6_ASAP7_75t_L g1222 ( 
.A(n_1121),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_1114),
.B(n_644),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_1012),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1114),
.B(n_647),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1013),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1060),
.B(n_594),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1062),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1081),
.B(n_606),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1094),
.Y(n_1230)
);

BUFx5_ASAP7_75t_L g1231 ( 
.A(n_1109),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1031),
.B(n_656),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1050),
.B(n_657),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1118),
.B(n_667),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1053),
.B(n_672),
.Y(n_1235)
);

BUFx5_ASAP7_75t_L g1236 ( 
.A(n_1112),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1118),
.B(n_1100),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1057),
.B(n_677),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1058),
.B(n_684),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1095),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1061),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1100),
.B(n_692),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_SL g1243 ( 
.A(n_1106),
.B(n_734),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1092),
.A2(n_757),
.B1(n_802),
.B2(n_755),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1108),
.B(n_701),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1082),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1009),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1124),
.B(n_703),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1128),
.B(n_633),
.C(n_616),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_966),
.B(n_705),
.Y(n_1250)
);

NOR3xp33_ASAP7_75t_L g1251 ( 
.A(n_1003),
.B(n_854),
.C(n_747),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_973),
.Y(n_1252)
);

NOR2xp67_ASAP7_75t_L g1253 ( 
.A(n_981),
.B(n_640),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_984),
.B(n_709),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1093),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1009),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_984),
.B(n_724),
.Y(n_1257)
);

NAND2xp33_ASAP7_75t_L g1258 ( 
.A(n_987),
.B(n_727),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1015),
.B(n_750),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1016),
.B(n_761),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1068),
.B(n_762),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1122),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1017),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1018),
.Y(n_1264)
);

NAND2xp33_ASAP7_75t_L g1265 ( 
.A(n_987),
.B(n_768),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_994),
.B(n_741),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1123),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1019),
.B(n_671),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1022),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1026),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1023),
.B(n_802),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1028),
.B(n_769),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1029),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_L g1274 ( 
.A(n_1101),
.B(n_687),
.C(n_679),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1030),
.B(n_782),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1069),
.B(n_783),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_983),
.B(n_784),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1032),
.B(n_793),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1034),
.B(n_807),
.Y(n_1279)
);

NOR3xp33_ASAP7_75t_L g1280 ( 
.A(n_1067),
.B(n_545),
.C(n_544),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_982),
.B(n_985),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1084),
.B(n_816),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1125),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1085),
.B(n_826),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_989),
.B(n_827),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1064),
.B(n_838),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_993),
.B(n_546),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_R g1288 ( 
.A(n_995),
.B(n_821),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_976),
.B(n_839),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1127),
.Y(n_1290)
);

AOI221xp5_ASAP7_75t_L g1291 ( 
.A1(n_977),
.A2(n_548),
.B1(n_555),
.B2(n_537),
.C(n_533),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1130),
.Y(n_1292)
);

AND2x4_ASAP7_75t_L g1293 ( 
.A(n_967),
.B(n_821),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1131),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_998),
.B(n_840),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_971),
.B(n_972),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1133),
.B(n_844),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1136),
.B(n_856),
.Y(n_1298)
);

NAND2xp33_ASAP7_75t_L g1299 ( 
.A(n_970),
.B(n_857),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1115),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1107),
.B(n_860),
.Y(n_1301)
);

XNOR2x2_ASAP7_75t_L g1302 ( 
.A(n_979),
.B(n_685),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_975),
.B(n_550),
.Y(n_1303)
);

CKINVDCx16_ASAP7_75t_R g1304 ( 
.A(n_978),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_978),
.B(n_861),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1120),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1072),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1129),
.B(n_543),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1132),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1059),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1059),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1134),
.B(n_699),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1135),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1113),
.B(n_553),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1119),
.B(n_556),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1024),
.A2(n_841),
.B1(n_562),
.B2(n_563),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1059),
.B(n_720),
.C(n_717),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1024),
.B(n_557),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1025),
.B(n_726),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1090),
.B(n_728),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1090),
.B(n_729),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1027),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1027),
.B(n_742),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1090),
.B(n_797),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1090),
.B(n_822),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1036),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1036),
.A2(n_572),
.B1(n_574),
.B2(n_559),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1039),
.B(n_565),
.Y(n_1328)
);

NOR2xp67_ASAP7_75t_L g1329 ( 
.A(n_1039),
.B(n_15),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1104),
.B(n_850),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1086),
.B(n_573),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1086),
.B(n_852),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1104),
.B(n_660),
.Y(n_1333)
);

XNOR2x2_ASAP7_75t_L g1334 ( 
.A(n_1111),
.B(n_560),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1111),
.B(n_725),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1078),
.B(n_716),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1091),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_999),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_L g1339 ( 
.A(n_1083),
.B(n_582),
.C(n_577),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1066),
.B(n_576),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1091),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1071),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1078),
.B(n_716),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1066),
.B(n_845),
.Y(n_1344)
);

NAND2xp33_ASAP7_75t_L g1345 ( 
.A(n_1110),
.B(n_841),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_997),
.B(n_845),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1091),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1091),
.Y(n_1348)
);

INVxp33_ASAP7_75t_L g1349 ( 
.A(n_1006),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1038),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1091),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1000),
.B(n_579),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1066),
.B(n_593),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1091),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_L g1355 ( 
.A(n_1083),
.B(n_585),
.C(n_584),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1091),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1002),
.A2(n_588),
.B(n_592),
.C(n_586),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1066),
.B(n_599),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1000),
.B(n_604),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1078),
.B(n_694),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1066),
.B(n_611),
.Y(n_1361)
);

INVxp33_ASAP7_75t_L g1362 ( 
.A(n_1006),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_996),
.B(n_614),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1091),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1002),
.A2(n_612),
.B(n_615),
.C(n_603),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1066),
.B(n_621),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1035),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1035),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1035),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1035),
.Y(n_1370)
);

INVx5_ASAP7_75t_L g1371 ( 
.A(n_1014),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1078),
.B(n_698),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1035),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1000),
.B(n_622),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1078),
.B(n_623),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1091),
.Y(n_1376)
);

INVx5_ASAP7_75t_L g1377 ( 
.A(n_1222),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1222),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1207),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1152),
.B(n_628),
.Y(n_1380)
);

AND2x6_ASAP7_75t_L g1381 ( 
.A(n_1218),
.B(n_625),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1339),
.A2(n_597),
.B1(n_601),
.B2(n_590),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1152),
.B(n_629),
.Y(n_1383)
);

BUFx8_ASAP7_75t_L g1384 ( 
.A(n_1168),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1213),
.A2(n_632),
.B(n_650),
.C(n_626),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1371),
.B(n_631),
.Y(n_1386)
);

INVx5_ASAP7_75t_L g1387 ( 
.A(n_1371),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1150),
.B(n_637),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1350),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1176),
.A2(n_652),
.B(n_655),
.C(n_651),
.Y(n_1390)
);

AND2x6_ASAP7_75t_SL g1391 ( 
.A(n_1170),
.B(n_1266),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1204),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1153),
.B(n_639),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1158),
.B(n_641),
.Y(n_1394)
);

O2A1O1Ixp5_ASAP7_75t_L g1395 ( 
.A1(n_1162),
.A2(n_1186),
.B(n_1256),
.C(n_1247),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1350),
.Y(n_1396)
);

AND2x2_ASAP7_75t_SL g1397 ( 
.A(n_1243),
.B(n_849),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1167),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1339),
.A2(n_1355),
.B1(n_1274),
.B2(n_1249),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1146),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1355),
.A2(n_601),
.B1(n_646),
.B2(n_597),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1274),
.A2(n_658),
.B1(n_666),
.B2(n_646),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1371),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1204),
.Y(n_1404)
);

AO22x1_ASAP7_75t_L g1405 ( 
.A1(n_1293),
.A2(n_674),
.B1(n_676),
.B2(n_666),
.Y(n_1405)
);

NOR3xp33_ASAP7_75t_SL g1406 ( 
.A(n_1307),
.B(n_643),
.C(n_642),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1167),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1371),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1175),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1295),
.B(n_1286),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1282),
.B(n_674),
.Y(n_1411)
);

INVx2_ASAP7_75t_SL g1412 ( 
.A(n_1138),
.Y(n_1412)
);

NOR3xp33_ASAP7_75t_SL g1413 ( 
.A(n_1164),
.B(n_648),
.C(n_645),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1288),
.Y(n_1414)
);

NOR2x1_ASAP7_75t_R g1415 ( 
.A(n_1293),
.B(n_649),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1337),
.B(n_659),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1341),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1347),
.B(n_663),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1252),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1241),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1284),
.B(n_676),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1244),
.B(n_1199),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1143),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1348),
.B(n_664),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1351),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1154),
.Y(n_1426)
);

NAND2xp33_ASAP7_75t_SL g1427 ( 
.A(n_1168),
.B(n_683),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1217),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1375),
.B(n_683),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1249),
.A2(n_693),
.B1(n_697),
.B2(n_690),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1354),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1338),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1203),
.A2(n_693),
.B1(n_697),
.B2(n_690),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1143),
.B(n_669),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1356),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1363),
.B(n_700),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1262),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1172),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1364),
.Y(n_1439)
);

AND3x2_ASAP7_75t_SL g1440 ( 
.A(n_1271),
.B(n_704),
.C(n_700),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1197),
.B(n_675),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1376),
.B(n_678),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1177),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1224),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1263),
.B(n_661),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1167),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1304),
.A2(n_753),
.B1(n_772),
.B2(n_704),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1346),
.A2(n_772),
.B1(n_776),
.B2(n_753),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1264),
.B(n_668),
.Y(n_1449)
);

AND2x4_ASAP7_75t_L g1450 ( 
.A(n_1269),
.B(n_681),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1137),
.B(n_682),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1182),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1137),
.B(n_691),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1193),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_R g1455 ( 
.A(n_1243),
.B(n_776),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1344),
.B(n_707),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1270),
.B(n_702),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1190),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1344),
.B(n_708),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1340),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1346),
.B(n_781),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1358),
.B(n_1209),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1191),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1228),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1198),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1305),
.B(n_781),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1194),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1226),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_1353),
.Y(n_1469)
);

AND2x6_ASAP7_75t_L g1470 ( 
.A(n_1218),
.B(n_711),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1262),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1230),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1273),
.B(n_714),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1346),
.A2(n_796),
.B1(n_825),
.B2(n_791),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1178),
.B(n_723),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1328),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1214),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1334),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1331),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1361),
.B(n_712),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1262),
.B(n_1294),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1267),
.B(n_718),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1345),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1267),
.Y(n_1484)
);

INVx4_ASAP7_75t_L g1485 ( 
.A(n_1267),
.Y(n_1485)
);

NOR2x2_ASAP7_75t_L g1486 ( 
.A(n_1266),
.B(n_791),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1200),
.Y(n_1487)
);

NOR2x2_ASAP7_75t_L g1488 ( 
.A(n_1266),
.B(n_1302),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1145),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1366),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1296),
.B(n_732),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1287),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1161),
.B(n_722),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1151),
.B(n_730),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1357),
.B(n_731),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1294),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1214),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1277),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1365),
.B(n_739),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1147),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_SL g1501 ( 
.A(n_1166),
.B(n_796),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1303),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1214),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1221),
.A2(n_737),
.B(n_744),
.C(n_735),
.Y(n_1504)
);

OAI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1221),
.A2(n_825),
.B1(n_751),
.B2(n_758),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1157),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1342),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1316),
.A2(n_745),
.B1(n_748),
.B2(n_740),
.Y(n_1508)
);

NOR2x2_ASAP7_75t_L g1509 ( 
.A(n_1261),
.B(n_754),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1169),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1174),
.B(n_756),
.Y(n_1511)
);

AND2x6_ASAP7_75t_L g1512 ( 
.A(n_1246),
.B(n_749),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1156),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_SL g1514 ( 
.A(n_1255),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1336),
.B(n_759),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1276),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1179),
.B(n_760),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1171),
.Y(n_1518)
);

AND2x6_ASAP7_75t_L g1519 ( 
.A(n_1294),
.B(n_766),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1181),
.A2(n_786),
.B1(n_787),
.B2(n_777),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1233),
.B(n_767),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1205),
.A2(n_795),
.B1(n_801),
.B2(n_790),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1227),
.A2(n_817),
.B1(n_820),
.B2(n_804),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1248),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1281),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1183),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1240),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1367),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1279),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1180),
.B(n_770),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1227),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1229),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1229),
.Y(n_1533)
);

NAND3xp33_ASAP7_75t_SL g1534 ( 
.A(n_1251),
.B(n_778),
.C(n_774),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1162),
.A2(n_824),
.B(n_823),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1311),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1368),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1343),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1238),
.B(n_788),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1139),
.B(n_831),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1291),
.A2(n_1327),
.B1(n_1184),
.B2(n_1185),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1188),
.B(n_792),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1311),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1292),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1369),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1370),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1373),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_L g1548 ( 
.A(n_1186),
.B(n_794),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1202),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1140),
.B(n_1142),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1219),
.A2(n_803),
.B1(n_805),
.B2(n_798),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_SL g1552 ( 
.A(n_1211),
.B(n_806),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1159),
.B(n_810),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1292),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1285),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1235),
.B(n_811),
.Y(n_1556)
);

O2A1O1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1250),
.A2(n_846),
.B(n_848),
.C(n_842),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1163),
.B(n_812),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1253),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1192),
.B(n_851),
.Y(n_1560)
);

AND3x2_ASAP7_75t_SL g1561 ( 
.A(n_1280),
.B(n_814),
.C(n_813),
.Y(n_1561)
);

XOR2x2_ASAP7_75t_L g1562 ( 
.A(n_1360),
.B(n_14),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1208),
.A2(n_859),
.B1(n_863),
.B2(n_853),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1210),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1352),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1359),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1319),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1319),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1374),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1333),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1289),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1165),
.B(n_819),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1323),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1212),
.A2(n_830),
.B(n_832),
.C(n_828),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1283),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1323),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1215),
.A2(n_834),
.B1(n_835),
.B2(n_833),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1239),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1216),
.A2(n_837),
.B1(n_843),
.B2(n_836),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1332),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1173),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1144),
.B(n_847),
.Y(n_1582)
);

INVx5_ASAP7_75t_L g1583 ( 
.A(n_1290),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1318),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1314),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1254),
.B(n_855),
.Y(n_1586)
);

NOR2x2_ASAP7_75t_L g1587 ( 
.A(n_1299),
.B(n_16),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1220),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1148),
.B(n_17),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1189),
.B(n_17),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1195),
.B(n_18),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_SL g1592 ( 
.A1(n_1349),
.A2(n_21),
.B1(n_18),
.B2(n_19),
.Y(n_1592)
);

CKINVDCx6p67_ASAP7_75t_R g1593 ( 
.A(n_1257),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1187),
.B(n_19),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1196),
.B(n_22),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1362),
.B(n_964),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1315),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1201),
.B(n_1141),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1268),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1372),
.B(n_964),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1232),
.B(n_23),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1149),
.B(n_24),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1329),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1308),
.Y(n_1604)
);

AO22x1_ASAP7_75t_L g1605 ( 
.A1(n_1297),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1160),
.B(n_27),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1231),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1320),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1325),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1223),
.B(n_28),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1225),
.B(n_28),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1275),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1259),
.Y(n_1613)
);

AOI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1234),
.A2(n_880),
.B1(n_881),
.B2(n_874),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1312),
.A2(n_880),
.B1(n_881),
.B2(n_874),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1330),
.Y(n_1616)
);

BUFx12f_ASAP7_75t_L g1617 ( 
.A(n_1258),
.Y(n_1617)
);

AND2x2_ASAP7_75t_SL g1618 ( 
.A(n_1265),
.B(n_29),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1321),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1260),
.B(n_30),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1272),
.B(n_30),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1237),
.A2(n_884),
.B1(n_885),
.B2(n_881),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1301),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1324),
.Y(n_1624)
);

NOR3xp33_ASAP7_75t_SL g1625 ( 
.A(n_1278),
.B(n_32),
.C(n_33),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1242),
.B(n_32),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1310),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1298),
.B(n_33),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1245),
.B(n_34),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1155),
.B(n_34),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1317),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1310),
.Y(n_1632)
);

A2O1A1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1206),
.A2(n_885),
.B(n_891),
.C(n_884),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1313),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1634)
);

OR2x6_ASAP7_75t_L g1635 ( 
.A(n_1335),
.B(n_37),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1326),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1236),
.B(n_38),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1300),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1306),
.Y(n_1639)
);

NAND3xp33_ASAP7_75t_SL g1640 ( 
.A(n_1309),
.B(n_38),
.C(n_39),
.Y(n_1640)
);

AND3x2_ASAP7_75t_SL g1641 ( 
.A(n_1322),
.B(n_41),
.C(n_42),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1236),
.B(n_41),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1339),
.A2(n_915),
.B1(n_885),
.B2(n_891),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1167),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1532),
.B(n_42),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1387),
.B(n_884),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1448),
.A2(n_46),
.B1(n_43),
.B2(n_44),
.Y(n_1647)
);

OR2x6_ASAP7_75t_L g1648 ( 
.A(n_1405),
.B(n_43),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1536),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1443),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1409),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1395),
.A2(n_885),
.B(n_884),
.Y(n_1652)
);

BUFx12f_ASAP7_75t_L g1653 ( 
.A(n_1384),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1550),
.A2(n_1548),
.B(n_1533),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_SL g1655 ( 
.A1(n_1574),
.A2(n_336),
.B(n_337),
.C(n_334),
.Y(n_1655)
);

AO21x2_ASAP7_75t_L g1656 ( 
.A1(n_1535),
.A2(n_896),
.B(n_891),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1436),
.B(n_1422),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1417),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1387),
.B(n_896),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1531),
.A2(n_1599),
.B1(n_1568),
.B2(n_1573),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1462),
.B(n_47),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1425),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1387),
.B(n_47),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1567),
.A2(n_898),
.B1(n_915),
.B2(n_896),
.Y(n_1664)
);

AO21x1_ASAP7_75t_L g1665 ( 
.A1(n_1637),
.A2(n_1642),
.B(n_1643),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1576),
.A2(n_1580),
.B(n_1588),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1466),
.B(n_49),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1431),
.B(n_49),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1411),
.B(n_50),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1435),
.B(n_52),
.Y(n_1670)
);

INVx3_ASAP7_75t_L g1671 ( 
.A(n_1403),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1384),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1391),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1439),
.B(n_1554),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1468),
.B(n_898),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1448),
.A2(n_52),
.B(n_53),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1536),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1455),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1618),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_R g1680 ( 
.A(n_1427),
.B(n_54),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1598),
.B(n_55),
.C(n_57),
.Y(n_1681)
);

O2A1O1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1504),
.A2(n_60),
.B(n_57),
.C(n_59),
.Y(n_1682)
);

AND2x4_ASAP7_75t_SL g1683 ( 
.A(n_1444),
.B(n_59),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1400),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1433),
.B(n_60),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1472),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1397),
.B(n_1552),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1389),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1464),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_R g1690 ( 
.A(n_1419),
.B(n_61),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1476),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1390),
.A2(n_1385),
.B(n_1505),
.C(n_1469),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1529),
.B(n_62),
.Y(n_1693)
);

O2A1O1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1460),
.A2(n_66),
.B(n_62),
.C(n_65),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1420),
.B(n_67),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_R g1696 ( 
.A(n_1501),
.B(n_70),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1541),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1402),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.C(n_74),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1410),
.B(n_73),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1403),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1479),
.B(n_74),
.Y(n_1701)
);

BUFx4f_ASAP7_75t_L g1702 ( 
.A(n_1617),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1421),
.A2(n_79),
.B1(n_75),
.B2(n_76),
.C(n_80),
.Y(n_1703)
);

HB1xp67_ASAP7_75t_L g1704 ( 
.A(n_1396),
.Y(n_1704)
);

AOI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1584),
.A2(n_343),
.B(n_341),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1490),
.B(n_75),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1597),
.A2(n_347),
.B(n_346),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1452),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1428),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1461),
.B(n_76),
.Y(n_1710)
);

INVx4_ASAP7_75t_L g1711 ( 
.A(n_1377),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1458),
.Y(n_1712)
);

A2O1A1Ixp33_ASAP7_75t_SL g1713 ( 
.A1(n_1539),
.A2(n_349),
.B(n_352),
.C(n_348),
.Y(n_1713)
);

BUFx4f_ASAP7_75t_L g1714 ( 
.A(n_1519),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1541),
.B(n_80),
.Y(n_1715)
);

INVx5_ASAP7_75t_L g1716 ( 
.A(n_1519),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1609),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1474),
.B(n_1382),
.Y(n_1718)
);

NOR3xp33_ASAP7_75t_L g1719 ( 
.A(n_1498),
.B(n_81),
.C(n_82),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1380),
.B(n_84),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1429),
.A2(n_89),
.B1(n_84),
.B2(n_87),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1612),
.B(n_87),
.Y(n_1722)
);

INVx5_ASAP7_75t_L g1723 ( 
.A(n_1519),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1543),
.A2(n_1530),
.B(n_1517),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1383),
.B(n_91),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1519),
.Y(n_1726)
);

CKINVDCx14_ASAP7_75t_R g1727 ( 
.A(n_1447),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1463),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1542),
.A2(n_373),
.B(n_372),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1492),
.B(n_91),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1438),
.B(n_93),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1570),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1613),
.B(n_93),
.Y(n_1733)
);

NOR3xp33_ASAP7_75t_L g1734 ( 
.A(n_1566),
.B(n_94),
.C(n_95),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1549),
.Y(n_1735)
);

OR2x6_ASAP7_75t_L g1736 ( 
.A(n_1414),
.B(n_1426),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1379),
.Y(n_1737)
);

A2O1A1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1616),
.A2(n_1557),
.B(n_1595),
.C(n_1399),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1553),
.A2(n_375),
.B(n_374),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1631),
.A2(n_380),
.B(n_379),
.Y(n_1740)
);

INVx3_ASAP7_75t_SL g1741 ( 
.A(n_1486),
.Y(n_1741)
);

BUFx12f_ASAP7_75t_L g1742 ( 
.A(n_1432),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1558),
.A2(n_383),
.B(n_381),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1378),
.B(n_94),
.Y(n_1744)
);

CKINVDCx20_ASAP7_75t_R g1745 ( 
.A(n_1377),
.Y(n_1745)
);

BUFx2_ASAP7_75t_L g1746 ( 
.A(n_1381),
.Y(n_1746)
);

A2O1A1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1590),
.A2(n_100),
.B(n_97),
.C(n_99),
.Y(n_1747)
);

OAI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1483),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1581),
.B(n_1523),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1551),
.B(n_102),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1527),
.B(n_103),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1523),
.B(n_104),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1412),
.B(n_104),
.Y(n_1753)
);

AO32x1_ASAP7_75t_L g1754 ( 
.A1(n_1594),
.A2(n_107),
.A3(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1636),
.A2(n_399),
.B(n_398),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_SL g1756 ( 
.A(n_1607),
.B(n_105),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1398),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1474),
.A2(n_109),
.B1(n_106),
.B2(n_108),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1398),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1569),
.B(n_109),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1478),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_1761)
);

A2O1A1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1591),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1398),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1475),
.B(n_113),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1638),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1407),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1511),
.A2(n_403),
.B(n_402),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1639),
.A2(n_409),
.B(n_405),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1564),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1377),
.Y(n_1770)
);

INVx4_ASAP7_75t_L g1771 ( 
.A(n_1485),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1524),
.B(n_119),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1522),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1564),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1585),
.B(n_1575),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1381),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1522),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1415),
.B(n_124),
.Y(n_1778)
);

BUFx12f_ASAP7_75t_L g1779 ( 
.A(n_1525),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1382),
.B(n_125),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1475),
.B(n_126),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1451),
.B(n_126),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1437),
.Y(n_1783)
);

AO32x1_ASAP7_75t_L g1784 ( 
.A1(n_1603),
.A2(n_127),
.A3(n_128),
.B1(n_129),
.B2(n_132),
.Y(n_1784)
);

AOI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1480),
.A2(n_413),
.B(n_412),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1471),
.Y(n_1786)
);

NAND2x1p5_ASAP7_75t_L g1787 ( 
.A(n_1484),
.B(n_128),
.Y(n_1787)
);

BUFx4f_ASAP7_75t_L g1788 ( 
.A(n_1593),
.Y(n_1788)
);

AOI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1520),
.A2(n_136),
.B1(n_133),
.B2(n_135),
.Y(n_1789)
);

INVxp67_ASAP7_75t_SL g1790 ( 
.A(n_1433),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1456),
.A2(n_1459),
.B(n_1601),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1607),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1508),
.B(n_135),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1415),
.B(n_137),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1453),
.B(n_137),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1520),
.B(n_138),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1441),
.B(n_139),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1485),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1540),
.B(n_139),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_1571),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1540),
.B(n_140),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1430),
.B(n_1401),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1578),
.B(n_140),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1623),
.B(n_141),
.Y(n_1804)
);

INVx5_ASAP7_75t_L g1805 ( 
.A(n_1381),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1445),
.A2(n_147),
.B1(n_143),
.B2(n_144),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1445),
.B(n_143),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1629),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_1808)
);

O2A1O1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1495),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_1809)
);

O2A1O1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1499),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1586),
.B(n_151),
.Y(n_1811)
);

OAI22x1_ASAP7_75t_L g1812 ( 
.A1(n_1440),
.A2(n_1587),
.B1(n_1491),
.B2(n_1641),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1408),
.B(n_153),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1454),
.Y(n_1814)
);

A2O1A1Ixp33_ASAP7_75t_L g1815 ( 
.A1(n_1628),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_1815)
);

CKINVDCx16_ASAP7_75t_R g1816 ( 
.A(n_1514),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_1381),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1572),
.A2(n_417),
.B(n_416),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1537),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_1407),
.Y(n_1820)
);

O2A1O1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1589),
.A2(n_157),
.B(n_154),
.C(n_156),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1407),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1521),
.B(n_158),
.Y(n_1823)
);

AO32x2_ASAP7_75t_L g1824 ( 
.A1(n_1634),
.A2(n_158),
.A3(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1545),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1423),
.B(n_160),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1565),
.B(n_162),
.Y(n_1827)
);

BUFx10_ASAP7_75t_L g1828 ( 
.A(n_1514),
.Y(n_1828)
);

OAI22x1_ASAP7_75t_L g1829 ( 
.A1(n_1516),
.A2(n_166),
.B1(n_163),
.B2(n_164),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1556),
.B(n_164),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1577),
.B(n_167),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1467),
.Y(n_1832)
);

CKINVDCx8_ASAP7_75t_R g1833 ( 
.A(n_1586),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1413),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1465),
.Y(n_1835)
);

NOR2xp67_ASAP7_75t_L g1836 ( 
.A(n_1640),
.B(n_419),
.Y(n_1836)
);

NOR3xp33_ASAP7_75t_L g1837 ( 
.A(n_1534),
.B(n_168),
.C(n_169),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1449),
.B(n_169),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1577),
.B(n_170),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1449),
.B(n_171),
.Y(n_1840)
);

CKINVDCx8_ASAP7_75t_R g1841 ( 
.A(n_1470),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1547),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1579),
.B(n_171),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1446),
.Y(n_1844)
);

A2O1A1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1620),
.A2(n_172),
.B(n_173),
.C(n_174),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1487),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1450),
.B(n_174),
.Y(n_1847)
);

A2O1A1Ixp33_ASAP7_75t_L g1848 ( 
.A1(n_1621),
.A2(n_175),
.B(n_176),
.C(n_178),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1450),
.B(n_1457),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1579),
.B(n_175),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1489),
.A2(n_427),
.B(n_426),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_SL g1852 ( 
.A1(n_1634),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_1852)
);

O2A1O1Ixp33_ASAP7_75t_SL g1853 ( 
.A1(n_1633),
.A2(n_515),
.B(n_513),
.C(n_512),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1457),
.B(n_1473),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1500),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1506),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1446),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1473),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1496),
.B(n_183),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_SL g1860 ( 
.A(n_1555),
.B(n_1512),
.Y(n_1860)
);

A2O1A1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1602),
.A2(n_185),
.B(n_186),
.C(n_187),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1513),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1583),
.Y(n_1863)
);

BUFx6f_ASAP7_75t_L g1864 ( 
.A(n_1446),
.Y(n_1864)
);

NOR3xp33_ASAP7_75t_L g1865 ( 
.A(n_1592),
.B(n_187),
.C(n_188),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1560),
.B(n_188),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1560),
.B(n_189),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1512),
.Y(n_1868)
);

INVx6_ASAP7_75t_L g1869 ( 
.A(n_1583),
.Y(n_1869)
);

BUFx2_ASAP7_75t_L g1870 ( 
.A(n_1512),
.Y(n_1870)
);

BUFx6f_ASAP7_75t_L g1871 ( 
.A(n_1497),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1528),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1538),
.B(n_189),
.Y(n_1873)
);

NOR2x1_ASAP7_75t_L g1874 ( 
.A(n_1630),
.B(n_190),
.Y(n_1874)
);

O2A1O1Ixp33_ASAP7_75t_L g1875 ( 
.A1(n_1494),
.A2(n_191),
.B(n_192),
.C(n_193),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1510),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1388),
.A2(n_447),
.B(n_446),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1512),
.B(n_1393),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1497),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1518),
.Y(n_1880)
);

O2A1O1Ixp33_ASAP7_75t_L g1881 ( 
.A1(n_1493),
.A2(n_191),
.B(n_194),
.C(n_196),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1526),
.Y(n_1882)
);

BUFx6f_ASAP7_75t_L g1883 ( 
.A(n_1497),
.Y(n_1883)
);

AND2x2_ASAP7_75t_SL g1884 ( 
.A(n_1509),
.B(n_194),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1559),
.B(n_196),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1546),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1544),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_SL g1888 ( 
.A1(n_1488),
.A2(n_198),
.B1(n_199),
.B2(n_201),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1608),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1515),
.B(n_203),
.Y(n_1890)
);

OAI22x1_ASAP7_75t_L g1891 ( 
.A1(n_1583),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1394),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1582),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1635),
.Y(n_1894)
);

A2O1A1Ixp33_ASAP7_75t_L g1895 ( 
.A1(n_1610),
.A2(n_208),
.B(n_209),
.C(n_210),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1503),
.B(n_211),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1416),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1418),
.B(n_211),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1644),
.B(n_212),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1424),
.B(n_212),
.Y(n_1900)
);

BUFx3_ASAP7_75t_L g1901 ( 
.A(n_1600),
.Y(n_1901)
);

CKINVDCx5p33_ASAP7_75t_R g1902 ( 
.A(n_1406),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1442),
.B(n_1563),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1644),
.B(n_213),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1434),
.B(n_218),
.Y(n_1905)
);

INVx4_ASAP7_75t_L g1906 ( 
.A(n_1644),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1606),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1482),
.B(n_220),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1604),
.B(n_1392),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1477),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1546),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1386),
.B(n_221),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1611),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1635),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1404),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_L g1916 ( 
.A(n_1625),
.B(n_222),
.C(n_223),
.Y(n_1916)
);

OAI21xp33_ASAP7_75t_L g1917 ( 
.A1(n_1626),
.A2(n_224),
.B(n_225),
.Y(n_1917)
);

O2A1O1Ixp33_ASAP7_75t_L g1918 ( 
.A1(n_1481),
.A2(n_226),
.B(n_230),
.C(n_231),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1600),
.B(n_231),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1619),
.B(n_232),
.Y(n_1920)
);

OAI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1624),
.A2(n_510),
.B(n_508),
.Y(n_1921)
);

BUFx3_ASAP7_75t_L g1922 ( 
.A(n_1562),
.Y(n_1922)
);

BUFx8_ASAP7_75t_L g1923 ( 
.A(n_1561),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1605),
.B(n_232),
.Y(n_1924)
);

O2A1O1Ixp33_ASAP7_75t_L g1925 ( 
.A1(n_1596),
.A2(n_233),
.B(n_234),
.C(n_235),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1614),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1507),
.B(n_233),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1507),
.B(n_234),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1627),
.B(n_236),
.Y(n_1929)
);

INVx3_ASAP7_75t_L g1930 ( 
.A(n_1632),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1614),
.B(n_237),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1622),
.B(n_238),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1622),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_1933)
);

OR2x6_ASAP7_75t_L g1934 ( 
.A(n_1615),
.B(n_239),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1615),
.B(n_242),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1387),
.B(n_243),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1532),
.B(n_243),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1536),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1532),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1502),
.B(n_244),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1422),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1532),
.B(n_247),
.Y(n_1942)
);

OR2x6_ASAP7_75t_L g1943 ( 
.A(n_1405),
.B(n_248),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1532),
.B(n_248),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1409),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1502),
.B(n_249),
.Y(n_1946)
);

OR2x6_ASAP7_75t_SL g1947 ( 
.A(n_1419),
.B(n_250),
.Y(n_1947)
);

NOR2xp33_ASAP7_75t_SL g1948 ( 
.A(n_1397),
.B(n_250),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1389),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1395),
.A2(n_500),
.B(n_496),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1395),
.A2(n_495),
.B(n_494),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1387),
.B(n_252),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1384),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1409),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1532),
.B(n_253),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1387),
.B(n_254),
.Y(n_1956)
);

NOR2x1_ASAP7_75t_SL g1957 ( 
.A(n_1387),
.B(n_254),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1599),
.A2(n_255),
.B1(n_257),
.B2(n_260),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1532),
.B(n_255),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1443),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1599),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1502),
.B(n_261),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1409),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1502),
.B(n_262),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1384),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1387),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1532),
.B(n_263),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1387),
.B(n_263),
.Y(n_1968)
);

BUFx3_ASAP7_75t_L g1969 ( 
.A(n_1384),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_R g1970 ( 
.A(n_1427),
.B(n_264),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1387),
.B(n_264),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1387),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1532),
.B(n_265),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_SL g1974 ( 
.A(n_1387),
.B(n_266),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1532),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_1975)
);

OR2x6_ASAP7_75t_L g1976 ( 
.A(n_1405),
.B(n_268),
.Y(n_1976)
);

CKINVDCx20_ASAP7_75t_R g1977 ( 
.A(n_1384),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1502),
.B(n_269),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1387),
.B(n_270),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1422),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1536),
.Y(n_1981)
);

AOI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1395),
.A2(n_457),
.B(n_471),
.Y(n_1982)
);

NOR3xp33_ASAP7_75t_L g1983 ( 
.A(n_1498),
.B(n_271),
.C(n_272),
.Y(n_1983)
);

O2A1O1Ixp33_ASAP7_75t_L g1984 ( 
.A1(n_1504),
.A2(n_275),
.B(n_276),
.C(n_277),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1395),
.A2(n_456),
.B(n_466),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1805),
.Y(n_1986)
);

AO21x2_ASAP7_75t_L g1987 ( 
.A1(n_1652),
.A2(n_472),
.B(n_460),
.Y(n_1987)
);

BUFx2_ASAP7_75t_R g1988 ( 
.A(n_1672),
.Y(n_1988)
);

OAI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1654),
.A2(n_275),
.B(n_276),
.Y(n_1989)
);

BUFx12f_ASAP7_75t_L g1990 ( 
.A(n_1653),
.Y(n_1990)
);

AOI22x1_ASAP7_75t_L g1991 ( 
.A1(n_1791),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_1991)
);

AO21x2_ASAP7_75t_L g1992 ( 
.A1(n_1740),
.A2(n_451),
.B(n_449),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1788),
.Y(n_1993)
);

INVxp67_ASAP7_75t_SL g1994 ( 
.A(n_1660),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1718),
.B(n_282),
.Y(n_1995)
);

AOI22x1_ASAP7_75t_L g1996 ( 
.A1(n_1724),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1651),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1658),
.Y(n_1998)
);

BUFx3_ASAP7_75t_L g1999 ( 
.A(n_1745),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1649),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1742),
.Y(n_2001)
);

OAI21x1_ASAP7_75t_L g2002 ( 
.A1(n_1950),
.A2(n_286),
.B(n_287),
.Y(n_2002)
);

NAND2x1p5_ASAP7_75t_L g2003 ( 
.A(n_1805),
.B(n_286),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1662),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1945),
.Y(n_2005)
);

BUFx12f_ASAP7_75t_L g2006 ( 
.A(n_1828),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1649),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1657),
.B(n_288),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1684),
.Y(n_2009)
);

INVx8_ASAP7_75t_L g2010 ( 
.A(n_1805),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1788),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1954),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1977),
.Y(n_2013)
);

CKINVDCx8_ASAP7_75t_R g2014 ( 
.A(n_1816),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1732),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1749),
.B(n_288),
.Y(n_2016)
);

AO21x2_ASAP7_75t_L g2017 ( 
.A1(n_1985),
.A2(n_290),
.B(n_291),
.Y(n_2017)
);

AO21x2_ASAP7_75t_L g2018 ( 
.A1(n_1951),
.A2(n_292),
.B(n_293),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1963),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1790),
.B(n_293),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1650),
.Y(n_2021)
);

BUFx2_ASAP7_75t_R g2022 ( 
.A(n_1969),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1738),
.A2(n_1666),
.B(n_1903),
.Y(n_2023)
);

INVx2_ASAP7_75t_SL g2024 ( 
.A(n_1702),
.Y(n_2024)
);

INVx3_ASAP7_75t_L g2025 ( 
.A(n_1841),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1960),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1688),
.B(n_1849),
.Y(n_2027)
);

INVx4_ASAP7_75t_L g2028 ( 
.A(n_1716),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1802),
.B(n_295),
.Y(n_2029)
);

AOI22x1_ASAP7_75t_L g2030 ( 
.A1(n_1767),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_2030)
);

INVx4_ASAP7_75t_L g2031 ( 
.A(n_1716),
.Y(n_2031)
);

OAI21x1_ASAP7_75t_L g2032 ( 
.A1(n_1982),
.A2(n_298),
.B(n_299),
.Y(n_2032)
);

NAND2x1p5_ASAP7_75t_L g2033 ( 
.A(n_1714),
.B(n_302),
.Y(n_2033)
);

INVx4_ASAP7_75t_L g2034 ( 
.A(n_1716),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1723),
.B(n_305),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1854),
.B(n_306),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1686),
.Y(n_2037)
);

INVx1_ASAP7_75t_SL g2038 ( 
.A(n_1800),
.Y(n_2038)
);

BUFx2_ASAP7_75t_SL g2039 ( 
.A(n_1953),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1860),
.A2(n_308),
.B1(n_311),
.B2(n_312),
.Y(n_2040)
);

BUFx4_ASAP7_75t_SL g2041 ( 
.A(n_1648),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1689),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1966),
.Y(n_2043)
);

BUFx3_ASAP7_75t_L g2044 ( 
.A(n_1972),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1708),
.Y(n_2045)
);

BUFx4f_ASAP7_75t_L g2046 ( 
.A(n_1943),
.Y(n_2046)
);

INVx3_ASAP7_75t_L g2047 ( 
.A(n_1972),
.Y(n_2047)
);

INVx3_ASAP7_75t_SL g2048 ( 
.A(n_1965),
.Y(n_2048)
);

CKINVDCx14_ASAP7_75t_R g2049 ( 
.A(n_1680),
.Y(n_2049)
);

NAND2x1p5_ASAP7_75t_L g2050 ( 
.A(n_1714),
.B(n_1723),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1677),
.Y(n_2051)
);

BUFx12f_ASAP7_75t_L g2052 ( 
.A(n_1828),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1938),
.Y(n_2053)
);

BUFx3_ASAP7_75t_L g2054 ( 
.A(n_1869),
.Y(n_2054)
);

INVx3_ASAP7_75t_L g2055 ( 
.A(n_1792),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1869),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1712),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1892),
.B(n_1897),
.Y(n_2058)
);

AO21x2_ASAP7_75t_L g2059 ( 
.A1(n_1656),
.A2(n_1926),
.B(n_1661),
.Y(n_2059)
);

INVx4_ASAP7_75t_L g2060 ( 
.A(n_1702),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1728),
.Y(n_2061)
);

AO21x2_ASAP7_75t_L g2062 ( 
.A1(n_1656),
.A2(n_1851),
.B(n_1921),
.Y(n_2062)
);

INVx1_ASAP7_75t_SL g2063 ( 
.A(n_1775),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1938),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_1863),
.Y(n_2065)
);

INVx4_ASAP7_75t_L g2066 ( 
.A(n_1936),
.Y(n_2066)
);

INVxp67_ASAP7_75t_L g2067 ( 
.A(n_1949),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1691),
.Y(n_2068)
);

NAND2x1_ASAP7_75t_L g2069 ( 
.A(n_1906),
.B(n_1938),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1770),
.Y(n_2070)
);

INVxp67_ASAP7_75t_SL g2071 ( 
.A(n_1981),
.Y(n_2071)
);

AO21x2_ASAP7_75t_L g2072 ( 
.A1(n_1713),
.A2(n_1715),
.B(n_1836),
.Y(n_2072)
);

OR2x6_ASAP7_75t_L g2073 ( 
.A(n_1943),
.B(n_1648),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1735),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1836),
.B(n_1679),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1819),
.Y(n_2076)
);

OA21x2_ASAP7_75t_L g2077 ( 
.A1(n_1917),
.A2(n_1705),
.B(n_1755),
.Y(n_2077)
);

INVx6_ASAP7_75t_SL g2078 ( 
.A(n_1936),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1825),
.Y(n_2079)
);

BUFx3_ASAP7_75t_L g2080 ( 
.A(n_1771),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1692),
.B(n_1737),
.Y(n_2081)
);

INVx1_ASAP7_75t_SL g2082 ( 
.A(n_1775),
.Y(n_2082)
);

BUFx12f_ASAP7_75t_L g2083 ( 
.A(n_1923),
.Y(n_2083)
);

AOI22x1_ASAP7_75t_L g2084 ( 
.A1(n_1785),
.A2(n_1743),
.B1(n_1739),
.B2(n_1729),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_1833),
.B(n_1914),
.Y(n_2085)
);

AO21x2_ASAP7_75t_L g2086 ( 
.A1(n_1932),
.A2(n_1655),
.B(n_1917),
.Y(n_2086)
);

AO21x2_ASAP7_75t_L g2087 ( 
.A1(n_1931),
.A2(n_1927),
.B(n_1899),
.Y(n_2087)
);

INVx3_ASAP7_75t_L g2088 ( 
.A(n_1771),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_1736),
.Y(n_2089)
);

AO21x2_ASAP7_75t_L g2090 ( 
.A1(n_1896),
.A2(n_1904),
.B(n_1645),
.Y(n_2090)
);

BUFx12f_ASAP7_75t_L g2091 ( 
.A(n_1923),
.Y(n_2091)
);

OAI21xp5_ASAP7_75t_L g2092 ( 
.A1(n_1699),
.A2(n_1725),
.B(n_1720),
.Y(n_2092)
);

NAND2x1_ASAP7_75t_L g2093 ( 
.A(n_1906),
.B(n_1757),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1976),
.B(n_1850),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1852),
.A2(n_1780),
.B1(n_1685),
.B2(n_1812),
.Y(n_2095)
);

INVx3_ASAP7_75t_L g2096 ( 
.A(n_1956),
.Y(n_2096)
);

CKINVDCx6p67_ASAP7_75t_R g2097 ( 
.A(n_1741),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1709),
.Y(n_2098)
);

INVxp67_ASAP7_75t_L g2099 ( 
.A(n_1704),
.Y(n_2099)
);

OA21x2_ASAP7_75t_L g2100 ( 
.A1(n_1707),
.A2(n_1877),
.B(n_1768),
.Y(n_2100)
);

INVx3_ASAP7_75t_L g2101 ( 
.A(n_1956),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1842),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1835),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_SL g2104 ( 
.A1(n_1888),
.A2(n_1852),
.B1(n_1884),
.B2(n_1970),
.Y(n_2104)
);

AO21x2_ASAP7_75t_L g2105 ( 
.A1(n_1937),
.A2(n_1944),
.B(n_1942),
.Y(n_2105)
);

BUFx3_ASAP7_75t_L g2106 ( 
.A(n_1746),
.Y(n_2106)
);

AOI21x1_ASAP7_75t_L g2107 ( 
.A1(n_1878),
.A2(n_1659),
.B(n_1646),
.Y(n_2107)
);

BUFx12f_ASAP7_75t_L g2108 ( 
.A(n_1673),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1855),
.Y(n_2109)
);

NAND2x1p5_ASAP7_75t_L g2110 ( 
.A(n_1776),
.B(n_1817),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_L g2111 ( 
.A(n_1894),
.B(n_1913),
.Y(n_2111)
);

BUFx2_ASAP7_75t_SL g2112 ( 
.A(n_1711),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1710),
.B(n_1823),
.Y(n_2113)
);

AOI22x1_ASAP7_75t_L g2114 ( 
.A1(n_1818),
.A2(n_1891),
.B1(n_1870),
.B2(n_1829),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1856),
.Y(n_2115)
);

OAI21x1_ASAP7_75t_L g2116 ( 
.A1(n_1874),
.A2(n_1664),
.B(n_1925),
.Y(n_2116)
);

INVx3_ASAP7_75t_L g2117 ( 
.A(n_1798),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1862),
.Y(n_2118)
);

INVx6_ASAP7_75t_L g2119 ( 
.A(n_1711),
.Y(n_2119)
);

OAI21x1_ASAP7_75t_L g2120 ( 
.A1(n_1874),
.A2(n_1959),
.B(n_1955),
.Y(n_2120)
);

OAI21x1_ASAP7_75t_L g2121 ( 
.A1(n_1967),
.A2(n_1973),
.B(n_1929),
.Y(n_2121)
);

AO21x2_ASAP7_75t_L g2122 ( 
.A1(n_1681),
.A2(n_1853),
.B(n_1920),
.Y(n_2122)
);

AO21x2_ASAP7_75t_L g2123 ( 
.A1(n_1924),
.A2(n_1839),
.B(n_1831),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_1876),
.B(n_1880),
.Y(n_2124)
);

OAI21xp5_ASAP7_75t_L g2125 ( 
.A1(n_1782),
.A2(n_1795),
.B(n_1898),
.Y(n_2125)
);

INVx4_ASAP7_75t_L g2126 ( 
.A(n_1753),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1882),
.Y(n_2127)
);

OAI21x1_ASAP7_75t_L g2128 ( 
.A1(n_1952),
.A2(n_1971),
.B(n_1968),
.Y(n_2128)
);

INVx8_ASAP7_75t_L g2129 ( 
.A(n_1753),
.Y(n_2129)
);

AO21x2_ASAP7_75t_L g2130 ( 
.A1(n_1668),
.A2(n_1670),
.B(n_1747),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_1701),
.A2(n_1706),
.B(n_1797),
.Y(n_2131)
);

INVx6_ASAP7_75t_L g2132 ( 
.A(n_1736),
.Y(n_2132)
);

AND2x4_ASAP7_75t_L g2133 ( 
.A(n_1911),
.B(n_1671),
.Y(n_2133)
);

AO21x2_ASAP7_75t_L g2134 ( 
.A1(n_1762),
.A2(n_1845),
.B(n_1815),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1830),
.B(n_1760),
.Y(n_2135)
);

BUFx10_ASAP7_75t_L g2136 ( 
.A(n_1751),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1826),
.Y(n_2137)
);

INVx3_ASAP7_75t_L g2138 ( 
.A(n_1798),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1872),
.Y(n_2139)
);

HB1xp67_ASAP7_75t_L g2140 ( 
.A(n_1751),
.Y(n_2140)
);

AO21x2_ASAP7_75t_L g2141 ( 
.A1(n_1848),
.A2(n_1861),
.B(n_1717),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1826),
.Y(n_2142)
);

INVx3_ASAP7_75t_L g2143 ( 
.A(n_1759),
.Y(n_2143)
);

INVx8_ASAP7_75t_L g2144 ( 
.A(n_1744),
.Y(n_2144)
);

CKINVDCx16_ASAP7_75t_R g2145 ( 
.A(n_1690),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1846),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_1843),
.B(n_1676),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_1922),
.B(n_1783),
.Y(n_2148)
);

AO21x2_ASAP7_75t_L g2149 ( 
.A1(n_1928),
.A2(n_1979),
.B(n_1974),
.Y(n_2149)
);

CKINVDCx20_ASAP7_75t_R g2150 ( 
.A(n_1678),
.Y(n_2150)
);

BUFx2_ASAP7_75t_L g2151 ( 
.A(n_1726),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1759),
.Y(n_2152)
);

BUFx12f_ASAP7_75t_L g2153 ( 
.A(n_1779),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_1759),
.Y(n_2154)
);

OR3x4_ASAP7_75t_SL g2155 ( 
.A(n_1947),
.B(n_1888),
.C(n_1727),
.Y(n_2155)
);

BUFx2_ASAP7_75t_L g2156 ( 
.A(n_1696),
.Y(n_2156)
);

OA21x2_ASAP7_75t_L g2157 ( 
.A1(n_1895),
.A2(n_1808),
.B(n_1958),
.Y(n_2157)
);

AOI22x1_ASAP7_75t_L g2158 ( 
.A1(n_1663),
.A2(n_1935),
.B1(n_1844),
.B2(n_1820),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1763),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_L g2160 ( 
.A(n_1763),
.Y(n_2160)
);

BUFx2_ASAP7_75t_L g2161 ( 
.A(n_1744),
.Y(n_2161)
);

INVx6_ASAP7_75t_L g2162 ( 
.A(n_1674),
.Y(n_2162)
);

INVx1_ASAP7_75t_SL g2163 ( 
.A(n_1786),
.Y(n_2163)
);

AOI21xp5_ASAP7_75t_L g2164 ( 
.A1(n_1900),
.A2(n_1750),
.B(n_1675),
.Y(n_2164)
);

OAI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_1890),
.A2(n_1667),
.B(n_1799),
.Y(n_2165)
);

OAI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_1801),
.A2(n_1867),
.B(n_1866),
.Y(n_2166)
);

AO21x2_ASAP7_75t_L g2167 ( 
.A1(n_1859),
.A2(n_1919),
.B(n_1961),
.Y(n_2167)
);

BUFx2_ASAP7_75t_L g2168 ( 
.A(n_1674),
.Y(n_2168)
);

BUFx12f_ASAP7_75t_L g2169 ( 
.A(n_1834),
.Y(n_2169)
);

BUFx2_ASAP7_75t_R g2170 ( 
.A(n_1902),
.Y(n_2170)
);

INVx1_ASAP7_75t_SL g2171 ( 
.A(n_1683),
.Y(n_2171)
);

AO21x2_ASAP7_75t_L g2172 ( 
.A1(n_1958),
.A2(n_1961),
.B(n_1756),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_1766),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_1671),
.B(n_1700),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1669),
.B(n_1752),
.Y(n_2175)
);

INVx5_ASAP7_75t_L g2176 ( 
.A(n_1766),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_1730),
.B(n_1811),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1766),
.Y(n_2178)
);

INVx1_ASAP7_75t_SL g2179 ( 
.A(n_1772),
.Y(n_2179)
);

INVx5_ASAP7_75t_L g2180 ( 
.A(n_1820),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_1807),
.B(n_1838),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1822),
.Y(n_2182)
);

AO21x2_ASAP7_75t_L g2183 ( 
.A1(n_1813),
.A2(n_1809),
.B(n_1810),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1844),
.Y(n_2184)
);

OA21x2_ASAP7_75t_L g2185 ( 
.A1(n_1679),
.A2(n_1907),
.B(n_1941),
.Y(n_2185)
);

OAI21x1_ASAP7_75t_L g2186 ( 
.A1(n_1918),
.A2(n_1930),
.B(n_1821),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1840),
.B(n_1847),
.Y(n_2187)
);

AO21x2_ASAP7_75t_L g2188 ( 
.A1(n_1697),
.A2(n_1837),
.B(n_1875),
.Y(n_2188)
);

INVx8_ASAP7_75t_L g2189 ( 
.A(n_1934),
.Y(n_2189)
);

AO21x2_ASAP7_75t_L g2190 ( 
.A1(n_1881),
.A2(n_1907),
.B(n_1764),
.Y(n_2190)
);

CKINVDCx20_ASAP7_75t_R g2191 ( 
.A(n_1687),
.Y(n_2191)
);

OAI21x1_ASAP7_75t_L g2192 ( 
.A1(n_1787),
.A2(n_1984),
.B(n_1682),
.Y(n_2192)
);

AND2x2_ASAP7_75t_L g2193 ( 
.A(n_1940),
.B(n_1946),
.Y(n_2193)
);

OAI21xp5_ASAP7_75t_L g2194 ( 
.A1(n_1781),
.A2(n_1796),
.B(n_1793),
.Y(n_2194)
);

OR2x2_ASAP7_75t_L g2195 ( 
.A(n_1803),
.B(n_1962),
.Y(n_2195)
);

HB1xp67_ASAP7_75t_L g2196 ( 
.A(n_1934),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1857),
.Y(n_2197)
);

AO21x2_ASAP7_75t_L g2198 ( 
.A1(n_1933),
.A2(n_1693),
.B(n_1734),
.Y(n_2198)
);

INVx4_ASAP7_75t_L g2199 ( 
.A(n_1857),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1864),
.Y(n_2200)
);

OAI21x1_ASAP7_75t_SL g2201 ( 
.A1(n_1957),
.A2(n_1789),
.B(n_1773),
.Y(n_2201)
);

INVx6_ASAP7_75t_L g2202 ( 
.A(n_1910),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_1804),
.B(n_1909),
.Y(n_2203)
);

BUFx8_ASAP7_75t_SL g2204 ( 
.A(n_1722),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_L g2205 ( 
.A(n_1873),
.B(n_1978),
.Y(n_2205)
);

BUFx4_ASAP7_75t_SL g2206 ( 
.A(n_1901),
.Y(n_2206)
);

OAI21x1_ASAP7_75t_L g2207 ( 
.A1(n_1761),
.A2(n_1886),
.B(n_1694),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1722),
.Y(n_2208)
);

OAI21x1_ASAP7_75t_L g2209 ( 
.A1(n_1748),
.A2(n_1814),
.B(n_1832),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1772),
.Y(n_2210)
);

OAI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_1868),
.A2(n_1893),
.B(n_1905),
.Y(n_2211)
);

BUFx4f_ASAP7_75t_L g2212 ( 
.A(n_1864),
.Y(n_2212)
);

CKINVDCx6p67_ASAP7_75t_R g2213 ( 
.A(n_1827),
.Y(n_2213)
);

INVx2_ASAP7_75t_SL g2214 ( 
.A(n_1733),
.Y(n_2214)
);

AO21x2_ASAP7_75t_L g2215 ( 
.A1(n_1719),
.A2(n_1983),
.B(n_1647),
.Y(n_2215)
);

INVx1_ASAP7_75t_SL g2216 ( 
.A(n_1964),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1789),
.Y(n_2217)
);

CKINVDCx11_ASAP7_75t_R g2218 ( 
.A(n_1758),
.Y(n_2218)
);

OAI22xp33_ASAP7_75t_SL g2219 ( 
.A1(n_1948),
.A2(n_1777),
.B1(n_1773),
.B2(n_1698),
.Y(n_2219)
);

BUFx3_ASAP7_75t_L g2220 ( 
.A(n_1864),
.Y(n_2220)
);

AO21x2_ASAP7_75t_L g2221 ( 
.A1(n_1777),
.A2(n_1695),
.B(n_1731),
.Y(n_2221)
);

NAND2x1p5_ASAP7_75t_L g2222 ( 
.A(n_1871),
.B(n_1883),
.Y(n_2222)
);

INVx2_ASAP7_75t_SL g2223 ( 
.A(n_1915),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1939),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_1879),
.B(n_1883),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1975),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1865),
.B(n_1885),
.Y(n_2227)
);

OAI21x1_ASAP7_75t_SL g2228 ( 
.A1(n_1769),
.A2(n_1774),
.B(n_1887),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1765),
.Y(n_2229)
);

OAI21x1_ASAP7_75t_SL g2230 ( 
.A1(n_1889),
.A2(n_1806),
.B(n_1858),
.Y(n_2230)
);

AO21x2_ASAP7_75t_L g2231 ( 
.A1(n_1916),
.A2(n_1912),
.B(n_1908),
.Y(n_2231)
);

INVx8_ASAP7_75t_L g2232 ( 
.A(n_1778),
.Y(n_2232)
);

OAI21x1_ASAP7_75t_L g2233 ( 
.A1(n_1980),
.A2(n_1721),
.B(n_1703),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_1754),
.A2(n_1784),
.B(n_1794),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_1824),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1824),
.B(n_1754),
.Y(n_2236)
);

BUFx6f_ASAP7_75t_L g2237 ( 
.A(n_1824),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_1784),
.Y(n_2238)
);

OA21x2_ASAP7_75t_L g2239 ( 
.A1(n_1652),
.A2(n_1395),
.B(n_1162),
.Y(n_2239)
);

INVx2_ASAP7_75t_SL g2240 ( 
.A(n_1653),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_1718),
.B(n_1790),
.Y(n_2241)
);

AO21x2_ASAP7_75t_L g2242 ( 
.A1(n_1652),
.A2(n_1665),
.B(n_1186),
.Y(n_2242)
);

BUFx3_ASAP7_75t_L g2243 ( 
.A(n_1745),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_1666),
.B(n_1532),
.Y(n_2244)
);

NAND2x1p5_ASAP7_75t_L g2245 ( 
.A(n_1805),
.B(n_1387),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1651),
.Y(n_2246)
);

INVx5_ASAP7_75t_SL g2247 ( 
.A(n_1648),
.Y(n_2247)
);

OAI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_1654),
.A2(n_1249),
.B(n_1339),
.Y(n_2248)
);

OAI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_1654),
.A2(n_1249),
.B(n_1339),
.Y(n_2249)
);

AO21x2_ASAP7_75t_L g2250 ( 
.A1(n_1652),
.A2(n_1665),
.B(n_1186),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1651),
.Y(n_2251)
);

INVx2_ASAP7_75t_SL g2252 ( 
.A(n_1653),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_1666),
.B(n_1532),
.Y(n_2253)
);

INVx1_ASAP7_75t_SL g2254 ( 
.A(n_1684),
.Y(n_2254)
);

AOI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_2218),
.A2(n_2147),
.B1(n_2189),
.B2(n_2073),
.Y(n_2255)
);

INVx2_ASAP7_75t_SL g2256 ( 
.A(n_1990),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2068),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_2212),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1997),
.Y(n_2259)
);

BUFx3_ASAP7_75t_L g2260 ( 
.A(n_1990),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1998),
.Y(n_2261)
);

OAI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_2046),
.A2(n_2073),
.B1(n_2189),
.B2(n_2196),
.Y(n_2262)
);

BUFx3_ASAP7_75t_L g2263 ( 
.A(n_2001),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_2073),
.B(n_2066),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2004),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_SL g2266 ( 
.A1(n_2201),
.A2(n_2066),
.B(n_2158),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_2083),
.Y(n_2267)
);

NAND2x1p5_ASAP7_75t_L g2268 ( 
.A(n_2060),
.B(n_2046),
.Y(n_2268)
);

OAI22xp33_ASAP7_75t_SL g2269 ( 
.A1(n_2196),
.A2(n_2075),
.B1(n_2147),
.B2(n_2033),
.Y(n_2269)
);

BUFx3_ASAP7_75t_L g2270 ( 
.A(n_2001),
.Y(n_2270)
);

OAI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2189),
.A2(n_2095),
.B1(n_1994),
.B2(n_2247),
.Y(n_2271)
);

NAND2x1p5_ASAP7_75t_L g2272 ( 
.A(n_2060),
.B(n_2080),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2005),
.Y(n_2273)
);

INVx3_ASAP7_75t_L g2274 ( 
.A(n_2245),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_2212),
.Y(n_2275)
);

INVx1_ASAP7_75t_SL g2276 ( 
.A(n_2078),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2217),
.B(n_2241),
.Y(n_2277)
);

CKINVDCx11_ASAP7_75t_R g2278 ( 
.A(n_2083),
.Y(n_2278)
);

AOI22xp33_ASAP7_75t_L g2279 ( 
.A1(n_2218),
.A2(n_2095),
.B1(n_2104),
.B2(n_2094),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2012),
.Y(n_2280)
);

NAND2x1p5_ASAP7_75t_L g2281 ( 
.A(n_2176),
.B(n_2180),
.Y(n_2281)
);

OAI22xp33_ASAP7_75t_L g2282 ( 
.A1(n_2129),
.A2(n_2144),
.B1(n_2126),
.B2(n_2156),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2058),
.B(n_1995),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2058),
.B(n_2124),
.Y(n_2284)
);

BUFx2_ASAP7_75t_L g2285 ( 
.A(n_2078),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2019),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2124),
.B(n_2021),
.Y(n_2287)
);

AOI22xp33_ASAP7_75t_SL g2288 ( 
.A1(n_2247),
.A2(n_2129),
.B1(n_2144),
.B2(n_2049),
.Y(n_2288)
);

AOI22xp33_ASAP7_75t_L g2289 ( 
.A1(n_2104),
.A2(n_2215),
.B1(n_2185),
.B2(n_2247),
.Y(n_2289)
);

BUFx2_ASAP7_75t_L g2290 ( 
.A(n_2078),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2015),
.Y(n_2291)
);

OAI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_1994),
.A2(n_2140),
.B1(n_2253),
.B2(n_2244),
.Y(n_2292)
);

INVx2_ASAP7_75t_SL g2293 ( 
.A(n_2006),
.Y(n_2293)
);

BUFx3_ASAP7_75t_L g2294 ( 
.A(n_2006),
.Y(n_2294)
);

INVx6_ASAP7_75t_L g2295 ( 
.A(n_2052),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2037),
.Y(n_2296)
);

AOI22xp33_ASAP7_75t_SL g2297 ( 
.A1(n_2129),
.A2(n_2144),
.B1(n_2049),
.B2(n_2219),
.Y(n_2297)
);

CKINVDCx20_ASAP7_75t_R g2298 ( 
.A(n_2013),
.Y(n_2298)
);

BUFx6f_ASAP7_75t_L g2299 ( 
.A(n_2010),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2098),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2081),
.B(n_2244),
.Y(n_2301)
);

INVxp33_ASAP7_75t_L g2302 ( 
.A(n_2204),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2042),
.Y(n_2303)
);

INVx4_ASAP7_75t_L g2304 ( 
.A(n_2010),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2038),
.B(n_2204),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2045),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2244),
.B(n_2253),
.Y(n_2307)
);

INVx6_ASAP7_75t_L g2308 ( 
.A(n_2052),
.Y(n_2308)
);

INVx2_ASAP7_75t_SL g2309 ( 
.A(n_2206),
.Y(n_2309)
);

BUFx2_ASAP7_75t_SL g2310 ( 
.A(n_2014),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2057),
.Y(n_2311)
);

CKINVDCx8_ASAP7_75t_R g2312 ( 
.A(n_2013),
.Y(n_2312)
);

BUFx2_ASAP7_75t_L g2313 ( 
.A(n_2065),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2061),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_2009),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2246),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2251),
.Y(n_2317)
);

BUFx3_ASAP7_75t_L g2318 ( 
.A(n_2048),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_2215),
.A2(n_2185),
.B1(n_2205),
.B2(n_2177),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2074),
.Y(n_2320)
);

OAI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_2145),
.A2(n_2161),
.B1(n_2140),
.B2(n_2179),
.Y(n_2321)
);

INVx6_ASAP7_75t_L g2322 ( 
.A(n_2091),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2103),
.Y(n_2323)
);

INVx4_ASAP7_75t_L g2324 ( 
.A(n_2010),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2076),
.Y(n_2325)
);

BUFx2_ASAP7_75t_SL g2326 ( 
.A(n_2024),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2079),
.Y(n_2327)
);

OAI21x1_ASAP7_75t_SL g2328 ( 
.A1(n_2228),
.A2(n_2114),
.B(n_1989),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2102),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2253),
.B(n_2023),
.Y(n_2330)
);

OAI22x1_ASAP7_75t_L g2331 ( 
.A1(n_2041),
.A2(n_2155),
.B1(n_2033),
.B2(n_2171),
.Y(n_2331)
);

OAI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_2185),
.A2(n_2016),
.B1(n_2101),
.B2(n_2096),
.Y(n_2332)
);

OR2x6_ASAP7_75t_L g2333 ( 
.A(n_2050),
.B(n_2112),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2109),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2224),
.B(n_2226),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2115),
.Y(n_2336)
);

OR2x6_ASAP7_75t_L g2337 ( 
.A(n_2050),
.B(n_2003),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2127),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2026),
.B(n_2067),
.Y(n_2339)
);

INVx2_ASAP7_75t_SL g2340 ( 
.A(n_2206),
.Y(n_2340)
);

BUFx3_ASAP7_75t_L g2341 ( 
.A(n_2048),
.Y(n_2341)
);

CKINVDCx11_ASAP7_75t_R g2342 ( 
.A(n_2091),
.Y(n_2342)
);

AOI22xp33_ASAP7_75t_SL g2343 ( 
.A1(n_2172),
.A2(n_1991),
.B1(n_2191),
.B2(n_2041),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2146),
.Y(n_2344)
);

AOI22xp33_ASAP7_75t_L g2345 ( 
.A1(n_2205),
.A2(n_2177),
.B1(n_2227),
.B2(n_2193),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2118),
.Y(n_2346)
);

BUFx6f_ASAP7_75t_L g2347 ( 
.A(n_2176),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2139),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2139),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2254),
.Y(n_2350)
);

HB1xp67_ASAP7_75t_L g2351 ( 
.A(n_2071),
.Y(n_2351)
);

BUFx2_ASAP7_75t_L g2352 ( 
.A(n_2065),
.Y(n_2352)
);

BUFx10_ASAP7_75t_L g2353 ( 
.A(n_2252),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_1996),
.Y(n_2354)
);

AOI22xp33_ASAP7_75t_L g2355 ( 
.A1(n_2230),
.A2(n_2229),
.B1(n_2172),
.B2(n_2165),
.Y(n_2355)
);

OAI22xp33_ASAP7_75t_L g2356 ( 
.A1(n_2213),
.A2(n_2191),
.B1(n_2099),
.B2(n_2113),
.Y(n_2356)
);

BUFx2_ASAP7_75t_L g2357 ( 
.A(n_2070),
.Y(n_2357)
);

AOI22xp33_ASAP7_75t_L g2358 ( 
.A1(n_2175),
.A2(n_2232),
.B1(n_2198),
.B2(n_2195),
.Y(n_2358)
);

OAI22xp5_ASAP7_75t_L g2359 ( 
.A1(n_2096),
.A2(n_2101),
.B1(n_2003),
.B2(n_2029),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2111),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2111),
.Y(n_2361)
);

CKINVDCx12_ASAP7_75t_R g2362 ( 
.A(n_1988),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2099),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2130),
.B(n_2105),
.Y(n_2364)
);

NOR2x1_ASAP7_75t_R g2365 ( 
.A(n_2153),
.B(n_2039),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2137),
.Y(n_2366)
);

INVxp33_ASAP7_75t_L g2367 ( 
.A(n_2085),
.Y(n_2367)
);

AOI21x1_ASAP7_75t_L g2368 ( 
.A1(n_2077),
.A2(n_2239),
.B(n_2120),
.Y(n_2368)
);

INVx8_ASAP7_75t_L g2369 ( 
.A(n_2153),
.Y(n_2369)
);

AOI22xp33_ASAP7_75t_L g2370 ( 
.A1(n_2232),
.A2(n_2198),
.B1(n_2181),
.B2(n_2187),
.Y(n_2370)
);

NAND2x1p5_ASAP7_75t_L g2371 ( 
.A(n_2176),
.B(n_2180),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2142),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2027),
.Y(n_2373)
);

BUFx3_ASAP7_75t_L g2374 ( 
.A(n_1999),
.Y(n_2374)
);

BUFx2_ASAP7_75t_L g2375 ( 
.A(n_1999),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2168),
.B(n_2020),
.Y(n_2376)
);

AOI22xp33_ASAP7_75t_L g2377 ( 
.A1(n_2232),
.A2(n_2181),
.B1(n_2187),
.B2(n_2216),
.Y(n_2377)
);

CKINVDCx11_ASAP7_75t_R g2378 ( 
.A(n_2108),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2223),
.Y(n_2379)
);

BUFx12f_ASAP7_75t_L g2380 ( 
.A(n_2240),
.Y(n_2380)
);

BUFx2_ASAP7_75t_L g2381 ( 
.A(n_2243),
.Y(n_2381)
);

AOI22xp33_ASAP7_75t_L g2382 ( 
.A1(n_2008),
.A2(n_2231),
.B1(n_2203),
.B2(n_2221),
.Y(n_2382)
);

OAI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_2235),
.A2(n_2157),
.B1(n_2135),
.B2(n_2208),
.Y(n_2383)
);

BUFx3_ASAP7_75t_L g2384 ( 
.A(n_2243),
.Y(n_2384)
);

AOI22xp33_ASAP7_75t_SL g2385 ( 
.A1(n_2136),
.A2(n_2132),
.B1(n_2157),
.B2(n_2155),
.Y(n_2385)
);

INVx1_ASAP7_75t_SL g2386 ( 
.A(n_2063),
.Y(n_2386)
);

HB1xp67_ASAP7_75t_L g2387 ( 
.A(n_2071),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_2082),
.B(n_2163),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2210),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2235),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2036),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2036),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2136),
.B(n_2162),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2130),
.B(n_2105),
.Y(n_2394)
);

INVx8_ASAP7_75t_L g2395 ( 
.A(n_2176),
.Y(n_2395)
);

BUFx2_ASAP7_75t_L g2396 ( 
.A(n_2088),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2237),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2162),
.B(n_2054),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2237),
.Y(n_2399)
);

INVx3_ASAP7_75t_L g2400 ( 
.A(n_2028),
.Y(n_2400)
);

AOI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2203),
.A2(n_2157),
.B1(n_2221),
.B2(n_2190),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_2108),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2237),
.Y(n_2403)
);

INVx3_ASAP7_75t_L g2404 ( 
.A(n_2028),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2190),
.B(n_2194),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2035),
.Y(n_2406)
);

INVxp67_ASAP7_75t_L g2407 ( 
.A(n_2035),
.Y(n_2407)
);

INVx1_ASAP7_75t_SL g2408 ( 
.A(n_2151),
.Y(n_2408)
);

AOI22xp33_ASAP7_75t_L g2409 ( 
.A1(n_2231),
.A2(n_2211),
.B1(n_2214),
.B2(n_2167),
.Y(n_2409)
);

INVx3_ASAP7_75t_L g2410 ( 
.A(n_2031),
.Y(n_2410)
);

AOI21x1_ASAP7_75t_L g2411 ( 
.A1(n_2077),
.A2(n_2239),
.B(n_2236),
.Y(n_2411)
);

CKINVDCx14_ASAP7_75t_R g2412 ( 
.A(n_2097),
.Y(n_2412)
);

BUFx4f_ASAP7_75t_L g2413 ( 
.A(n_1993),
.Y(n_2413)
);

BUFx2_ASAP7_75t_R g2414 ( 
.A(n_2025),
.Y(n_2414)
);

AOI21x1_ASAP7_75t_L g2415 ( 
.A1(n_2236),
.A2(n_2131),
.B(n_2107),
.Y(n_2415)
);

INVx2_ASAP7_75t_SL g2416 ( 
.A(n_2119),
.Y(n_2416)
);

INVxp67_ASAP7_75t_L g2417 ( 
.A(n_1986),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2047),
.Y(n_2418)
);

NAND2x1p5_ASAP7_75t_L g2419 ( 
.A(n_2031),
.B(n_2034),
.Y(n_2419)
);

CKINVDCx6p67_ASAP7_75t_R g2420 ( 
.A(n_2169),
.Y(n_2420)
);

NOR2xp33_ASAP7_75t_L g2421 ( 
.A(n_2148),
.B(n_2085),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2119),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2119),
.Y(n_2423)
);

INVx6_ASAP7_75t_L g2424 ( 
.A(n_2132),
.Y(n_2424)
);

AOI22xp33_ASAP7_75t_L g2425 ( 
.A1(n_2167),
.A2(n_2188),
.B1(n_2166),
.B2(n_2092),
.Y(n_2425)
);

AOI22xp33_ASAP7_75t_SL g2426 ( 
.A1(n_2030),
.A2(n_2188),
.B1(n_2134),
.B2(n_2141),
.Y(n_2426)
);

OAI22xp33_ASAP7_75t_L g2427 ( 
.A1(n_2040),
.A2(n_2025),
.B1(n_2162),
.B2(n_2089),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_2043),
.B(n_2044),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2043),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2044),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_1986),
.Y(n_2431)
);

AOI22xp33_ASAP7_75t_L g2432 ( 
.A1(n_2134),
.A2(n_2125),
.B1(n_2141),
.B2(n_2233),
.Y(n_2432)
);

BUFx10_ASAP7_75t_L g2433 ( 
.A(n_2011),
.Y(n_2433)
);

BUFx4_ASAP7_75t_SL g2434 ( 
.A(n_2150),
.Y(n_2434)
);

BUFx3_ASAP7_75t_L g2435 ( 
.A(n_2054),
.Y(n_2435)
);

INVx11_ASAP7_75t_L g2436 ( 
.A(n_2169),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_2150),
.B(n_2056),
.Y(n_2437)
);

AOI21x1_ASAP7_75t_L g2438 ( 
.A1(n_2164),
.A2(n_2234),
.B(n_2100),
.Y(n_2438)
);

INVx1_ASAP7_75t_SL g2439 ( 
.A(n_2106),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2284),
.B(n_2117),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2390),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2257),
.Y(n_2442)
);

BUFx6f_ASAP7_75t_L g2443 ( 
.A(n_2395),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2259),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_2278),
.Y(n_2445)
);

AOI22xp33_ASAP7_75t_L g2446 ( 
.A1(n_2271),
.A2(n_2233),
.B1(n_2123),
.B2(n_2183),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_2342),
.Y(n_2447)
);

OR2x6_ASAP7_75t_L g2448 ( 
.A(n_2369),
.B(n_2022),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2261),
.Y(n_2449)
);

BUFx3_ASAP7_75t_L g2450 ( 
.A(n_2318),
.Y(n_2450)
);

CKINVDCx14_ASAP7_75t_R g2451 ( 
.A(n_2412),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2283),
.B(n_2138),
.Y(n_2452)
);

BUFx3_ASAP7_75t_L g2453 ( 
.A(n_2341),
.Y(n_2453)
);

OR2x6_ASAP7_75t_L g2454 ( 
.A(n_2369),
.B(n_2110),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2373),
.B(n_2133),
.Y(n_2455)
);

AO31x2_ASAP7_75t_L g2456 ( 
.A1(n_2364),
.A2(n_2184),
.A3(n_2064),
.B(n_2159),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2265),
.Y(n_2457)
);

NOR2xp33_ASAP7_75t_R g2458 ( 
.A(n_2369),
.B(n_2138),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2339),
.B(n_2174),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2360),
.B(n_2174),
.Y(n_2460)
);

HB1xp67_ASAP7_75t_L g2461 ( 
.A(n_2315),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_2267),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_R g2463 ( 
.A(n_2298),
.B(n_2143),
.Y(n_2463)
);

NOR2x1p5_ASAP7_75t_L g2464 ( 
.A(n_2304),
.B(n_2238),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2287),
.B(n_2174),
.Y(n_2465)
);

OR2x6_ASAP7_75t_L g2466 ( 
.A(n_2333),
.B(n_2055),
.Y(n_2466)
);

HB1xp67_ASAP7_75t_L g2467 ( 
.A(n_2350),
.Y(n_2467)
);

CKINVDCx5p33_ASAP7_75t_R g2468 ( 
.A(n_2434),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2273),
.Y(n_2469)
);

AND2x2_ASAP7_75t_SL g2470 ( 
.A(n_2255),
.B(n_2199),
.Y(n_2470)
);

CKINVDCx5p33_ASAP7_75t_R g2471 ( 
.A(n_2434),
.Y(n_2471)
);

NAND2xp33_ASAP7_75t_R g2472 ( 
.A(n_2333),
.B(n_2238),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2280),
.Y(n_2473)
);

OAI22xp33_ASAP7_75t_L g2474 ( 
.A1(n_2271),
.A2(n_2055),
.B1(n_2248),
.B2(n_2249),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_2378),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_SL g2476 ( 
.A(n_2269),
.B(n_2000),
.Y(n_2476)
);

INVx2_ASAP7_75t_SL g2477 ( 
.A(n_2295),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2361),
.B(n_2234),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2286),
.Y(n_2479)
);

NAND3xp33_ASAP7_75t_SL g2480 ( 
.A(n_2312),
.B(n_2069),
.C(n_2093),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2345),
.B(n_2207),
.Y(n_2481)
);

NAND2xp33_ASAP7_75t_R g2482 ( 
.A(n_2333),
.B(n_2225),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2296),
.Y(n_2483)
);

AOI22xp33_ASAP7_75t_L g2484 ( 
.A1(n_2279),
.A2(n_2123),
.B1(n_2183),
.B2(n_2192),
.Y(n_2484)
);

OR2x2_ASAP7_75t_L g2485 ( 
.A(n_2277),
.B(n_2197),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2303),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2306),
.Y(n_2487)
);

INVxp67_ASAP7_75t_L g2488 ( 
.A(n_2365),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2311),
.Y(n_2489)
);

OAI21xp5_ASAP7_75t_SL g2490 ( 
.A1(n_2297),
.A2(n_2222),
.B(n_2154),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_2263),
.Y(n_2491)
);

CKINVDCx5p33_ASAP7_75t_R g2492 ( 
.A(n_2260),
.Y(n_2492)
);

BUFx12f_ASAP7_75t_L g2493 ( 
.A(n_2322),
.Y(n_2493)
);

NAND2xp33_ASAP7_75t_R g2494 ( 
.A(n_2264),
.B(n_2154),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2322),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2314),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2291),
.Y(n_2497)
);

OR2x6_ASAP7_75t_L g2498 ( 
.A(n_2268),
.B(n_2202),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2376),
.B(n_2207),
.Y(n_2499)
);

OR2x2_ASAP7_75t_L g2500 ( 
.A(n_2277),
.B(n_2053),
.Y(n_2500)
);

CKINVDCx20_ASAP7_75t_R g2501 ( 
.A(n_2362),
.Y(n_2501)
);

NAND2xp33_ASAP7_75t_R g2502 ( 
.A(n_2365),
.B(n_2313),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2380),
.Y(n_2503)
);

BUFx6f_ASAP7_75t_L g2504 ( 
.A(n_2395),
.Y(n_2504)
);

NOR2x1_ASAP7_75t_R g2505 ( 
.A(n_2295),
.B(n_2170),
.Y(n_2505)
);

OR2x6_ASAP7_75t_L g2506 ( 
.A(n_2310),
.B(n_2202),
.Y(n_2506)
);

OR2x2_ASAP7_75t_L g2507 ( 
.A(n_2408),
.B(n_2388),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2316),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2352),
.B(n_2192),
.Y(n_2509)
);

AOI21xp5_ASAP7_75t_L g2510 ( 
.A1(n_2359),
.A2(n_2086),
.B(n_2072),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2391),
.B(n_2149),
.Y(n_2511)
);

AO31x2_ASAP7_75t_L g2512 ( 
.A1(n_2364),
.A2(n_2159),
.A3(n_2064),
.B(n_2182),
.Y(n_2512)
);

NOR3xp33_ASAP7_75t_SL g2513 ( 
.A(n_2402),
.B(n_2128),
.C(n_2149),
.Y(n_2513)
);

BUFx3_ASAP7_75t_L g2514 ( 
.A(n_2270),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2367),
.B(n_2202),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2357),
.B(n_2220),
.Y(n_2516)
);

NAND2xp33_ASAP7_75t_R g2517 ( 
.A(n_2337),
.B(n_2274),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2392),
.B(n_2209),
.Y(n_2518)
);

AO32x2_ASAP7_75t_L g2519 ( 
.A1(n_2383),
.A2(n_2250),
.A3(n_2242),
.B1(n_2059),
.B2(n_2018),
.Y(n_2519)
);

AOI22xp33_ASAP7_75t_L g2520 ( 
.A1(n_2289),
.A2(n_2090),
.B1(n_2087),
.B2(n_2186),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_2436),
.Y(n_2521)
);

NAND2xp33_ASAP7_75t_R g2522 ( 
.A(n_2337),
.B(n_2274),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2301),
.Y(n_2523)
);

NAND3xp33_ASAP7_75t_SL g2524 ( 
.A(n_2297),
.B(n_2197),
.C(n_2051),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2317),
.Y(n_2525)
);

NOR2x1p5_ASAP7_75t_L g2526 ( 
.A(n_2304),
.B(n_2173),
.Y(n_2526)
);

AO21x2_ASAP7_75t_L g2527 ( 
.A1(n_2328),
.A2(n_2250),
.B(n_2242),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_2294),
.Y(n_2528)
);

CKINVDCx20_ASAP7_75t_R g2529 ( 
.A(n_2420),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2320),
.B(n_2209),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2325),
.Y(n_2531)
);

CKINVDCx16_ASAP7_75t_R g2532 ( 
.A(n_2309),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_2308),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_L g2534 ( 
.A(n_2356),
.B(n_2152),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_R g2535 ( 
.A(n_2308),
.B(n_2152),
.Y(n_2535)
);

NOR3xp33_ASAP7_75t_SL g2536 ( 
.A(n_2282),
.B(n_2128),
.C(n_2017),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_2256),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_2353),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2327),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2421),
.B(n_2173),
.Y(n_2540)
);

O2A1O1Ixp33_ASAP7_75t_SL g2541 ( 
.A1(n_2262),
.A2(n_2143),
.B(n_2200),
.C(n_1992),
.Y(n_2541)
);

CKINVDCx5p33_ASAP7_75t_R g2542 ( 
.A(n_2353),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2329),
.B(n_2090),
.Y(n_2543)
);

NAND3xp33_ASAP7_75t_SL g2544 ( 
.A(n_2288),
.B(n_2385),
.C(n_2262),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2300),
.Y(n_2545)
);

CKINVDCx14_ASAP7_75t_R g2546 ( 
.A(n_2305),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2336),
.Y(n_2547)
);

AOI22xp33_ASAP7_75t_L g2548 ( 
.A1(n_2331),
.A2(n_2087),
.B1(n_2186),
.B2(n_2017),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2363),
.B(n_2377),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2398),
.B(n_2121),
.Y(n_2550)
);

OR2x2_ASAP7_75t_L g2551 ( 
.A(n_2386),
.B(n_2439),
.Y(n_2551)
);

AOI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2370),
.A2(n_2122),
.B1(n_2086),
.B2(n_2116),
.Y(n_2552)
);

A2O1A1Ixp33_ASAP7_75t_L g2553 ( 
.A1(n_2343),
.A2(n_2385),
.B(n_2407),
.C(n_2417),
.Y(n_2553)
);

AND2x2_ASAP7_75t_SL g2554 ( 
.A(n_2324),
.B(n_2178),
.Y(n_2554)
);

NAND2xp33_ASAP7_75t_R g2555 ( 
.A(n_2337),
.B(n_2100),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2355),
.A2(n_2358),
.B1(n_2319),
.B2(n_2321),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_2340),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2338),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2344),
.Y(n_2559)
);

NAND2xp33_ASAP7_75t_SL g2560 ( 
.A(n_2324),
.B(n_2302),
.Y(n_2560)
);

BUFx3_ASAP7_75t_L g2561 ( 
.A(n_2299),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2366),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2293),
.Y(n_2563)
);

CKINVDCx5p33_ASAP7_75t_R g2564 ( 
.A(n_2374),
.Y(n_2564)
);

HB1xp67_ASAP7_75t_L g2565 ( 
.A(n_2351),
.Y(n_2565)
);

OR2x2_ASAP7_75t_L g2566 ( 
.A(n_2439),
.B(n_2178),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2379),
.B(n_2178),
.Y(n_2567)
);

INVxp67_ASAP7_75t_L g2568 ( 
.A(n_2326),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_R g2569 ( 
.A(n_2395),
.B(n_2160),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2372),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_2396),
.B(n_2375),
.Y(n_2571)
);

HB1xp67_ASAP7_75t_L g2572 ( 
.A(n_2351),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2384),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_R g2574 ( 
.A(n_2299),
.B(n_2160),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_2299),
.Y(n_2575)
);

OAI21xp5_ASAP7_75t_L g2576 ( 
.A1(n_2425),
.A2(n_2032),
.B(n_2002),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2389),
.Y(n_2577)
);

INVxp67_ASAP7_75t_L g2578 ( 
.A(n_2435),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2431),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2323),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2335),
.B(n_2059),
.Y(n_2581)
);

HB1xp67_ASAP7_75t_L g2582 ( 
.A(n_2387),
.Y(n_2582)
);

AO31x2_ASAP7_75t_L g2583 ( 
.A1(n_2394),
.A2(n_2062),
.A3(n_2122),
.B(n_1992),
.Y(n_2583)
);

AO31x2_ASAP7_75t_L g2584 ( 
.A1(n_2394),
.A2(n_2062),
.A3(n_1987),
.B(n_2002),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2346),
.Y(n_2585)
);

AOI22xp33_ASAP7_75t_L g2586 ( 
.A1(n_2269),
.A2(n_2084),
.B1(n_1987),
.B2(n_2007),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2348),
.Y(n_2587)
);

INVx8_ASAP7_75t_L g2588 ( 
.A(n_2428),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2349),
.Y(n_2589)
);

BUFx4f_ASAP7_75t_SL g2590 ( 
.A(n_2433),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2550),
.B(n_2464),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2441),
.Y(n_2592)
);

INVx3_ASAP7_75t_L g2593 ( 
.A(n_2554),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2459),
.B(n_2387),
.Y(n_2594)
);

AOI22xp33_ASAP7_75t_L g2595 ( 
.A1(n_2544),
.A2(n_2343),
.B1(n_2332),
.B2(n_2292),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2442),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2456),
.Y(n_2597)
);

OAI21xp5_ASAP7_75t_SL g2598 ( 
.A1(n_2451),
.A2(n_2288),
.B(n_2272),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2444),
.B(n_2301),
.Y(n_2599)
);

A2O1A1Ixp33_ASAP7_75t_L g2600 ( 
.A1(n_2553),
.A2(n_2292),
.B(n_2417),
.C(n_2332),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2452),
.B(n_2381),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2465),
.B(n_2440),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2449),
.B(n_2432),
.Y(n_2603)
);

BUFx6f_ASAP7_75t_L g2604 ( 
.A(n_2443),
.Y(n_2604)
);

AOI221xp5_ASAP7_75t_L g2605 ( 
.A1(n_2474),
.A2(n_2383),
.B1(n_2382),
.B2(n_2409),
.C(n_2427),
.Y(n_2605)
);

HB1xp67_ASAP7_75t_L g2606 ( 
.A(n_2565),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2457),
.Y(n_2607)
);

HB1xp67_ASAP7_75t_L g2608 ( 
.A(n_2572),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2469),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2549),
.B(n_2428),
.Y(n_2610)
);

OR2x2_ASAP7_75t_L g2611 ( 
.A(n_2507),
.B(n_2307),
.Y(n_2611)
);

HB1xp67_ASAP7_75t_L g2612 ( 
.A(n_2582),
.Y(n_2612)
);

OR2x2_ASAP7_75t_L g2613 ( 
.A(n_2551),
.B(n_2307),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2473),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2479),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2483),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2486),
.Y(n_2617)
);

BUFx6f_ASAP7_75t_L g2618 ( 
.A(n_2443),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2487),
.Y(n_2619)
);

INVx4_ASAP7_75t_L g2620 ( 
.A(n_2466),
.Y(n_2620)
);

INVx4_ASAP7_75t_L g2621 ( 
.A(n_2443),
.Y(n_2621)
);

AND2x4_ASAP7_75t_L g2622 ( 
.A(n_2523),
.B(n_2397),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_L g2623 ( 
.A1(n_2481),
.A2(n_2330),
.B1(n_2406),
.B2(n_2426),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2489),
.B(n_2401),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2496),
.Y(n_2625)
);

HB1xp67_ASAP7_75t_L g2626 ( 
.A(n_2512),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2508),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2525),
.Y(n_2628)
);

AOI22xp33_ASAP7_75t_L g2629 ( 
.A1(n_2448),
.A2(n_2330),
.B1(n_2426),
.B2(n_2354),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2531),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2539),
.Y(n_2631)
);

BUFx2_ASAP7_75t_L g2632 ( 
.A(n_2569),
.Y(n_2632)
);

HB1xp67_ASAP7_75t_L g2633 ( 
.A(n_2512),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2512),
.Y(n_2634)
);

INVx3_ASAP7_75t_L g2635 ( 
.A(n_2588),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2547),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_L g2637 ( 
.A(n_2461),
.B(n_2467),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2558),
.Y(n_2638)
);

BUFx3_ASAP7_75t_L g2639 ( 
.A(n_2504),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2571),
.B(n_2429),
.Y(n_2640)
);

BUFx2_ASAP7_75t_L g2641 ( 
.A(n_2458),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2540),
.B(n_2430),
.Y(n_2642)
);

HB1xp67_ASAP7_75t_L g2643 ( 
.A(n_2555),
.Y(n_2643)
);

BUFx2_ASAP7_75t_L g2644 ( 
.A(n_2535),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2559),
.B(n_2401),
.Y(n_2645)
);

CKINVDCx20_ASAP7_75t_R g2646 ( 
.A(n_2529),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2579),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2499),
.B(n_2334),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2562),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2509),
.B(n_2399),
.Y(n_2650)
);

AND2x4_ASAP7_75t_L g2651 ( 
.A(n_2478),
.B(n_2403),
.Y(n_2651)
);

BUFx2_ASAP7_75t_L g2652 ( 
.A(n_2574),
.Y(n_2652)
);

AOI22xp33_ASAP7_75t_L g2653 ( 
.A1(n_2448),
.A2(n_2266),
.B1(n_2424),
.B2(n_2290),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2570),
.Y(n_2654)
);

INVx5_ASAP7_75t_SL g2655 ( 
.A(n_2454),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2577),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2585),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2516),
.B(n_2567),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2587),
.Y(n_2659)
);

INVx2_ASAP7_75t_SL g2660 ( 
.A(n_2588),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2589),
.Y(n_2661)
);

HB1xp67_ASAP7_75t_L g2662 ( 
.A(n_2497),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2485),
.Y(n_2663)
);

NOR2x1_ASAP7_75t_SL g2664 ( 
.A(n_2466),
.B(n_2347),
.Y(n_2664)
);

INVxp67_ASAP7_75t_L g2665 ( 
.A(n_2472),
.Y(n_2665)
);

OR2x2_ASAP7_75t_L g2666 ( 
.A(n_2500),
.B(n_2405),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2460),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2455),
.Y(n_2668)
);

HB1xp67_ASAP7_75t_L g2669 ( 
.A(n_2545),
.Y(n_2669)
);

INVx3_ASAP7_75t_L g2670 ( 
.A(n_2504),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2502),
.A2(n_2276),
.B1(n_2424),
.B2(n_2285),
.Y(n_2671)
);

INVx8_ASAP7_75t_L g2672 ( 
.A(n_2504),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_2580),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2543),
.Y(n_2674)
);

OR2x2_ASAP7_75t_L g2675 ( 
.A(n_2532),
.B(n_2405),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2511),
.Y(n_2676)
);

AND2x4_ASAP7_75t_L g2677 ( 
.A(n_2530),
.B(n_2415),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2518),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2581),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2597),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2592),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2648),
.B(n_2527),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2679),
.B(n_2676),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2663),
.B(n_2556),
.Y(n_2684)
);

HB1xp67_ASAP7_75t_L g2685 ( 
.A(n_2606),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2674),
.B(n_2552),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2592),
.Y(n_2687)
);

AND2x4_ASAP7_75t_L g2688 ( 
.A(n_2591),
.B(n_2438),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2651),
.B(n_2678),
.Y(n_2689)
);

HB1xp67_ASAP7_75t_L g2690 ( 
.A(n_2606),
.Y(n_2690)
);

INVxp67_ASAP7_75t_SL g2691 ( 
.A(n_2662),
.Y(n_2691)
);

HB1xp67_ASAP7_75t_L g2692 ( 
.A(n_2608),
.Y(n_2692)
);

AND2x4_ASAP7_75t_L g2693 ( 
.A(n_2591),
.B(n_2510),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2667),
.B(n_2484),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2651),
.B(n_2411),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2651),
.B(n_2519),
.Y(n_2696)
);

OR2x2_ASAP7_75t_L g2697 ( 
.A(n_2611),
.B(n_2566),
.Y(n_2697)
);

INVx2_ASAP7_75t_SL g2698 ( 
.A(n_2652),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2650),
.B(n_2446),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2668),
.B(n_2534),
.Y(n_2700)
);

AND2x4_ASAP7_75t_L g2701 ( 
.A(n_2591),
.B(n_2643),
.Y(n_2701)
);

AOI211xp5_ASAP7_75t_L g2702 ( 
.A1(n_2598),
.A2(n_2505),
.B(n_2560),
.C(n_2488),
.Y(n_2702)
);

AND2x2_ASAP7_75t_L g2703 ( 
.A(n_2650),
.B(n_2520),
.Y(n_2703)
);

HB1xp67_ASAP7_75t_L g2704 ( 
.A(n_2608),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2650),
.B(n_2584),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2622),
.B(n_2584),
.Y(n_2706)
);

OR2x2_ASAP7_75t_L g2707 ( 
.A(n_2613),
.B(n_2476),
.Y(n_2707)
);

NAND2x1p5_ASAP7_75t_L g2708 ( 
.A(n_2620),
.B(n_2526),
.Y(n_2708)
);

OAI21xp5_ASAP7_75t_L g2709 ( 
.A1(n_2600),
.A2(n_2524),
.B(n_2536),
.Y(n_2709)
);

AND2x4_ASAP7_75t_SL g2710 ( 
.A(n_2620),
.B(n_2454),
.Y(n_2710)
);

AND3x2_ASAP7_75t_L g2711 ( 
.A(n_2641),
.B(n_2568),
.C(n_2578),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2622),
.B(n_2658),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2637),
.B(n_2470),
.Y(n_2713)
);

HB1xp67_ASAP7_75t_L g2714 ( 
.A(n_2612),
.Y(n_2714)
);

OR2x2_ASAP7_75t_L g2715 ( 
.A(n_2666),
.B(n_2584),
.Y(n_2715)
);

NOR3xp33_ASAP7_75t_L g2716 ( 
.A(n_2600),
.B(n_2515),
.C(n_2480),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2622),
.B(n_2368),
.Y(n_2717)
);

OR2x2_ASAP7_75t_L g2718 ( 
.A(n_2612),
.B(n_2675),
.Y(n_2718)
);

HB1xp67_ASAP7_75t_L g2719 ( 
.A(n_2662),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2677),
.B(n_2576),
.Y(n_2720)
);

OR2x2_ASAP7_75t_L g2721 ( 
.A(n_2624),
.B(n_2548),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2677),
.B(n_2583),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_2669),
.Y(n_2723)
);

AND3x1_ASAP7_75t_L g2724 ( 
.A(n_2702),
.B(n_2635),
.C(n_2660),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2682),
.B(n_2643),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2682),
.B(n_2677),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_SL g2727 ( 
.A(n_2702),
.B(n_2644),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2681),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2681),
.Y(n_2729)
);

INVxp67_ASAP7_75t_SL g2730 ( 
.A(n_2719),
.Y(n_2730)
);

AND2x4_ASAP7_75t_L g2731 ( 
.A(n_2701),
.B(n_2665),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2687),
.Y(n_2732)
);

HB1xp67_ASAP7_75t_L g2733 ( 
.A(n_2723),
.Y(n_2733)
);

AND2x4_ASAP7_75t_SL g2734 ( 
.A(n_2698),
.B(n_2620),
.Y(n_2734)
);

AND2x4_ASAP7_75t_L g2735 ( 
.A(n_2701),
.B(n_2665),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2720),
.B(n_2623),
.Y(n_2736)
);

NAND4xp25_ASAP7_75t_L g2737 ( 
.A(n_2716),
.B(n_2629),
.C(n_2595),
.D(n_2623),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2720),
.B(n_2626),
.Y(n_2738)
);

INVxp67_ASAP7_75t_L g2739 ( 
.A(n_2698),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2689),
.B(n_2626),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2689),
.B(n_2633),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2701),
.Y(n_2742)
);

OR2x2_ASAP7_75t_L g2743 ( 
.A(n_2718),
.B(n_2645),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2696),
.B(n_2633),
.Y(n_2744)
);

INVxp33_ASAP7_75t_L g2745 ( 
.A(n_2708),
.Y(n_2745)
);

INVx2_ASAP7_75t_L g2746 ( 
.A(n_2680),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2696),
.B(n_2610),
.Y(n_2747)
);

AND2x4_ASAP7_75t_L g2748 ( 
.A(n_2701),
.B(n_2634),
.Y(n_2748)
);

NAND5xp2_ASAP7_75t_L g2749 ( 
.A(n_2709),
.B(n_2629),
.C(n_2595),
.D(n_2605),
.E(n_2653),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2684),
.B(n_2637),
.Y(n_2750)
);

INVx3_ASAP7_75t_L g2751 ( 
.A(n_2688),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2688),
.B(n_2669),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2695),
.B(n_2640),
.Y(n_2753)
);

OR2x2_ASAP7_75t_L g2754 ( 
.A(n_2718),
.B(n_2673),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2695),
.B(n_2594),
.Y(n_2755)
);

OR2x2_ASAP7_75t_L g2756 ( 
.A(n_2685),
.B(n_2673),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2705),
.B(n_2596),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2683),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2683),
.Y(n_2759)
);

NOR3xp33_ASAP7_75t_SL g2760 ( 
.A(n_2709),
.B(n_2447),
.C(n_2445),
.Y(n_2760)
);

BUFx2_ASAP7_75t_L g2761 ( 
.A(n_2724),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2754),
.Y(n_2762)
);

XNOR2xp5_ASAP7_75t_L g2763 ( 
.A(n_2760),
.B(n_2475),
.Y(n_2763)
);

AOI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_2737),
.A2(n_2713),
.B1(n_2703),
.B2(n_2699),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2754),
.Y(n_2765)
);

OR2x2_ASAP7_75t_L g2766 ( 
.A(n_2743),
.B(n_2758),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_R g2767 ( 
.A(n_2736),
.B(n_2671),
.Y(n_2767)
);

AOI22xp33_ASAP7_75t_L g2768 ( 
.A1(n_2749),
.A2(n_2700),
.B1(n_2601),
.B2(n_2699),
.Y(n_2768)
);

AND2x4_ASAP7_75t_L g2769 ( 
.A(n_2731),
.B(n_2735),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2756),
.Y(n_2770)
);

OR2x2_ASAP7_75t_L g2771 ( 
.A(n_2743),
.B(n_2697),
.Y(n_2771)
);

O2A1O1Ixp5_ASAP7_75t_R g2772 ( 
.A1(n_2750),
.A2(n_2694),
.B(n_2603),
.C(n_2599),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2731),
.B(n_2712),
.Y(n_2773)
);

AOI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2727),
.A2(n_2703),
.B1(n_2686),
.B2(n_2710),
.Y(n_2774)
);

OR2x2_ASAP7_75t_L g2775 ( 
.A(n_2758),
.B(n_2697),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2733),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2734),
.B(n_2688),
.Y(n_2777)
);

HB1xp67_ASAP7_75t_L g2778 ( 
.A(n_2756),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2757),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2746),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2757),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2730),
.Y(n_2782)
);

OAI33xp33_ASAP7_75t_L g2783 ( 
.A1(n_2739),
.A2(n_2471),
.A3(n_2468),
.B1(n_2721),
.B2(n_2707),
.B3(n_2617),
.Y(n_2783)
);

AOI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2736),
.A2(n_2686),
.B1(n_2710),
.B2(n_2705),
.Y(n_2784)
);

AOI21x1_ASAP7_75t_L g2785 ( 
.A1(n_2742),
.A2(n_2632),
.B(n_2690),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2746),
.Y(n_2786)
);

NOR2xp67_ASAP7_75t_L g2787 ( 
.A(n_2751),
.B(n_2493),
.Y(n_2787)
);

INVx2_ASAP7_75t_SL g2788 ( 
.A(n_2734),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2759),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2731),
.B(n_2712),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2740),
.A2(n_2710),
.B1(n_2706),
.B2(n_2717),
.Y(n_2791)
);

NAND2xp33_ASAP7_75t_L g2792 ( 
.A(n_2745),
.B(n_2708),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2759),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2735),
.B(n_2692),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2744),
.B(n_2704),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2740),
.Y(n_2796)
);

NOR2xp67_ASAP7_75t_L g2797 ( 
.A(n_2751),
.B(n_2621),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2744),
.B(n_2714),
.Y(n_2798)
);

AOI21xp5_ASAP7_75t_L g2799 ( 
.A1(n_2752),
.A2(n_2541),
.B(n_2664),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2741),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2741),
.Y(n_2801)
);

AOI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2783),
.A2(n_2725),
.B1(n_2738),
.B2(n_2735),
.Y(n_2802)
);

OR2x2_ASAP7_75t_L g2803 ( 
.A(n_2771),
.B(n_2738),
.Y(n_2803)
);

OAI22xp33_ASAP7_75t_L g2804 ( 
.A1(n_2774),
.A2(n_2742),
.B1(n_2751),
.B2(n_2708),
.Y(n_2804)
);

NOR3xp33_ASAP7_75t_L g2805 ( 
.A(n_2783),
.B(n_2761),
.C(n_2772),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2778),
.Y(n_2806)
);

HB1xp67_ASAP7_75t_L g2807 ( 
.A(n_2778),
.Y(n_2807)
);

AOI221xp5_ASAP7_75t_L g2808 ( 
.A1(n_2768),
.A2(n_2725),
.B1(n_2627),
.B2(n_2619),
.C(n_2616),
.Y(n_2808)
);

NAND3xp33_ASAP7_75t_L g2809 ( 
.A(n_2764),
.B(n_2711),
.C(n_2513),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2794),
.B(n_2747),
.Y(n_2810)
);

O2A1O1Ixp33_ASAP7_75t_L g2811 ( 
.A1(n_2776),
.A2(n_2546),
.B(n_2501),
.C(n_2477),
.Y(n_2811)
);

OAI22xp33_ASAP7_75t_SL g2812 ( 
.A1(n_2777),
.A2(n_2752),
.B1(n_2593),
.B2(n_2660),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2766),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2785),
.Y(n_2814)
);

NAND3xp33_ASAP7_75t_L g2815 ( 
.A(n_2768),
.B(n_2653),
.C(n_2721),
.Y(n_2815)
);

NOR3xp33_ASAP7_75t_L g2816 ( 
.A(n_2777),
.B(n_2782),
.C(n_2792),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2795),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2795),
.Y(n_2818)
);

AOI21xp33_ASAP7_75t_L g2819 ( 
.A1(n_2763),
.A2(n_2537),
.B(n_2563),
.Y(n_2819)
);

AOI221xp5_ASAP7_75t_L g2820 ( 
.A1(n_2762),
.A2(n_2654),
.B1(n_2614),
.B2(n_2615),
.C(n_2625),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2798),
.Y(n_2821)
);

AOI22x1_ASAP7_75t_SL g2822 ( 
.A1(n_2767),
.A2(n_2646),
.B1(n_2495),
.B2(n_2533),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2798),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2775),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2779),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2780),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2781),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_2822),
.B(n_2646),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2807),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2826),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2817),
.B(n_2818),
.Y(n_2831)
);

NOR2x1_ASAP7_75t_L g2832 ( 
.A(n_2814),
.B(n_2491),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2808),
.B(n_2796),
.Y(n_2833)
);

O2A1O1Ixp33_ASAP7_75t_L g2834 ( 
.A1(n_2805),
.A2(n_2788),
.B(n_2450),
.C(n_2453),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2824),
.Y(n_2835)
);

AOI21xp33_ASAP7_75t_L g2836 ( 
.A1(n_2815),
.A2(n_2437),
.B(n_2492),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2813),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2803),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2806),
.Y(n_2839)
);

OAI31xp33_ASAP7_75t_L g2840 ( 
.A1(n_2812),
.A2(n_2769),
.A3(n_2799),
.B(n_2752),
.Y(n_2840)
);

NOR2xp33_ASAP7_75t_L g2841 ( 
.A(n_2819),
.B(n_2528),
.Y(n_2841)
);

NOR2xp33_ASAP7_75t_L g2842 ( 
.A(n_2819),
.B(n_2769),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_2825),
.Y(n_2843)
);

XNOR2x1_ASAP7_75t_L g2844 ( 
.A(n_2809),
.B(n_2503),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2808),
.B(n_2800),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2821),
.Y(n_2846)
);

OAI221xp5_ASAP7_75t_L g2847 ( 
.A1(n_2816),
.A2(n_2802),
.B1(n_2784),
.B2(n_2791),
.C(n_2811),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2823),
.B(n_2820),
.Y(n_2848)
);

INVxp67_ASAP7_75t_L g2849 ( 
.A(n_2820),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2827),
.B(n_2789),
.Y(n_2850)
);

OAI221xp5_ASAP7_75t_L g2851 ( 
.A1(n_2804),
.A2(n_2797),
.B1(n_2787),
.B2(n_2799),
.C(n_2770),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_SL g2852 ( 
.A(n_2810),
.B(n_2693),
.Y(n_2852)
);

AND2x4_ASAP7_75t_L g2853 ( 
.A(n_2816),
.B(n_2773),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_L g2854 ( 
.A(n_2822),
.B(n_2790),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2807),
.Y(n_2855)
);

OAI21xp33_ASAP7_75t_L g2856 ( 
.A1(n_2847),
.A2(n_2765),
.B(n_2793),
.Y(n_2856)
);

NAND3xp33_ASAP7_75t_L g2857 ( 
.A(n_2840),
.B(n_2557),
.C(n_2564),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2829),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2855),
.Y(n_2859)
);

NOR3x1_ASAP7_75t_L g2860 ( 
.A(n_2851),
.B(n_2848),
.C(n_2845),
.Y(n_2860)
);

AOI211xp5_ASAP7_75t_L g2861 ( 
.A1(n_2834),
.A2(n_2538),
.B(n_2542),
.C(n_2463),
.Y(n_2861)
);

NAND3xp33_ASAP7_75t_SL g2862 ( 
.A(n_2828),
.B(n_2573),
.C(n_2272),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2849),
.B(n_2753),
.Y(n_2863)
);

NOR2xp33_ASAP7_75t_L g2864 ( 
.A(n_2844),
.B(n_2462),
.Y(n_2864)
);

NAND3xp33_ASAP7_75t_L g2865 ( 
.A(n_2836),
.B(n_2514),
.C(n_2586),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2848),
.B(n_2753),
.Y(n_2866)
);

NAND3xp33_ASAP7_75t_L g2867 ( 
.A(n_2836),
.B(n_2786),
.C(n_2729),
.Y(n_2867)
);

NOR2x1_ASAP7_75t_L g2868 ( 
.A(n_2832),
.B(n_2635),
.Y(n_2868)
);

AOI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_2854),
.A2(n_2672),
.B(n_2521),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2835),
.B(n_2747),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2831),
.Y(n_2871)
);

NOR2x1_ASAP7_75t_SL g2872 ( 
.A(n_2852),
.B(n_2621),
.Y(n_2872)
);

NAND2x1p5_ASAP7_75t_L g2873 ( 
.A(n_2841),
.B(n_2561),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2831),
.Y(n_2874)
);

NAND3xp33_ASAP7_75t_L g2875 ( 
.A(n_2842),
.B(n_2729),
.C(n_2728),
.Y(n_2875)
);

AOI221xp5_ASAP7_75t_L g2876 ( 
.A1(n_2833),
.A2(n_2801),
.B1(n_2726),
.B2(n_2722),
.C(n_2656),
.Y(n_2876)
);

NOR2x1_ASAP7_75t_L g2877 ( 
.A(n_2857),
.B(n_2853),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2862),
.A2(n_2853),
.B(n_2839),
.Y(n_2878)
);

NAND3xp33_ASAP7_75t_L g2879 ( 
.A(n_2856),
.B(n_2846),
.C(n_2837),
.Y(n_2879)
);

AOI21xp5_ASAP7_75t_L g2880 ( 
.A1(n_2869),
.A2(n_2850),
.B(n_2843),
.Y(n_2880)
);

OAI22xp5_ASAP7_75t_L g2881 ( 
.A1(n_2866),
.A2(n_2838),
.B1(n_2830),
.B2(n_2850),
.Y(n_2881)
);

NOR2xp33_ASAP7_75t_L g2882 ( 
.A(n_2864),
.B(n_2590),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2858),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2859),
.Y(n_2884)
);

HB1xp67_ASAP7_75t_L g2885 ( 
.A(n_2871),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_SL g2886 ( 
.A(n_2868),
.B(n_2655),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_SL g2887 ( 
.A(n_2861),
.B(n_2655),
.Y(n_2887)
);

OA22x2_ASAP7_75t_L g2888 ( 
.A1(n_2874),
.A2(n_2693),
.B1(n_2276),
.B2(n_2688),
.Y(n_2888)
);

AOI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2861),
.A2(n_2672),
.B(n_2413),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2863),
.B(n_2655),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2876),
.B(n_2755),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_SL g2892 ( 
.A(n_2867),
.B(n_2604),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2860),
.B(n_2755),
.Y(n_2893)
);

OAI221xp5_ASAP7_75t_SL g2894 ( 
.A1(n_2893),
.A2(n_2875),
.B1(n_2865),
.B2(n_2870),
.C(n_2506),
.Y(n_2894)
);

AOI221xp5_ASAP7_75t_L g2895 ( 
.A1(n_2885),
.A2(n_2884),
.B1(n_2883),
.B2(n_2878),
.C(n_2879),
.Y(n_2895)
);

NOR2xp67_ASAP7_75t_L g2896 ( 
.A(n_2880),
.B(n_2872),
.Y(n_2896)
);

NAND3xp33_ASAP7_75t_L g2897 ( 
.A(n_2877),
.B(n_2423),
.C(n_2422),
.Y(n_2897)
);

AOI221xp5_ASAP7_75t_L g2898 ( 
.A1(n_2881),
.A2(n_2873),
.B1(n_2649),
.B2(n_2607),
.C(n_2628),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2892),
.Y(n_2899)
);

AOI21xp5_ASAP7_75t_L g2900 ( 
.A1(n_2887),
.A2(n_2886),
.B(n_2882),
.Y(n_2900)
);

AOI221xp5_ASAP7_75t_L g2901 ( 
.A1(n_2890),
.A2(n_2638),
.B1(n_2636),
.B2(n_2630),
.C(n_2609),
.Y(n_2901)
);

NAND3xp33_ASAP7_75t_L g2902 ( 
.A(n_2891),
.B(n_2889),
.C(n_2888),
.Y(n_2902)
);

XNOR2x1_ASAP7_75t_L g2903 ( 
.A(n_2877),
.B(n_2506),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2877),
.B(n_2726),
.Y(n_2904)
);

NOR3xp33_ASAP7_75t_L g2905 ( 
.A(n_2877),
.B(n_2416),
.C(n_2404),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2893),
.B(n_2722),
.Y(n_2906)
);

AOI221xp5_ASAP7_75t_SL g2907 ( 
.A1(n_2878),
.A2(n_2631),
.B1(n_2647),
.B2(n_2691),
.C(n_2707),
.Y(n_2907)
);

AOI221xp5_ASAP7_75t_SL g2908 ( 
.A1(n_2878),
.A2(n_2657),
.B1(n_2659),
.B2(n_2661),
.C(n_2642),
.Y(n_2908)
);

NOR2x1_ASAP7_75t_L g2909 ( 
.A(n_2903),
.B(n_2498),
.Y(n_2909)
);

AO22x1_ASAP7_75t_L g2910 ( 
.A1(n_2905),
.A2(n_2639),
.B1(n_2414),
.B2(n_2575),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2902),
.B(n_2414),
.Y(n_2911)
);

OR2x2_ASAP7_75t_L g2912 ( 
.A(n_2906),
.B(n_2715),
.Y(n_2912)
);

AOI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2896),
.A2(n_2517),
.B1(n_2522),
.B2(n_2693),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2899),
.Y(n_2914)
);

INVxp67_ASAP7_75t_L g2915 ( 
.A(n_2897),
.Y(n_2915)
);

AOI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2904),
.A2(n_2693),
.B1(n_2482),
.B2(n_2494),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2901),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2898),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_2895),
.B(n_2604),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2894),
.Y(n_2920)
);

HB1xp67_ASAP7_75t_L g2921 ( 
.A(n_2914),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2911),
.B(n_2900),
.Y(n_2922)
);

OAI321xp33_ASAP7_75t_L g2923 ( 
.A1(n_2920),
.A2(n_2907),
.A3(n_2908),
.B1(n_2371),
.B2(n_2281),
.C(n_2419),
.Y(n_2923)
);

NOR2x1_ASAP7_75t_L g2924 ( 
.A(n_2919),
.B(n_2498),
.Y(n_2924)
);

NOR3xp33_ASAP7_75t_L g2925 ( 
.A(n_2910),
.B(n_2404),
.C(n_2400),
.Y(n_2925)
);

AOI221xp5_ASAP7_75t_SL g2926 ( 
.A1(n_2915),
.A2(n_2918),
.B1(n_2917),
.B2(n_2909),
.C(n_2912),
.Y(n_2926)
);

AOI21xp5_ASAP7_75t_L g2927 ( 
.A1(n_2913),
.A2(n_2413),
.B(n_2672),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2916),
.B(n_2728),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2914),
.Y(n_2929)
);

OAI211xp5_ASAP7_75t_SL g2930 ( 
.A1(n_2914),
.A2(n_2490),
.B(n_2670),
.C(n_2593),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2914),
.Y(n_2931)
);

AOI211xp5_ASAP7_75t_L g2932 ( 
.A1(n_2920),
.A2(n_2575),
.B(n_2258),
.C(n_2275),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2911),
.B(n_2602),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2921),
.B(n_2732),
.Y(n_2934)
);

CKINVDCx5p33_ASAP7_75t_R g2935 ( 
.A(n_2929),
.Y(n_2935)
);

OR2x2_ASAP7_75t_L g2936 ( 
.A(n_2931),
.B(n_2715),
.Y(n_2936)
);

CKINVDCx20_ASAP7_75t_R g2937 ( 
.A(n_2922),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2932),
.B(n_2732),
.Y(n_2938)
);

INVx1_ASAP7_75t_SL g2939 ( 
.A(n_2924),
.Y(n_2939)
);

CKINVDCx5p33_ASAP7_75t_R g2940 ( 
.A(n_2933),
.Y(n_2940)
);

XOR2xp5_ASAP7_75t_L g2941 ( 
.A(n_2937),
.B(n_2927),
.Y(n_2941)
);

INVxp67_ASAP7_75t_L g2942 ( 
.A(n_2935),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2940),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2939),
.B(n_2923),
.Y(n_2944)
);

OAI22x1_ASAP7_75t_L g2945 ( 
.A1(n_2934),
.A2(n_2926),
.B1(n_2928),
.B2(n_2925),
.Y(n_2945)
);

AOI31xp33_ASAP7_75t_L g2946 ( 
.A1(n_2942),
.A2(n_2936),
.A3(n_2938),
.B(n_2930),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2944),
.A2(n_2433),
.B1(n_2575),
.B2(n_2639),
.Y(n_2947)
);

AOI221xp5_ASAP7_75t_L g2948 ( 
.A1(n_2945),
.A2(n_2410),
.B1(n_2400),
.B2(n_2393),
.C(n_2418),
.Y(n_2948)
);

AOI22xp33_ASAP7_75t_SL g2949 ( 
.A1(n_2943),
.A2(n_2258),
.B1(n_2275),
.B2(n_2618),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2941),
.Y(n_2950)
);

OAI21xp5_ASAP7_75t_SL g2951 ( 
.A1(n_2949),
.A2(n_2371),
.B(n_2281),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2950),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2947),
.B(n_2670),
.Y(n_2953)
);

HB1xp67_ASAP7_75t_L g2954 ( 
.A(n_2952),
.Y(n_2954)
);

OAI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2954),
.A2(n_2946),
.B1(n_2953),
.B2(n_2951),
.Y(n_2955)
);

AOI22xp5_ASAP7_75t_L g2956 ( 
.A1(n_2955),
.A2(n_2948),
.B1(n_2275),
.B2(n_2258),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2956),
.B(n_2410),
.Y(n_2957)
);

AOI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_2957),
.A2(n_2618),
.B1(n_2604),
.B2(n_2748),
.Y(n_2958)
);


endmodule