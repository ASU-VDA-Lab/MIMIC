module fake_jpeg_11892_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_5),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_1),
.B(n_2),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_58),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_50),
.Y(n_63)
);

NOR2xp67_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_3),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_41),
.B1(n_51),
.B2(n_40),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_74),
.B(n_54),
.C(n_44),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_73),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_8),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_54),
.B(n_60),
.C(n_48),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_11),
.B(n_12),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_54),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_3),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_89),
.Y(n_102)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_96)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_76),
.B1(n_78),
.B2(n_83),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_92),
.B1(n_25),
.B2(n_26),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_104),
.B(n_24),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_97),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_85),
.B(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_16),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_23),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_18),
.B(n_19),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_110),
.Y(n_117)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_103),
.B(n_99),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_112),
.B(n_113),
.Y(n_116)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_107),
.B(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_115),
.B1(n_104),
.B2(n_96),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_106),
.B(n_111),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_105),
.B1(n_102),
.B2(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_27),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_123),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_122),
.B(n_119),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_120),
.B(n_30),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_29),
.Y(n_129)
);


endmodule