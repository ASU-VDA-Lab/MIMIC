module fake_jpeg_21390_n_39 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_39);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_32;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_22),
.A2(n_23),
.B1(n_5),
.B2(n_18),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_26),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_30),
.Y(n_32)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2x1_ASAP7_75t_SL g34 ( 
.A(n_33),
.B(n_24),
.Y(n_34)
);

AOI31xp33_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_31),
.A3(n_28),
.B(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_36),
.B(n_32),
.Y(n_37)
);

OAI321xp33_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_30),
.A3(n_19),
.B1(n_14),
.B2(n_8),
.C(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_17),
.B1(n_19),
.B2(n_32),
.Y(n_39)
);


endmodule