module real_jpeg_17793_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_50;
wire n_38;
wire n_29;
wire n_55;
wire n_49;
wire n_52;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_47;
wire n_14;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_53;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_0),
.A2(n_3),
.B(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_2),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_3),
.A2(n_16),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_3),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_19),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_5),
.A2(n_17),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_7),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_9),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

OAI31xp33_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_29),
.A3(n_33),
.B(n_37),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_23),
.Y(n_13)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_24),
.A2(n_27),
.B(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_27),
.C(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_51),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_48),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);


endmodule