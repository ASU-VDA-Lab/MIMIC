module real_jpeg_18163_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_436),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_0),
.B(n_437),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_85),
.B1(n_89),
.B2(n_90),
.Y(n_84)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_1),
.A2(n_89),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22x1_ASAP7_75t_SL g314 ( 
.A1(n_1),
.A2(n_89),
.B1(n_315),
.B2(n_319),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_1),
.A2(n_89),
.B1(n_159),
.B2(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_2),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_2),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_3),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_3),
.A2(n_56),
.B1(n_171),
.B2(n_174),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_4),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_4),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_5),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_5),
.B(n_86),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_5),
.A2(n_26),
.B1(n_156),
.B2(n_159),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_5),
.A2(n_26),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_5),
.B(n_332),
.Y(n_331)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_5),
.A2(n_358),
.A3(n_360),
.B1(n_362),
.B2(n_364),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_5),
.B(n_306),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_5),
.B(n_179),
.Y(n_393)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_6),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_6),
.Y(n_306)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_7),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_7),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_7),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g321 ( 
.A(n_7),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_7),
.Y(n_367)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_8),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_9),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_10),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_10),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_10),
.A2(n_129),
.B1(n_193),
.B2(n_196),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_10),
.A2(n_129),
.B1(n_257),
.B2(n_260),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_12),
.Y(n_161)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_13),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_13),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_409),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_281),
.B(n_405),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_264),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_20),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_240),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_21),
.B(n_240),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_151),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_22),
.B(n_152),
.C(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_82),
.C(n_123),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_23),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_50),
.Y(n_23)
);

XOR2x2_ASAP7_75t_SL g269 ( 
.A(n_24),
.B(n_50),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B1(n_40),
.B2(n_43),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_26),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_26),
.B(n_108),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_26),
.A2(n_40),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_26),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_26),
.B(n_363),
.Y(n_362)
);

OAI32xp33_ASAP7_75t_L g289 ( 
.A1(n_27),
.A2(n_122),
.A3(n_290),
.B1(n_292),
.B2(n_297),
.Y(n_289)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_36),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_39),
.A2(n_134),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_42),
.Y(n_144)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_49),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_63),
.B(n_67),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_51),
.A2(n_73),
.B(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_55),
.Y(n_388)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_66),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_67),
.B(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_68),
.A2(n_154),
.B(n_162),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_69),
.A2(n_234),
.B(n_237),
.Y(n_233)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_73),
.B(n_155),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_73),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_73),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_75),
.Y(n_236)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_77),
.Y(n_187)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_82),
.A2(n_123),
.B1(n_124),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_82),
.Y(n_244)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_119),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_83),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_94),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_84),
.B(n_95),
.Y(n_254)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_109),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_94),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_94),
.B(n_256),
.Y(n_255)
);

NOR2x1p5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_107),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_95),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_95),
.B(n_256),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_95),
.Y(n_332)
);

AO22x2_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B1(n_102),
.B2(n_104),
.Y(n_95)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_102),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_103),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_103),
.Y(n_291)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_106),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_116),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_110),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_114),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_120),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_139),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_126),
.B(n_140),
.Y(n_219)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_129),
.B(n_235),
.Y(n_234)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_132),
.B(n_145),
.Y(n_218)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_132),
.Y(n_275)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_140),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_140),
.Y(n_428)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_145),
.Y(n_427)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_147),
.Y(n_252)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_211),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_168),
.Y(n_152)
);

AOI21x1_ASAP7_75t_L g424 ( 
.A1(n_153),
.A2(n_169),
.B(n_190),
.Y(n_424)
);

OA21x2_ASAP7_75t_L g302 ( 
.A1(n_154),
.A2(n_303),
.B(n_307),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_154),
.A2(n_335),
.B(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_183),
.B1(n_185),
.B2(n_188),
.Y(n_182)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_161),
.Y(n_340)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_161),
.Y(n_361)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp67_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_190),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_179),
.Y(n_169)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_170),
.Y(n_421)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_180),
.B(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_192),
.Y(n_230)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_181),
.A2(n_199),
.B(n_223),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_181),
.B(n_314),
.Y(n_353)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_182),
.B(n_200),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_201),
.B1(n_205),
.B2(n_209),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_186),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_189),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_191),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_199),
.B(n_314),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_199),
.Y(n_422)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_211),
.Y(n_412)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_220),
.Y(n_211)
);

XOR2x1_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_213),
.Y(n_415)
);

AOI21x1_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B(n_216),
.Y(n_213)
);

NOR2x1p5_ASAP7_75t_SL g349 ( 
.A(n_215),
.B(n_216),
.Y(n_349)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_217),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_220),
.B(n_415),
.C(n_416),
.Y(n_414)
);

NAND2x1p5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_231),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_231),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_222),
.B(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_223),
.Y(n_312)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_230),
.B(n_313),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_230),
.A2(n_421),
.B(n_422),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_233),
.B(n_336),
.Y(n_392)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_238),
.Y(n_335)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.C(n_263),
.Y(n_240)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_280),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_263),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.C(n_253),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_248),
.B1(n_253),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_249),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_251),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_254),
.B(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_279),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_265),
.B(n_279),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.C(n_270),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_266),
.B(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_269),
.Y(n_324)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.C(n_276),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_273),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_276),
.B1(n_277),
.B2(n_287),
.Y(n_286)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_274),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_275),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_426)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_278),
.B(n_378),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_325),
.B(n_404),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_322),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_284),
.B(n_322),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.C(n_308),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_285),
.B(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_288),
.A2(n_308),
.B1(n_309),
.B2(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_288),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_302),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_289),
.A2(n_302),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_289),
.Y(n_344)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_302),
.A2(n_343),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx12f_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_398),
.B(n_403),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_354),
.B(n_397),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_341),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_328),
.B(n_341),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.C(n_333),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_372),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_342),
.B(n_347),
.C(n_350),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_350),
.B2(n_351),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_349),
.B(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

AOI21x1_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_374),
.B(n_396),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_371),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_SL g396 ( 
.A(n_356),
.B(n_371),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_370),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_370),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_368),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_382),
.B(n_395),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_381),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_381),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_391),
.B(n_394),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_390),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_389),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_393),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_392),
.B(n_393),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_402),
.Y(n_403)
);

NAND2xp33_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_434),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_411),
.B(n_413),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_423),
.B1(n_432),
.B2(n_433),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_418),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_423),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_430),
.Y(n_425)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);


endmodule