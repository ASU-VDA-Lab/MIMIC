module real_jpeg_31146_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx3_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_0),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_0),
.A2(n_96),
.B1(n_165),
.B2(n_170),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_0),
.A2(n_96),
.B1(n_205),
.B2(n_208),
.Y(n_204)
);

AOI22x1_ASAP7_75t_L g246 ( 
.A1(n_0),
.A2(n_96),
.B1(n_247),
.B2(n_250),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_1),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_1),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_2),
.B(n_288),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_2),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_5),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_5),
.Y(n_199)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_5),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_6),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_6),
.A2(n_50),
.B1(n_228),
.B2(n_231),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_6),
.A2(n_50),
.B1(n_258),
.B2(n_261),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_6),
.A2(n_50),
.B1(n_247),
.B2(n_365),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_7),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_10),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_10),
.A2(n_108),
.B1(n_115),
.B2(n_119),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_10),
.A2(n_108),
.B1(n_197),
.B2(n_200),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_10),
.A2(n_108),
.B1(n_296),
.B2(n_300),
.Y(n_295)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_11),
.Y(n_127)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_12),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_13),
.Y(n_38)
);

OAI22x1_ASAP7_75t_SL g151 ( 
.A1(n_13),
.A2(n_38),
.B1(n_152),
.B2(n_156),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_13),
.A2(n_38),
.B1(n_214),
.B2(n_217),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_13),
.A2(n_38),
.B1(n_329),
.B2(n_331),
.Y(n_328)
);

INVx2_ASAP7_75t_R g355 ( 
.A(n_13),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_13),
.B(n_112),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_13),
.B(n_210),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_SL g431 ( 
.A(n_13),
.B(n_25),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_13),
.B(n_445),
.Y(n_444)
);

OAI311xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_281),
.A3(n_285),
.B1(n_306),
.C1(n_310),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_15),
.A2(n_286),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI21xp33_ASAP7_75t_SL g310 ( 
.A1(n_16),
.A2(n_311),
.B(n_530),
.Y(n_310)
);

AOI21xp33_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_177),
.B(n_279),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_17),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_158),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_18),
.B(n_158),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_141),
.C(n_146),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_20),
.A2(n_21),
.B1(n_141),
.B2(n_142),
.Y(n_275)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_65),
.B2(n_66),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_22),
.A2(n_23),
.B1(n_225),
.B2(n_432),
.Y(n_477)
);

OAI22x1_ASAP7_75t_L g506 ( 
.A1(n_22),
.A2(n_23),
.B1(n_242),
.B2(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

HB1xp67_ASAP7_75t_SL g175 ( 
.A(n_23),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_23),
.B(n_225),
.C(n_488),
.Y(n_487)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_36),
.B1(n_47),
.B2(n_54),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_24),
.A2(n_47),
.B(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_24),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_24),
.A2(n_36),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_25),
.B(n_56),
.Y(n_55)
);

AO22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_27),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_27),
.Y(n_461)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_37),
.B(n_55),
.Y(n_145)
);

OAI211xp5_ASAP7_75t_SL g335 ( 
.A1(n_38),
.A2(n_336),
.B(n_339),
.C(n_342),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_38),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_38),
.B(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_42),
.Y(n_299)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_46),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_46),
.Y(n_456)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_55),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_58),
.Y(n_304)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_63),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_64),
.Y(n_171)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_113),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_67),
.B(n_175),
.C(n_176),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_92),
.B1(n_104),
.B2(n_110),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_68),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_69),
.A2(n_111),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_69),
.A2(n_111),
.B1(n_226),
.B2(n_227),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g492 ( 
.A1(n_69),
.A2(n_111),
.B(n_226),
.Y(n_492)
);

NAND2x1p5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_83),
.Y(n_69)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

AOI22x1_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B1(n_78),
.B2(n_80),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_77),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_77),
.Y(n_219)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_91),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_90),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_96),
.B(n_97),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_101),
.Y(n_353)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_104),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_109),
.B(n_458),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_111),
.B(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_141),
.C(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_113),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_113),
.A2(n_147),
.B1(n_148),
.B2(n_176),
.Y(n_268)
);

NAND2x1_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_114),
.A2(n_204),
.B1(n_210),
.B2(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_115),
.B(n_355),
.Y(n_354)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_118),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_121),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_122),
.B(n_213),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_135),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_123),
.B(n_212),
.Y(n_211)
);

OAI21xp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_130),
.B(n_135),
.Y(n_123)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_124),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_129),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_129),
.Y(n_263)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_135)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_137),
.Y(n_251)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_138),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_138),
.Y(n_398)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_142),
.B(n_268),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_143),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_143),
.B(n_242),
.C(n_467),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_144),
.B(n_492),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

XOR2x2_ASAP7_75t_L g274 ( 
.A(n_146),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_154),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_155),
.Y(n_346)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_174),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_160),
.B(n_163),
.C(n_174),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_172),
.B(n_173),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_164),
.A2(n_172),
.B1(n_222),
.B2(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_273),
.B(n_278),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_264),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_179),
.B(n_264),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_223),
.C(n_239),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_180),
.A2(n_181),
.B1(n_223),
.B2(n_224),
.Y(n_514)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_220),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_203),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_183),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_183),
.A2(n_184),
.B1(n_271),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_196),
.Y(n_184)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_185),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_186),
.A2(n_246),
.B1(n_252),
.B2(n_253),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_186),
.Y(n_362)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_187),
.B(n_328),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_188),
.B(n_355),
.Y(n_404)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_192),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_192),
.Y(n_333)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_192),
.Y(n_391)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_194),
.Y(n_255)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp33_ASAP7_75t_SL g252 ( 
.A(n_196),
.Y(n_252)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_210),
.B(n_211),
.Y(n_203)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AO22x2_ASAP7_75t_L g256 ( 
.A1(n_210),
.A2(n_213),
.B1(n_234),
.B2(n_257),
.Y(n_256)
);

AO22x2_ASAP7_75t_L g320 ( 
.A1(n_210),
.A2(n_213),
.B1(n_234),
.B2(n_257),
.Y(n_320)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_214),
.Y(n_395)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_219),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_221),
.Y(n_272)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B(n_238),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_232),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_225),
.A2(n_428),
.B1(n_429),
.B2(n_432),
.Y(n_427)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_225),
.Y(n_432)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B(n_237),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_235),
.A2(n_387),
.B1(n_392),
.B2(n_396),
.Y(n_386)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_238),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_239),
.B(n_514),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_240),
.B(n_424),
.C(n_425),
.Y(n_423)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_242),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_242),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_242),
.A2(n_322),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_242),
.Y(n_507)
);

XNOR2x1_ASAP7_75t_L g505 ( 
.A(n_244),
.B(n_506),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_256),
.Y(n_244)
);

XOR2x2_ASAP7_75t_L g494 ( 
.A(n_245),
.B(n_374),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_246),
.A2(n_380),
.B(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_256),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_256),
.B(n_416),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_256),
.A2(n_374),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_256),
.B(n_435),
.C(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_270),
.C(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_271),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_276),
.Y(n_278)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_276),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_282),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_L g530 ( 
.A(n_282),
.B(n_308),
.C(n_531),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_290),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_305),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_312),
.Y(n_531)
);

NAND2x1p5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_522),
.Y(n_312)
);

AOI21x1_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_470),
.B(n_521),
.Y(n_313)
);

AO21x2_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_437),
.B(n_469),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_422),
.B(n_436),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_375),
.B(n_421),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_358),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_318),
.B(n_358),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.Y(n_318)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_320),
.A2(n_321),
.B1(n_385),
.B2(n_386),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_320),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_320),
.A2(n_321),
.B1(n_479),
.B2(n_483),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_320),
.B(n_479),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_321),
.B(n_385),
.Y(n_414)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_323),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_356),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_335),
.C(n_347),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g356 ( 
.A1(n_326),
.A2(n_348),
.B(n_357),
.Y(n_356)
);

OAI21xp33_ASAP7_75t_SL g434 ( 
.A1(n_326),
.A2(n_348),
.B(n_357),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_334),
.Y(n_326)
);

OA22x2_ASAP7_75t_L g417 ( 
.A1(n_327),
.A2(n_362),
.B1(n_363),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_328),
.B(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_335),
.Y(n_357)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_345),
.Y(n_449)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_354),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_373),
.C(n_374),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_401),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_360),
.B(n_401),
.Y(n_411)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_L g442 ( 
.A1(n_361),
.A2(n_443),
.B(n_462),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_361),
.B(n_443),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B(n_368),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_364),
.B(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_372),
.Y(n_383)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_372),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_373),
.B(n_417),
.Y(n_416)
);

AOI21x1_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_413),
.B(n_420),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_399),
.B(n_412),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_384),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_384),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_378),
.A2(n_379),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_378),
.B(n_430),
.C(n_432),
.Y(n_463)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_403),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx2_ASAP7_75t_R g419 ( 
.A(n_383),
.Y(n_419)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_402),
.B(n_411),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_414),
.B(n_415),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_426),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_433),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_427),
.Y(n_439)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_434),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_440),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_464),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_463),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

AO22x1_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_447),
.B1(n_453),
.B2(n_457),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_446),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_450),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx11_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

BUFx12f_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_462),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_463),
.Y(n_500)
);

MAJx2_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_499),
.C(n_500),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_465),
.B(n_492),
.C(n_493),
.Y(n_512)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_467),
.Y(n_468)
);

NOR2x1_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_501),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_495),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_472),
.B(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_486),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_473),
.B(n_486),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_478),
.C(n_484),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_497),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_476),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_485),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_479),
.Y(n_483)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_517),
.C(n_518),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_494),
.Y(n_489)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_490),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_494),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_498),
.Y(n_495)
);

NOR2x1_ASAP7_75t_L g527 ( 
.A(n_496),
.B(n_498),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_515),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_502),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_513),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_503),
.B(n_513),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_508),
.C(n_511),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_505),
.B(n_509),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g511 ( 
.A(n_512),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_515),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_519),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_519),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_524),
.Y(n_522)
);

A2O1A1Ixp33_ASAP7_75t_L g524 ( 
.A1(n_525),
.A2(n_526),
.B(n_528),
.C(n_529),
.Y(n_524)
);


endmodule