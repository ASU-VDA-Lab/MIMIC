module fake_jpeg_30534_n_139 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_139);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_22),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_0),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_57),
.CI(n_49),
.CON(n_77),
.SN(n_77)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_0),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_63),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_71),
.Y(n_79)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_50),
.B1(n_51),
.B2(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_51),
.B1(n_50),
.B2(n_43),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_49),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_7),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_53),
.C(n_52),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_81),
.C(n_90),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_94),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_87),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_93),
.B1(n_1),
.B2(n_2),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_48),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_2),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_46),
.B1(n_42),
.B2(n_21),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_104),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_108),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_4),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_5),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_6),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_111),
.B(n_113),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_7),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

XNOR2x1_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_9),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_111),
.B(n_110),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_10),
.B(n_12),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_13),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_127),
.B(n_128),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_109),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_114),
.B1(n_122),
.B2(n_115),
.Y(n_131)
);

AOI321xp33_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_114),
.A3(n_118),
.B1(n_120),
.B2(n_116),
.C(n_119),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_132),
.B1(n_97),
.B2(n_130),
.Y(n_134)
);

OAI31xp33_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_14),
.A3(n_17),
.B(n_19),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_23),
.B(n_25),
.C(n_26),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_137),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_27),
.Y(n_139)
);


endmodule