module fake_jpeg_4076_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_37),
.Y(n_55)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_23),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_50),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_45),
.B(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_22),
.Y(n_77)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_17),
.B(n_18),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_15),
.C(n_20),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_24),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_25),
.B1(n_17),
.B2(n_21),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_15),
.B1(n_20),
.B2(n_29),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_37),
.B(n_35),
.C(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_64),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_25),
.B1(n_35),
.B2(n_16),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_19),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_76),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_48),
.B1(n_58),
.B2(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_30),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_34),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_82),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_42),
.A2(n_25),
.B1(n_29),
.B2(n_33),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_58),
.B1(n_56),
.B2(n_42),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_52),
.C(n_48),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_92),
.C(n_101),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_67),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_93),
.B1(n_96),
.B2(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_62),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_45),
.C(n_59),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_75),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_68),
.B1(n_44),
.B2(n_65),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_100),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_34),
.B(n_33),
.C(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_44),
.B1(n_20),
.B2(n_15),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_69),
.B1(n_66),
.B2(n_72),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_106),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_74),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_79),
.C(n_76),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_66),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_92),
.C(n_87),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_123),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_90),
.B(n_99),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_138),
.B(n_142),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_136),
.C(n_110),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_99),
.B1(n_102),
.B2(n_93),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_104),
.C(n_86),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_86),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_98),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_98),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_144),
.C(n_150),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_112),
.C(n_106),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_118),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_152),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_121),
.B1(n_123),
.B2(n_122),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_121),
.C(n_109),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_114),
.C(n_27),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_153),
.C(n_129),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_27),
.B1(n_22),
.B2(n_14),
.C(n_13),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_27),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_27),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_157),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_127),
.B1(n_125),
.B2(n_130),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_133),
.B(n_147),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_166),
.B(n_170),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_133),
.B1(n_130),
.B2(n_137),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_161),
.A2(n_163),
.B1(n_22),
.B2(n_2),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_138),
.B1(n_137),
.B2(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_158),
.Y(n_173)
);

XOR2x2_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_138),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_22),
.C(n_12),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_142),
.B(n_22),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_142),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_179),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_173),
.A2(n_178),
.B(n_167),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_176),
.C(n_180),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_11),
.C(n_10),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_162),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_10),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_1),
.C(n_2),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_179),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_184),
.B(n_175),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_167),
.B(n_163),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_186),
.C(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_172),
.B(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_169),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_180),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_190),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_4),
.C(n_5),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_193),
.C(n_181),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_4),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_194),
.A2(n_7),
.B1(n_9),
.B2(n_188),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_185),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_SL g199 ( 
.A(n_197),
.B(n_191),
.C(n_7),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g201 ( 
.A(n_198),
.B(n_9),
.CI(n_195),
.CON(n_201),
.SN(n_201)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_199),
.A2(n_197),
.B(n_200),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_196),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule