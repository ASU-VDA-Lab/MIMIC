module real_jpeg_24073_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_0),
.B(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_0),
.B(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_0),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_0),
.B(n_17),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_0),
.B(n_32),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_0),
.B(n_53),
.Y(n_288)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_2),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_2),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_2),
.B(n_48),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_2),
.B(n_67),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_2),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_5),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_5),
.B(n_32),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_5),
.B(n_53),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_5),
.B(n_36),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_5),
.B(n_50),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_5),
.B(n_48),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_5),
.B(n_67),
.Y(n_289)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_7),
.B(n_53),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_7),
.B(n_50),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_7),
.B(n_32),
.Y(n_183)
);

NAND2x1_ASAP7_75t_SL g198 ( 
.A(n_7),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_7),
.B(n_48),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_7),
.B(n_67),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_7),
.B(n_92),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_8),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_8),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_8),
.B(n_36),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_8),
.B(n_32),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_8),
.B(n_53),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_9),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_9),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_32),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_9),
.B(n_53),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_9),
.B(n_50),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_9),
.B(n_48),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_9),
.B(n_67),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_11),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_11),
.B(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_11),
.B(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_11),
.B(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_11),
.B(n_261),
.Y(n_260)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_11),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_11),
.B(n_53),
.Y(n_323)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_13),
.B(n_48),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_13),
.B(n_67),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_13),
.B(n_50),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_13),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_13),
.B(n_32),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_13),
.B(n_92),
.Y(n_233)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_14),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_14),
.B(n_48),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_16),
.B(n_50),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_16),
.B(n_48),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_16),
.B(n_53),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_16),
.B(n_32),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_16),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_16),
.B(n_67),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_16),
.B(n_92),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_16),
.B(n_128),
.Y(n_303)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_17),
.Y(n_166)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_17),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_139),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_97),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_21),
.B(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.C(n_71),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_22),
.B(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.C(n_46),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_23),
.B(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_29),
.C(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_61),
.Y(n_82)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_29),
.B(n_85),
.C(n_96),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_29),
.A2(n_39),
.B1(n_84),
.B2(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_30),
.B(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_31),
.B(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_34),
.A2(n_38),
.B1(n_41),
.B2(n_316),
.Y(n_315)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_37),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_41),
.C(n_42),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_40),
.B(n_46),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_41),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_42),
.A2(n_43),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_46),
.Y(n_356)
);

FAx1_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.CI(n_52),
.CON(n_46),
.SN(n_46)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_49),
.C(n_52),
.Y(n_101)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_54),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_55),
.B(n_71),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.C(n_70),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_56),
.A2(n_57),
.B1(n_339),
.B2(n_341),
.Y(n_338)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.C(n_63),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_58),
.B(n_60),
.CI(n_63),
.CON(n_310),
.SN(n_310)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_62),
.B(n_64),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_75),
.C(n_77),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_66),
.A2(n_70),
.B1(n_76),
.B2(n_340),
.Y(n_339)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_70),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_73),
.Y(n_75)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_74),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_78),
.A2(n_79),
.B1(n_97),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_88),
.B2(n_89),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_90),
.C(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g125 ( 
.A(n_82),
.B(n_85),
.C(n_86),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_86),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_86),
.A2(n_87),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.C(n_94),
.Y(n_90)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_93),
.CI(n_94),
.CON(n_102),
.SN(n_102)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_97),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_104),
.C(n_107),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.C(n_102),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_99),
.B(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_101),
.B(n_102),
.Y(n_347)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_102),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_111),
.C(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_113),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g357 ( 
.A(n_120),
.Y(n_357)
);

FAx1_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_122),
.CI(n_123),
.CON(n_120),
.SN(n_120)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_127),
.Y(n_134)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_351),
.C(n_352),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_343),
.C(n_344),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_328),
.C(n_329),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_305),
.C(n_306),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_272),
.C(n_273),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_240),
.C(n_241),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_215),
.C(n_216),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_176),
.C(n_187),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_161),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_149),
.B(n_156),
.C(n_161),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_154),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_151),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_159),
.C(n_160),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_169),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_162),
.B(n_170),
.C(n_171),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_163),
.A2(n_164),
.B1(n_167),
.B2(n_168),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_166),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_172),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_173),
.B(n_175),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.C(n_186),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_181),
.B1(n_186),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_191)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_211),
.C(n_212),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_196),
.C(n_202),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_194),
.C(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.C(n_206),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_205),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_210),
.B(n_302),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_229),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_230),
.C(n_239),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_225),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_224),
.C(n_225),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_220),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_223),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_225),
.Y(n_359)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.CI(n_228),
.CON(n_225),
.SN(n_225)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_227),
.C(n_228),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_239),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_237),
.B2(n_238),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_233),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_236),
.C(n_238),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_256),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_245),
.C(n_256),
.Y(n_272)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_247),
.B(n_252),
.C(n_255),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g358 ( 
.A(n_247),
.Y(n_358)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.CI(n_250),
.CON(n_247),
.SN(n_247)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_248),
.B(n_249),
.C(n_250),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_264),
.C(n_270),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_264),
.B1(n_270),
.B2(n_271),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_259),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_262),
.B(n_263),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_262),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_263),
.B(n_296),
.C(n_297),
.Y(n_318)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_292),
.B2(n_304),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_293),
.C(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_278),
.C(n_285),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_285),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_281),
.C(n_284),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_290),
.C(n_291),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_303),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_301),
.C(n_303),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_326),
.B2(n_327),
.Y(n_306)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_317),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_317),
.C(n_326),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g362 ( 
.A(n_310),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_320),
.C(n_321),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_332),
.C(n_342),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_335),
.B2(n_342),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_335),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_335),
.Y(n_355)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.CI(n_338),
.CON(n_335),
.SN(n_335)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_336),
.B(n_337),
.C(n_338),
.Y(n_350)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_348),
.C(n_350),
.Y(n_351)
);


endmodule