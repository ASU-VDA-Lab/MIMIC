module fake_jpeg_18534_n_163 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_163);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_31),
.Y(n_60)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_22),
.Y(n_66)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_18),
.B1(n_15),
.B2(n_23),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_10),
.B1(n_60),
.B2(n_63),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_23),
.B1(n_18),
.B2(n_15),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_53),
.B1(n_56),
.B2(n_65),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_30),
.B(n_21),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_57),
.B(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_51),
.B(n_55),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_30),
.B1(n_20),
.B2(n_21),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_30),
.B(n_20),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_19),
.B1(n_28),
.B2(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_69),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_15),
.B1(n_22),
.B2(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_35),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_25),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_34),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_4),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_24),
.A3(n_19),
.B1(n_22),
.B2(n_12),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_82),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_85),
.B1(n_88),
.B2(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_71),
.B1(n_60),
.B2(n_47),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_4),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_5),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_8),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_91),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_9),
.B1(n_10),
.B2(n_71),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_9),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_89),
.B(n_94),
.Y(n_111)
);

OAI22x1_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_50),
.B1(n_70),
.B2(n_52),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_58),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_10),
.B(n_69),
.C(n_56),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_76),
.B(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_66),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_113),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_62),
.B1(n_73),
.B2(n_50),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_108),
.A2(n_109),
.B(n_110),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_62),
.B(n_70),
.Y(n_109)
);

OA21x2_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_92),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_73),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_92),
.B1(n_64),
.B2(n_47),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_99),
.C(n_101),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_108),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_76),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_122),
.B(n_110),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_93),
.C(n_80),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_120),
.C(n_102),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_85),
.C(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_102),
.Y(n_131)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

AO221x1_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_92),
.B1(n_116),
.B2(n_114),
.C(n_118),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_135),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_134),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_131),
.A2(n_133),
.B(n_127),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_137),
.B(n_115),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_112),
.C(n_77),
.Y(n_133)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_113),
.B1(n_103),
.B2(n_88),
.C(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_97),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_105),
.C(n_104),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_114),
.C(n_120),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_92),
.B(n_96),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_119),
.B1(n_64),
.B2(n_127),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_145),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_136),
.A2(n_121),
.B1(n_125),
.B2(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_146),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_135),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_140),
.C(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_137),
.B1(n_128),
.B2(n_146),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_152),
.A2(n_144),
.B(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_144),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_159),
.B(n_145),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_154),
.A2(n_152),
.B(n_148),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_161),
.B(n_130),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_153),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_129),
.B(n_52),
.Y(n_163)
);


endmodule