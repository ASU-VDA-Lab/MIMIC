module fake_jpeg_26171_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_30)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_4),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_44),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g71 ( 
.A(n_48),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_50),
.B(n_54),
.Y(n_74)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_41),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_56),
.B(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_19),
.B1(n_28),
.B2(n_32),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_29),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_19),
.B1(n_32),
.B2(n_23),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_31),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_63),
.B(n_71),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_35),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_30),
.B1(n_19),
.B2(n_18),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_66),
.B1(n_17),
.B2(n_34),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_37),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

BUFx24_ASAP7_75t_SL g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_89),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_29),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_18),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_35),
.Y(n_78)
);

AO21x2_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_35),
.B(n_29),
.Y(n_79)
);

OR2x6_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_22),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_22),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_26),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_78),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_104),
.Y(n_112)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_60),
.B(n_24),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_31),
.C(n_71),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_46),
.C(n_69),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_51),
.B(n_53),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_105),
.B(n_56),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_67),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_107),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_24),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_108),
.Y(n_111)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_52),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_23),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_20),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_107),
.A2(n_83),
.B1(n_76),
.B2(n_79),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_101),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_76),
.B(n_87),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_120),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_87),
.B1(n_58),
.B2(n_81),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_87),
.B1(n_40),
.B2(n_80),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_99),
.B(n_105),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_122),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_69),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_93),
.Y(n_138)
);

OAI31xp33_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_24),
.A3(n_16),
.B(n_20),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_104),
.C(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_134),
.Y(n_140)
);

XNOR2x1_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_131),
.A2(n_133),
.B1(n_111),
.B2(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_132),
.B(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_97),
.C(n_98),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_135),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_123),
.B(n_118),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_147),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_136),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_4),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_131),
.B1(n_128),
.B2(n_115),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_150),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_127),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_126),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_15),
.B(n_14),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_145),
.A2(n_126),
.B1(n_15),
.B2(n_14),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_5),
.B(n_6),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_157),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_153),
.A2(n_6),
.B(n_8),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_16),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_150),
.C(n_152),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_159),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_161),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_167),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_166),
.B(n_164),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_11),
.B(n_12),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_12),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_168),
.B(n_13),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_24),
.Y(n_172)
);


endmodule