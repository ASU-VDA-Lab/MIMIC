module real_jpeg_16130_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_47;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_48;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI22xp5_ASAP7_75t_L g10 ( 
.A1(n_0),
.A2(n_11),
.B1(n_12),
.B2(n_17),
.Y(n_10)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_15),
.Y(n_32)
);

OR2x4_ASAP7_75t_L g7 ( 
.A(n_1),
.B(n_8),
.Y(n_7)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_10),
.Y(n_9)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_2),
.B(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_3),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_3),
.B(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_5),
.B(n_25),
.Y(n_42)
);

OAI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_9),
.B(n_18),
.C(n_43),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_7),
.B(n_42),
.Y(n_41)
);

AND2x4_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_29),
.Y(n_28)
);

OR2x4_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

NAND3xp33_ASAP7_75t_SL g47 ( 
.A(n_13),
.B(n_34),
.C(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

AOI211xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_24),
.B(n_26),
.C(n_41),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B(n_35),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_27),
.A2(n_37),
.B1(n_45),
.B2(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);


endmodule