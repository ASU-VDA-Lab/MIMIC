module real_aes_4984_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_17;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_20;
wire n_18;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
O2A1O1Ixp33_ASAP7_75t_SL g6 ( .A1(n_0), .A2(n_7), .B(n_16), .C(n_17), .Y(n_6) );
INVx1_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
BUFx2_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
AOI21xp33_ASAP7_75t_SL g16 ( .A1(n_2), .A2(n_3), .B(n_5), .Y(n_16) );
AND3x1_ASAP7_75t_L g21 ( .A(n_2), .B(n_11), .C(n_15), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_3), .B(n_20), .Y(n_19) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_4), .B(n_12), .Y(n_15) );
INVx1_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_5), .A2(n_14), .B(n_15), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g7 ( .A(n_8), .Y(n_7) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_12), .B(n_13), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
BUFx8_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
AND2x4_ASAP7_75t_L g17 ( .A(n_18), .B(n_21), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_19), .Y(n_18) );
endmodule