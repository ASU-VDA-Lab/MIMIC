module fake_jpeg_23424_n_41 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_1),
.C(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_0),
.B(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

AND2x6_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_8),
.B1(n_14),
.B2(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_13),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_13),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_8),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_24),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_33),
.B1(n_26),
.B2(n_25),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_30),
.C(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_19),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_23),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_37),
.B(n_30),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_39),
.B1(n_34),
.B2(n_18),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_22),
.B(n_27),
.Y(n_41)
);


endmodule