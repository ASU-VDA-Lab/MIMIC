module fake_jpeg_16657_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_8),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_31),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_1),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_21),
.B1(n_20),
.B2(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_34),
.B1(n_21),
.B2(n_27),
.Y(n_59)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_72),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_51),
.C(n_44),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_19),
.C(n_50),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_17),
.B1(n_36),
.B2(n_26),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_37),
.B1(n_16),
.B2(n_27),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_78),
.B(n_83),
.Y(n_89)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_42),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_16),
.B1(n_36),
.B2(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_20),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_85),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_37),
.B1(n_26),
.B2(n_23),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_57),
.B1(n_56),
.B2(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_84),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_38),
.B1(n_28),
.B2(n_26),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_29),
.B(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_28),
.B1(n_29),
.B2(n_22),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_19),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_92),
.A2(n_95),
.B(n_106),
.C(n_25),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_19),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_105),
.Y(n_115)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_50),
.C(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_108),
.Y(n_136)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_50),
.Y(n_105)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_29),
.A3(n_19),
.B1(n_32),
.B2(n_28),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_28),
.B(n_32),
.C(n_22),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_95),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_80),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVxp67_ASAP7_75t_SL g111 ( 
.A(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_25),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_60),
.B1(n_83),
.B2(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_112),
.A2(n_123),
.B1(n_97),
.B2(n_107),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_59),
.B1(n_73),
.B2(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_114),
.B(n_131),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_85),
.A3(n_73),
.B1(n_72),
.B2(n_84),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_120),
.Y(n_140)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_132),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_128),
.C(n_130),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_69),
.B1(n_63),
.B2(n_68),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_3),
.B(n_4),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_1),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_127),
.A2(n_129),
.B(n_135),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_32),
.C(n_22),
.Y(n_128)
);

BUFx12f_ASAP7_75t_SL g129 ( 
.A(n_106),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_68),
.C(n_63),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_86),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_90),
.B(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_104),
.Y(n_148)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_113),
.B(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_143),
.B(n_158),
.Y(n_174)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_108),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_138),
.B(n_121),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_92),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_4),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_115),
.B(n_135),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_157),
.B(n_5),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_164),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_88),
.B(n_93),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_154),
.B(n_167),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_138),
.B1(n_5),
.B2(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_88),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_165),
.C(n_117),
.Y(n_172)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_103),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_96),
.B1(n_93),
.B2(n_86),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_185)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_25),
.B(n_2),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_101),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_9),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_134),
.B(n_133),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_4),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_8),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_178),
.C(n_186),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_179),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_156),
.B1(n_169),
.B2(n_148),
.Y(n_200)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_133),
.A3(n_134),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_194),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_182),
.B(n_184),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_149),
.A2(n_5),
.B(n_6),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_187),
.B(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_10),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_144),
.B(n_141),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_11),
.B(n_12),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_154),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_161),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_11),
.C(n_12),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_207),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_202),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_151),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_187),
.B1(n_176),
.B2(n_192),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_172),
.A2(n_168),
.B1(n_160),
.B2(n_150),
.Y(n_204)
);

AO21x2_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_155),
.B(n_167),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_153),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_208),
.A2(n_158),
.B(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_188),
.B(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_164),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_189),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_194),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_175),
.A2(n_154),
.B1(n_161),
.B2(n_167),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_215),
.A2(n_175),
.B1(n_173),
.B2(n_183),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_180),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_195),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_220),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_186),
.C(n_178),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_223),
.C(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_145),
.C(n_165),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_202),
.C(n_215),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_225),
.A2(n_157),
.B(n_185),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_229),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_142),
.B1(n_191),
.B2(n_182),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_230),
.B1(n_206),
.B2(n_196),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_210),
.B1(n_196),
.B2(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_235),
.C(n_239),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_228),
.A2(n_206),
.B1(n_197),
.B2(n_201),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_SL g237 ( 
.A(n_219),
.B(n_213),
.C(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_224),
.A2(n_212),
.B1(n_207),
.B2(n_205),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_220),
.B1(n_223),
.B2(n_216),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_229),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_199),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_159),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_245),
.B(n_247),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_216),
.C(n_217),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_254),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_241),
.B(n_230),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_218),
.B(n_227),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_163),
.C(n_184),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_234),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_256),
.B(n_261),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_253),
.A2(n_243),
.B(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_242),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_146),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_262),
.B(n_246),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_162),
.B1(n_14),
.B2(n_15),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_267),
.B(n_268),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_252),
.B1(n_262),
.B2(n_246),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_252),
.B(n_256),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_272),
.A2(n_266),
.B(n_13),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_273),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_276),
.B(n_274),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_13),
.C(n_14),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_14),
.Y(n_279)
);


endmodule