module fake_jpeg_29230_n_488 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_488);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_488;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_51),
.B(n_61),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx5_ASAP7_75t_SL g111 ( 
.A(n_54),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_17),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_60),
.B(n_69),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_0),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_62),
.Y(n_154)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_17),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_75),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_74),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_78),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_36),
.A2(n_14),
.B1(n_12),
.B2(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_79),
.A2(n_46),
.B1(n_20),
.B2(n_35),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_82),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_42),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_93),
.Y(n_104)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_30),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_37),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_96),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_14),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_99),
.Y(n_131)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_62),
.A2(n_40),
.B1(n_44),
.B2(n_39),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_105),
.A2(n_109),
.B1(n_117),
.B2(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_40),
.B1(n_37),
.B2(n_30),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_106),
.A2(n_119),
.B1(n_136),
.B2(n_143),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_35),
.B1(n_28),
.B2(n_20),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_SL g110 ( 
.A(n_51),
.B(n_46),
.C(n_44),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_50),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_90),
.A2(n_39),
.B1(n_34),
.B2(n_31),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_28),
.B1(n_41),
.B2(n_31),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_39),
.B1(n_47),
.B2(n_34),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_130),
.A2(n_144),
.B1(n_96),
.B2(n_111),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_61),
.B(n_47),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_132),
.B(n_141),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_67),
.A2(n_39),
.B1(n_19),
.B2(n_2),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_106),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_80),
.A2(n_14),
.B1(n_1),
.B2(n_3),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_60),
.B(n_0),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_92),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_152),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_88),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_52),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_92),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_89),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_155),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_157),
.Y(n_234)
);

INVx5_ASAP7_75t_SL g158 ( 
.A(n_115),
.Y(n_158)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_159),
.Y(n_214)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_161),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_169),
.Y(n_216)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_165),
.Y(n_256)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_102),
.B(n_84),
.C(n_98),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_194),
.C(n_154),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_103),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_57),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_171),
.B(n_190),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_176),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_173),
.A2(n_205),
.B1(n_211),
.B2(n_144),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_111),
.A2(n_54),
.B1(n_65),
.B2(n_55),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_113),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_96),
.B(n_64),
.C(n_70),
.Y(n_177)
);

XNOR2x2_ASAP7_75t_SL g237 ( 
.A(n_177),
.B(n_192),
.Y(n_237)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_183),
.Y(n_223)
);

OR2x2_ASAP7_75t_SL g180 ( 
.A(n_139),
.B(n_99),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_180),
.B(n_181),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_85),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_182),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_185),
.Y(n_250)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_108),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_104),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_196),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_56),
.Y(n_190)
);

NOR2x1_ASAP7_75t_R g192 ( 
.A(n_135),
.B(n_63),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_124),
.B(n_156),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_193),
.B(n_197),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_125),
.B(n_68),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_124),
.A2(n_6),
.B(n_8),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_100),
.B(n_94),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_200),
.B(n_203),
.Y(n_257)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_201),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_202),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_208),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_108),
.A2(n_76),
.B1(n_74),
.B2(n_73),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_145),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_128),
.A2(n_53),
.B1(n_76),
.B2(n_59),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_114),
.B1(n_128),
.B2(n_134),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_133),
.B(n_59),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_209),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_154),
.B(n_73),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_210),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_213),
.B(n_235),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_157),
.A2(n_115),
.B(n_130),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_222),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_224),
.A2(n_254),
.B1(n_194),
.B2(n_187),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_168),
.B(n_103),
.C(n_101),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_249),
.C(n_177),
.Y(n_258)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_190),
.A2(n_117),
.A3(n_74),
.B1(n_153),
.B2(n_151),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_199),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_162),
.A2(n_151),
.B(n_114),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_241),
.A2(n_169),
.B1(n_184),
.B2(n_182),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_162),
.A2(n_134),
.B1(n_138),
.B2(n_118),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_247),
.A2(n_255),
.B1(n_187),
.B2(n_209),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_167),
.B(n_180),
.C(n_171),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_192),
.A2(n_145),
.B(n_151),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_252),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_163),
.A2(n_138),
.B1(n_140),
.B2(n_149),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_181),
.A2(n_140),
.B1(n_149),
.B2(n_116),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_258),
.B(n_275),
.Y(n_316)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_228),
.B(n_191),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_261),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_250),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_262),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_234),
.A2(n_158),
.B1(n_165),
.B2(n_202),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_263),
.A2(n_221),
.B(n_242),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_SL g264 ( 
.A(n_237),
.B(n_181),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_264),
.A2(n_252),
.B(n_211),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_225),
.B(n_183),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_265),
.B(n_269),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_266),
.A2(n_292),
.B1(n_248),
.B2(n_243),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_166),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_268),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_239),
.B(n_208),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_227),
.B(n_172),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_159),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_270),
.B(n_274),
.Y(n_337)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_240),
.Y(n_271)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_272),
.Y(n_319)
);

AO21x2_ASAP7_75t_L g273 ( 
.A1(n_230),
.A2(n_222),
.B(n_252),
.Y(n_273)
);

OA22x2_ASAP7_75t_L g322 ( 
.A1(n_273),
.A2(n_253),
.B1(n_256),
.B2(n_236),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_199),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_229),
.B(n_164),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_227),
.B(n_175),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_276),
.B(n_280),
.Y(n_309)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_214),
.Y(n_277)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_278),
.A2(n_255),
.B1(n_241),
.B2(n_247),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_218),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_279),
.B(n_284),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_250),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_281),
.A2(n_285),
.B1(n_298),
.B2(n_242),
.Y(n_315)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_283),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_223),
.B(n_195),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_235),
.A2(n_185),
.B1(n_204),
.B2(n_198),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_232),
.B(n_160),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_288),
.B(n_290),
.Y(n_335)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_245),
.B(n_161),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_250),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_295),
.Y(n_336)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_294),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_245),
.B(n_179),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_232),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_296),
.Y(n_304)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g334 ( 
.A(n_297),
.B(n_299),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_215),
.B(n_170),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_215),
.B(n_201),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_249),
.C(n_213),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_300),
.B(n_301),
.C(n_307),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_246),
.C(n_216),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_303),
.A2(n_308),
.B1(n_315),
.B2(n_333),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_306),
.A2(n_310),
.B(n_273),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_258),
.B(n_246),
.C(n_216),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_274),
.A2(n_237),
.B1(n_221),
.B2(n_254),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_286),
.A2(n_216),
.B(n_246),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_317),
.B(n_220),
.Y(n_367)
);

AOI22x1_ASAP7_75t_SL g321 ( 
.A1(n_273),
.A2(n_226),
.B1(n_248),
.B2(n_243),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_321),
.A2(n_336),
.B(n_328),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_322),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_194),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_328),
.C(n_288),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_325),
.A2(n_260),
.B1(n_262),
.B2(n_280),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_231),
.C(n_212),
.Y(n_328)
);

BUFx10_ASAP7_75t_L g332 ( 
.A(n_272),
.Y(n_332)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_332),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_281),
.A2(n_178),
.B1(n_212),
.B2(n_226),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_269),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_338),
.B(n_350),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_341),
.A2(n_322),
.B(n_306),
.Y(n_370)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_319),
.Y(n_343)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_316),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_345),
.B(n_352),
.Y(n_393)
);

NOR2x1_ASAP7_75t_R g346 ( 
.A(n_321),
.B(n_264),
.Y(n_346)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_346),
.B(n_349),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_347),
.A2(n_348),
.B1(n_354),
.B2(n_359),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_326),
.A2(n_260),
.B1(n_267),
.B2(n_270),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_296),
.Y(n_350)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_316),
.B(n_268),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_325),
.A2(n_273),
.B1(n_291),
.B2(n_276),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_273),
.C(n_265),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_358),
.C(n_361),
.Y(n_376)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_356),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_330),
.B(n_261),
.C(n_259),
.Y(n_357)
);

NAND3xp33_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_311),
.C(n_327),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_294),
.C(n_293),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_317),
.A2(n_292),
.B1(n_283),
.B2(n_282),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_277),
.Y(n_360)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_360),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_297),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_302),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_362),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_289),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_363),
.B(n_368),
.Y(n_369)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_313),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_364),
.Y(n_374)
);

XNOR2x1_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_253),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_367),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_244),
.C(n_220),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_310),
.C(n_304),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_309),
.B(n_244),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_370),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_346),
.A2(n_322),
.B(n_335),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_372),
.A2(n_387),
.B(n_233),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_313),
.Y(n_373)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_373),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_368),
.B(n_363),
.Y(n_375)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_375),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_383),
.C(n_391),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_382),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_322),
.C(n_308),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_339),
.A2(n_319),
.B1(n_320),
.B2(n_329),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_386),
.A2(n_339),
.B1(n_342),
.B2(n_314),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_341),
.A2(n_334),
.B(n_333),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_343),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_389),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_353),
.A2(n_329),
.B1(n_318),
.B2(n_303),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_340),
.B(n_318),
.C(n_314),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_355),
.B(n_320),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_394),
.B(n_349),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_359),
.Y(n_395)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_395),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_351),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_406),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_399),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_340),
.C(n_366),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_408),
.C(n_416),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_354),
.Y(n_404)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_404),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_344),
.Y(n_405)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_405),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_352),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_385),
.A2(n_353),
.B1(n_383),
.B2(n_380),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_407),
.A2(n_409),
.B1(n_389),
.B2(n_388),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_358),
.C(n_361),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_378),
.B(n_365),
.Y(n_410)
);

XNOR2x1_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_411),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_378),
.B(n_367),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_415),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_332),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_377),
.C(n_381),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_384),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_417),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_332),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_387),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_371),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_423),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_404),
.A2(n_385),
.B1(n_392),
.B2(n_375),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_411),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_427),
.A2(n_414),
.B1(n_403),
.B2(n_369),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_407),
.A2(n_401),
.B1(n_396),
.B2(n_397),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_428),
.A2(n_433),
.B1(n_410),
.B2(n_256),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_405),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_431),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_371),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_372),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_415),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_374),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_408),
.C(n_416),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_436),
.C(n_398),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_369),
.C(n_370),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_439),
.Y(n_461)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_426),
.Y(n_440)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_440),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_434),
.A2(n_414),
.B(n_403),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_441),
.A2(n_420),
.B(n_432),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g442 ( 
.A1(n_424),
.A2(n_390),
.B1(n_379),
.B2(n_412),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_442),
.A2(n_449),
.B1(n_437),
.B2(n_10),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_443),
.B(n_446),
.Y(n_453)
);

XNOR2x1_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_421),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_436),
.A2(n_379),
.B(n_390),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_447),
.B(n_420),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_332),
.C(n_217),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_448),
.B(n_429),
.C(n_435),
.Y(n_457)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_233),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_424),
.A2(n_189),
.B1(n_186),
.B2(n_11),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_450),
.B(n_451),
.Y(n_455)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_425),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_457),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_459),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_421),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_460),
.A2(n_439),
.B(n_443),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_9),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_463),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_452),
.A2(n_437),
.B1(n_10),
.B2(n_11),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_464),
.B(n_450),
.C(n_438),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_454),
.A2(n_452),
.B(n_441),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_466),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_460),
.A2(n_451),
.B(n_440),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_453),
.B(n_448),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_471),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_469),
.B(n_473),
.Y(n_476)
);

NOR2x1_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_444),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_470),
.A2(n_457),
.B(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_475),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_472),
.B(n_455),
.Y(n_477)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_477),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_468),
.B(n_461),
.C(n_459),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_478),
.A2(n_473),
.B(n_461),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_480),
.B(n_476),
.Y(n_484)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_482),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_483),
.A2(n_484),
.B1(n_474),
.B2(n_481),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_479),
.C(n_472),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_486),
.B(n_9),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_487),
.B(n_9),
.Y(n_488)
);


endmodule