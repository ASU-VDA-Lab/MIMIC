module fake_netlist_6_2504_n_1717 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1717);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1717;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_40),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_84),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_87),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_41),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_6),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_48),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_88),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_57),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_48),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_51),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_128),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_42),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_51),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_97),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_103),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_55),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_2),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_28),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_65),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_70),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_29),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_89),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_67),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_15),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_43),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_45),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_109),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_96),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_0),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_59),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_91),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_105),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_123),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_38),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_7),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_23),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_72),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_47),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_61),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_113),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_21),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_81),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_56),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_7),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_131),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_28),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_124),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_5),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_39),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_90),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_22),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_56),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_92),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_69),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_117),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_17),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_62),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_22),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_60),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_66),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_54),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_49),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_99),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_148),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_144),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_58),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_130),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_46),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_14),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_114),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_2),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_0),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_59),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_94),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_37),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_102),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_135),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_119),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_53),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_140),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_26),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_55),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_30),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_82),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_54),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_58),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_19),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_57),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_79),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_40),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_156),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_46),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_98),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_14),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_146),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_17),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_73),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_43),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_74),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_100),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_93),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_42),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_12),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_95),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_6),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_125),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_3),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_5),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_60),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_23),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_118),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_13),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_10),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_39),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_129),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_52),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_21),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_127),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_47),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_27),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_33),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_8),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_108),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_80),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_104),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_120),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_115),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_52),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_76),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_153),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_112),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_45),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_25),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_38),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_71),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_75),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_160),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_267),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_205),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_158),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_267),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_267),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_161),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_170),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_203),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_164),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_267),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_169),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_205),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_203),
.B(n_1),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_1),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_209),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_188),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_267),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

BUFx2_ASAP7_75t_SL g334 ( 
.A(n_197),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_179),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_175),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_258),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_176),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_179),
.Y(n_339)
);

BUFx2_ASAP7_75t_SL g340 ( 
.A(n_197),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_212),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_282),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_253),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_199),
.B(n_3),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_212),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_212),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_177),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_183),
.Y(n_348)
);

AND2x6_ASAP7_75t_L g349 ( 
.A(n_163),
.B(n_151),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_187),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_212),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_212),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_190),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_273),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_201),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_273),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_209),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_251),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_199),
.B(n_4),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_202),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_273),
.Y(n_362)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_167),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_208),
.Y(n_364)
);

INVxp33_ASAP7_75t_SL g365 ( 
.A(n_157),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_211),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_273),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_213),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_216),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_287),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_159),
.B(n_4),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_265),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_251),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_218),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_219),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_282),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_226),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_227),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_287),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_230),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_287),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_162),
.B(n_171),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_228),
.B(n_8),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_233),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_165),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_287),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_167),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_340),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_385),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_330),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_335),
.B(n_287),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_312),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_346),
.B(n_162),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_351),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_313),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_351),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_352),
.B(n_354),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_352),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_355),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_355),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_357),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_325),
.A2(n_280),
.B1(n_166),
.B2(n_174),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_339),
.B(n_278),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_373),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_349),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_359),
.B(n_311),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_367),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_367),
.B(n_171),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_370),
.B(n_182),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_313),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_373),
.B(n_278),
.Y(n_429)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_316),
.B(n_163),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_316),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_370),
.B(n_236),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_317),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_379),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_317),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_321),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_349),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_321),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_349),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_182),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_386),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_386),
.B(n_283),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_323),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_328),
.B(n_168),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_334),
.B(n_237),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_323),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_325),
.A2(n_285),
.B1(n_220),
.B2(n_178),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_332),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_332),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_333),
.B(n_274),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_340),
.B(n_238),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_349),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_333),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_391),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_401),
.B(n_429),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_446),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_395),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_401),
.B(n_429),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_429),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_390),
.B(n_318),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_391),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_390),
.B(n_319),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_401),
.B(n_336),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

AO22x2_ASAP7_75t_L g468 ( 
.A1(n_447),
.A2(n_320),
.B1(n_360),
.B2(n_185),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_446),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_447),
.B(n_365),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_395),
.Y(n_472)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_403),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_399),
.B(n_338),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_451),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_423),
.B(n_348),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

INVx6_ASAP7_75t_L g480 ( 
.A(n_405),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_405),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_410),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_410),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

BUFx4f_ASAP7_75t_L g486 ( 
.A(n_405),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_419),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_350),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_419),
.B(n_382),
.C(n_371),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_399),
.B(n_353),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

CKINVDCx6p67_ASAP7_75t_R g492 ( 
.A(n_448),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_420),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_454),
.B(n_356),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_419),
.B(n_372),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_454),
.B(n_361),
.Y(n_497)
);

BUFx4f_ASAP7_75t_L g498 ( 
.A(n_405),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_420),
.B(n_364),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_391),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_L g501 ( 
.A1(n_396),
.A2(n_342),
.B1(n_327),
.B2(n_329),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_422),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_451),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_422),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_422),
.B(n_274),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_423),
.B(n_366),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_432),
.B(n_369),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_452),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_400),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_396),
.B(n_374),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_452),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_400),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_456),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_422),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_432),
.B(n_377),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_422),
.B(n_360),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_398),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_456),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_445),
.B(n_378),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_398),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_398),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_453),
.A2(n_382),
.B(n_181),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_415),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_398),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_391),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_407),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_445),
.Y(n_531)
);

BUFx10_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

AO21x2_ASAP7_75t_L g533 ( 
.A1(n_453),
.A2(n_181),
.B(n_159),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_438),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_453),
.A2(n_314),
.B1(n_358),
.B2(n_344),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_428),
.B(n_384),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_445),
.B(n_347),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_438),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_428),
.B(n_268),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_438),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_398),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_417),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_453),
.A2(n_358),
.B1(n_344),
.B2(n_383),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_428),
.B(n_368),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_422),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_428),
.B(n_240),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_450),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

AO22x1_ASAP7_75t_L g549 ( 
.A1(n_453),
.A2(n_242),
.B1(n_246),
.B2(n_262),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_422),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_428),
.B(n_243),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_425),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_391),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_436),
.B(n_249),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_450),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_440),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_409),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_440),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_440),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_394),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_449),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_404),
.A2(n_383),
.B1(n_269),
.B2(n_228),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_455),
.B(n_343),
.Y(n_563)
);

BUFx6f_ASAP7_75t_SL g564 ( 
.A(n_425),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_415),
.B(n_342),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_404),
.A2(n_269),
.B1(n_294),
.B2(n_296),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_L g568 ( 
.A1(n_425),
.A2(n_241),
.B1(n_173),
.B2(n_214),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_415),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_404),
.B(n_194),
.C(n_191),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_436),
.B(n_375),
.Y(n_571)
);

AND2x2_ASAP7_75t_SL g572 ( 
.A(n_425),
.B(n_163),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_455),
.B(n_380),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_409),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_394),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_436),
.B(n_266),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_394),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_415),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_449),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_449),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_436),
.B(n_363),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_404),
.B(n_387),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_394),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_425),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_388),
.B(n_387),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_394),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_394),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_436),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_404),
.A2(n_427),
.B1(n_426),
.B2(n_443),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_426),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_431),
.B(n_434),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_426),
.A2(n_294),
.B1(n_296),
.B2(n_283),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_426),
.B(n_191),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_431),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_426),
.A2(n_246),
.B1(n_308),
.B2(n_291),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_431),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_394),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_394),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_427),
.B(n_194),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_402),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_431),
.B(n_270),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_388),
.B(n_315),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_425),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_434),
.B(n_409),
.Y(n_604)
);

INVxp33_ASAP7_75t_L g605 ( 
.A(n_427),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_427),
.B(n_198),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_474),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_487),
.B(n_466),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_572),
.B(n_475),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_L g610 ( 
.A(n_471),
.B(n_489),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_462),
.B(n_180),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_572),
.B(n_425),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_566),
.B(n_184),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_508),
.A2(n_322),
.B1(n_324),
.B2(n_331),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_491),
.B(n_425),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_468),
.A2(n_349),
.B1(n_427),
.B2(n_443),
.Y(n_616)
);

BUFx5_ASAP7_75t_L g617 ( 
.A(n_481),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_526),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_459),
.Y(n_619)
);

BUFx6f_ASAP7_75t_SL g620 ( 
.A(n_467),
.Y(n_620)
);

NOR3xp33_ASAP7_75t_L g621 ( 
.A(n_501),
.B(n_189),
.C(n_186),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_581),
.B(n_434),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_475),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_517),
.B(n_434),
.Y(n_624)
);

AO22x2_ASAP7_75t_L g625 ( 
.A1(n_547),
.A2(n_198),
.B1(n_250),
.B2(n_310),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_557),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_458),
.B(n_402),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_458),
.B(n_402),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_531),
.B(n_337),
.Y(n_629)
);

O2A1O1Ixp5_ASAP7_75t_L g630 ( 
.A1(n_605),
.A2(n_443),
.B(n_409),
.C(n_229),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_569),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_475),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_569),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_461),
.B(n_488),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_459),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_565),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_468),
.A2(n_306),
.B1(n_272),
.B2(n_305),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_468),
.A2(n_443),
.B1(n_455),
.B2(n_442),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_495),
.B(n_402),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_478),
.B(n_402),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_566),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_470),
.B(n_402),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_475),
.Y(n_643)
);

NOR2x1p5_ASAP7_75t_L g644 ( 
.A(n_492),
.B(n_192),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_470),
.B(n_402),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_572),
.B(n_437),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_483),
.B(n_193),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_477),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_475),
.B(n_437),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_475),
.B(n_479),
.Y(n_651)
);

BUFx5_ASAP7_75t_L g652 ( 
.A(n_481),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_467),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_585),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_565),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_574),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_504),
.B(n_510),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_504),
.B(n_443),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_510),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_513),
.B(n_389),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_574),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_SL g662 ( 
.A1(n_542),
.A2(n_264),
.B1(n_168),
.B2(n_265),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_479),
.B(n_437),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_513),
.B(n_389),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_515),
.B(n_392),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_590),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_515),
.B(n_392),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_489),
.A2(n_250),
.B1(n_310),
.B2(n_206),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_483),
.B(n_196),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_468),
.A2(n_518),
.B1(n_492),
.B2(n_509),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_590),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_520),
.B(n_522),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_520),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_537),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_526),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_473),
.A2(n_235),
.B(n_239),
.C(n_232),
.Y(n_676)
);

NOR2x1_ASAP7_75t_L g677 ( 
.A(n_573),
.B(n_206),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_479),
.B(n_437),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_511),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_496),
.B(n_265),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_518),
.A2(n_222),
.B1(n_229),
.B2(n_281),
.Y(n_681)
);

BUFx6f_ASAP7_75t_SL g682 ( 
.A(n_467),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_518),
.A2(n_455),
.B1(n_442),
.B2(n_439),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_496),
.B(n_265),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_511),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_536),
.B(n_393),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_526),
.Y(n_687)
);

BUFx8_ASAP7_75t_L g688 ( 
.A(n_542),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_588),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_486),
.A2(n_455),
.B(n_437),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_518),
.A2(n_533),
.B1(n_599),
.B2(n_593),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_479),
.B(n_437),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_539),
.B(n_393),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_588),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_502),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_578),
.B(n_397),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_578),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_593),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_479),
.B(n_437),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_479),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_544),
.A2(n_571),
.B1(n_563),
.B2(n_497),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_511),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_463),
.B(n_200),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_582),
.B(n_397),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_582),
.B(n_406),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_514),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_601),
.B(n_406),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_494),
.B(n_437),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_482),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_465),
.B(n_204),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_589),
.B(n_500),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_518),
.A2(n_455),
.B1(n_442),
.B2(n_439),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_494),
.B(n_439),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_599),
.B(n_408),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_585),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_494),
.B(n_439),
.Y(n_716)
);

O2A1O1Ixp5_ASAP7_75t_L g717 ( 
.A1(n_486),
.A2(n_210),
.B(n_281),
.C(n_290),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_555),
.B(n_207),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_606),
.B(n_604),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_494),
.B(n_439),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_494),
.B(n_439),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_502),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_494),
.B(n_439),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_502),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_546),
.B(n_408),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_584),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_602),
.B(n_411),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_551),
.B(n_411),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_R g729 ( 
.A(n_493),
.B(n_275),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_521),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_535),
.B(n_215),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_554),
.B(n_412),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_576),
.B(n_412),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_512),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_548),
.B(n_413),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_584),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_603),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_514),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_514),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_SL g740 ( 
.A1(n_543),
.A2(n_277),
.B1(n_252),
.B2(n_245),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_499),
.A2(n_301),
.B1(n_302),
.B2(n_299),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_476),
.B(n_217),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_584),
.B(n_439),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_490),
.B(n_223),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_SL g745 ( 
.A(n_568),
.B(n_168),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_460),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_562),
.B(n_224),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_549),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_548),
.B(n_553),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_584),
.B(n_442),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_460),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_L g752 ( 
.A1(n_570),
.A2(n_247),
.B1(n_286),
.B2(n_290),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_529),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_584),
.B(n_603),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_530),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_584),
.B(n_442),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_603),
.B(n_442),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_548),
.B(n_413),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_469),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_533),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_530),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_603),
.B(n_442),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_592),
.B(n_231),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_595),
.B(n_234),
.C(n_309),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_603),
.B(n_442),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_549),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_553),
.B(n_414),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_603),
.B(n_244),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_570),
.B(n_414),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_534),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_553),
.B(n_560),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_486),
.B(n_455),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_498),
.B(n_455),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_498),
.A2(n_444),
.B(n_441),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_560),
.B(n_416),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_634),
.B(n_491),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_617),
.B(n_498),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_608),
.B(n_491),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_610),
.A2(n_567),
.B(n_289),
.C(n_172),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_626),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_608),
.B(n_491),
.Y(n_781)
);

BUFx2_ASAP7_75t_SL g782 ( 
.A(n_620),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_612),
.A2(n_552),
.B(n_591),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_615),
.A2(n_552),
.B(n_505),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_760),
.A2(n_533),
.B1(n_480),
.B2(n_564),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_615),
.A2(n_552),
.B(n_505),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_672),
.B(n_505),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_754),
.A2(n_505),
.B(n_503),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_623),
.A2(n_516),
.B(n_503),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_636),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_631),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_612),
.A2(n_525),
.B(n_594),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_655),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_736),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_701),
.A2(n_670),
.B1(n_677),
.B2(n_698),
.Y(n_795)
);

AND2x6_ASAP7_75t_L g796 ( 
.A(n_748),
.B(n_736),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_703),
.A2(n_291),
.B(n_289),
.C(n_288),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_654),
.B(n_525),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_674),
.B(n_480),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_623),
.A2(n_516),
.B(n_503),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_629),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_624),
.B(n_457),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_715),
.B(n_480),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_647),
.B(n_222),
.C(n_210),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_673),
.B(n_457),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_618),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_632),
.A2(n_726),
.B(n_643),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_656),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_611),
.B(n_255),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_R g810 ( 
.A(n_607),
.B(n_276),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_686),
.B(n_457),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_657),
.B(n_464),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_617),
.B(n_481),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_L g814 ( 
.A(n_617),
.B(n_506),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_661),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_653),
.B(n_560),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_711),
.B(n_464),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_614),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_646),
.A2(n_594),
.B(n_596),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_617),
.B(n_481),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_690),
.A2(n_771),
.B(n_749),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_663),
.A2(n_600),
.B(n_577),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_619),
.B(n_464),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_619),
.B(n_464),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_635),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_703),
.A2(n_710),
.B1(n_666),
.B2(n_671),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_709),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_710),
.A2(n_254),
.B(n_288),
.C(n_172),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_618),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_646),
.A2(n_596),
.B(n_534),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_734),
.B(n_480),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_617),
.B(n_652),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_632),
.A2(n_503),
.B(n_516),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_635),
.B(n_484),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_668),
.A2(n_538),
.B(n_580),
.C(n_579),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_609),
.A2(n_558),
.B(n_538),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_648),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_643),
.A2(n_516),
.B(n_503),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_653),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_637),
.A2(n_247),
.B(n_225),
.C(n_286),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_641),
.B(n_484),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_648),
.B(n_484),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_727),
.A2(n_564),
.B1(n_506),
.B2(n_597),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_676),
.A2(n_540),
.B(n_579),
.C(n_556),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_726),
.A2(n_628),
.B(n_627),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_639),
.A2(n_545),
.B(n_550),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_718),
.B(n_631),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_736),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_649),
.B(n_484),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_633),
.B(n_485),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_609),
.A2(n_540),
.B(n_556),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_737),
.A2(n_550),
.B(n_545),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_649),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_659),
.B(n_485),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_633),
.B(n_485),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_652),
.B(n_532),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_737),
.A2(n_550),
.B(n_545),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_691),
.A2(n_564),
.B1(n_506),
.B2(n_597),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_659),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_611),
.B(n_257),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_644),
.B(n_485),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_704),
.B(n_528),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_676),
.A2(n_256),
.B(n_185),
.C(n_195),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_736),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_683),
.A2(n_550),
.B(n_545),
.Y(n_865)
);

OAI21xp33_ASAP7_75t_L g866 ( 
.A1(n_647),
.A2(n_260),
.B(n_261),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_712),
.A2(n_640),
.B(n_719),
.Y(n_867)
);

OR2x2_ASAP7_75t_SL g868 ( 
.A(n_744),
.B(n_195),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_679),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_638),
.A2(n_564),
.B1(n_577),
.B2(n_587),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_768),
.A2(n_506),
.B1(n_598),
.B2(n_597),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_705),
.B(n_528),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_613),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_652),
.B(n_532),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_697),
.B(n_528),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_768),
.A2(n_506),
.B1(n_598),
.B2(n_597),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_772),
.A2(n_545),
.B(n_532),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_622),
.B(n_693),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_773),
.A2(n_532),
.B(n_600),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_689),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_773),
.A2(n_600),
.B(n_577),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_685),
.Y(n_882)
);

AO21x1_ASAP7_75t_L g883 ( 
.A1(n_681),
.A2(n_225),
.B(n_580),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_669),
.B(n_263),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_630),
.A2(n_558),
.B(n_559),
.Y(n_885)
);

NOR2x2_ASAP7_75t_L g886 ( 
.A(n_745),
.B(n_662),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_651),
.A2(n_587),
.B(n_586),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_707),
.B(n_598),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_725),
.B(n_598),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_731),
.A2(n_235),
.B(n_221),
.C(n_232),
.Y(n_890)
);

O2A1O1Ixp5_ASAP7_75t_L g891 ( 
.A1(n_717),
.A2(n_587),
.B(n_586),
.C(n_583),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_652),
.B(n_586),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_728),
.B(n_528),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_732),
.B(n_583),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_685),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_663),
.A2(n_561),
.B(n_559),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_752),
.A2(n_561),
.B(n_472),
.C(n_469),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_733),
.B(n_575),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_722),
.A2(n_506),
.B1(n_575),
.B2(n_583),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_SL g900 ( 
.A(n_620),
.B(n_264),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_651),
.A2(n_583),
.B(n_575),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_694),
.Y(n_902)
);

AOI21xp33_ASAP7_75t_L g903 ( 
.A1(n_747),
.A2(n_297),
.B(n_295),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_650),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_724),
.A2(n_575),
.B1(n_541),
.B2(n_527),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_678),
.A2(n_472),
.B(n_507),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_766),
.B(n_523),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_730),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_680),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_678),
.A2(n_541),
.B(n_527),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_675),
.B(n_507),
.Y(n_911)
);

AOI21xp33_ASAP7_75t_L g912 ( 
.A1(n_742),
.A2(n_271),
.B(n_292),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_702),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_702),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_687),
.A2(n_714),
.B1(n_616),
.B2(n_695),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_692),
.A2(n_721),
.B(n_723),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_684),
.B(n_523),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_692),
.A2(n_524),
.B(n_519),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_699),
.A2(n_716),
.B(n_743),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_699),
.A2(n_713),
.B(n_743),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_669),
.B(n_524),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_700),
.B(n_519),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_660),
.B(n_519),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_708),
.A2(n_506),
.B(n_430),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_664),
.B(n_416),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_708),
.A2(n_444),
.B(n_441),
.Y(n_926)
);

NAND2x1p5_ASAP7_75t_L g927 ( 
.A(n_700),
.B(n_163),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_706),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_713),
.A2(n_433),
.B(n_418),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_706),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_740),
.B(n_284),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_665),
.B(n_418),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_738),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_SL g934 ( 
.A(n_621),
.B(n_303),
.C(n_307),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_667),
.B(n_433),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_696),
.B(n_435),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_625),
.B(n_256),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_716),
.A2(n_421),
.B(n_424),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_720),
.A2(n_421),
.B(n_424),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_763),
.B(n_279),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_720),
.A2(n_435),
.B(n_163),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_729),
.B(n_264),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_753),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_721),
.A2(n_300),
.B(n_298),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_723),
.A2(n_430),
.B(n_293),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_769),
.B(n_221),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_750),
.A2(n_756),
.B(n_757),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_755),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_658),
.B(n_300),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_761),
.A2(n_304),
.B1(n_430),
.B2(n_300),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_750),
.A2(n_300),
.B(n_308),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_770),
.A2(n_430),
.B1(n_300),
.B2(n_262),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_738),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_756),
.A2(n_430),
.B(n_254),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_757),
.A2(n_248),
.B(n_242),
.C(n_239),
.Y(n_955)
);

AOI22x1_ASAP7_75t_L g956 ( 
.A1(n_746),
.A2(n_248),
.B1(n_430),
.B2(n_147),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_791),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_940),
.B(n_741),
.C(n_764),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_878),
.B(n_746),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_825),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_791),
.Y(n_961)
);

OAI21xp33_ASAP7_75t_L g962 ( 
.A1(n_903),
.A2(n_912),
.B(n_884),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_784),
.A2(n_765),
.B(n_762),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_786),
.A2(n_820),
.B(n_813),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_827),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_837),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_794),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_826),
.B(n_729),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_847),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_794),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_813),
.A2(n_765),
.B(n_762),
.Y(n_971)
);

OA22x2_ASAP7_75t_L g972 ( 
.A1(n_937),
.A2(n_625),
.B1(n_688),
.B2(n_682),
.Y(n_972)
);

CKINVDCx16_ASAP7_75t_R g973 ( 
.A(n_810),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_853),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_909),
.B(n_688),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_940),
.A2(n_804),
.B(n_795),
.C(n_921),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_794),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_778),
.B(n_759),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_859),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_804),
.A2(n_921),
.B(n_909),
.C(n_867),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_847),
.B(n_625),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_840),
.A2(n_642),
.B(n_645),
.C(n_767),
.Y(n_982)
);

AOI21x1_ASAP7_75t_L g983 ( 
.A1(n_892),
.A2(n_775),
.B(n_758),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_SL g984 ( 
.A1(n_797),
.A2(n_735),
.B(n_739),
.C(n_751),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_801),
.B(n_682),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_820),
.A2(n_650),
.B(n_774),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_873),
.B(n_688),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_908),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_781),
.B(n_759),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_797),
.A2(n_751),
.B(n_739),
.C(n_11),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_L g991 ( 
.A(n_796),
.B(n_650),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_856),
.A2(n_650),
.B(n_430),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_SL g993 ( 
.A1(n_799),
.A2(n_831),
.B(n_855),
.C(n_850),
.Y(n_993)
);

OAI21xp33_ASAP7_75t_SL g994 ( 
.A1(n_907),
.A2(n_650),
.B(n_10),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_856),
.A2(n_430),
.B(n_145),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_809),
.B(n_860),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_848),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_848),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_SL g999 ( 
.A(n_904),
.B(n_430),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_SL g1000 ( 
.A1(n_907),
.A2(n_9),
.B(n_11),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_942),
.B(n_9),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_810),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_785),
.A2(n_787),
.B1(n_890),
.B2(n_937),
.Y(n_1003)
);

O2A1O1Ixp5_ASAP7_75t_L g1004 ( 
.A1(n_949),
.A2(n_141),
.B(n_138),
.C(n_137),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_828),
.A2(n_12),
.B(n_13),
.C(n_16),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_799),
.B(n_430),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_874),
.A2(n_134),
.B(n_126),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_869),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_782),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_892),
.A2(n_122),
.B(n_121),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_882),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_874),
.A2(n_111),
.B(n_107),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_866),
.B(n_16),
.Y(n_1013)
);

OAI22x1_ASAP7_75t_SL g1014 ( 
.A1(n_818),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_1014)
);

NOR2x1_ASAP7_75t_L g1015 ( 
.A(n_839),
.B(n_106),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_776),
.B(n_101),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_816),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_946),
.B(n_18),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_890),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_828),
.A2(n_26),
.B(n_29),
.C(n_30),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_831),
.B(n_811),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_937),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_946),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_798),
.Y(n_1024)
);

AOI33xp33_ASAP7_75t_L g1025 ( 
.A1(n_943),
.A2(n_31),
.A3(n_32),
.B1(n_33),
.B2(n_34),
.B3(n_35),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_948),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_931),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_880),
.B(n_35),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_925),
.B(n_86),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_858),
.A2(n_36),
.B1(n_37),
.B2(n_41),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_794),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_902),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_931),
.A2(n_78),
.B1(n_77),
.B2(n_68),
.Y(n_1033)
);

OAI22x1_ASAP7_75t_L g1034 ( 
.A1(n_886),
.A2(n_36),
.B1(n_44),
.B2(n_49),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_777),
.A2(n_63),
.B(n_50),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_895),
.Y(n_1036)
);

AO32x2_ASAP7_75t_L g1037 ( 
.A1(n_915),
.A2(n_44),
.A3(n_50),
.B1(n_53),
.B2(n_870),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_816),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_913),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_949),
.A2(n_817),
.B(n_845),
.Y(n_1040)
);

NOR2xp67_ASAP7_75t_L g1041 ( 
.A(n_934),
.B(n_793),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_914),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_832),
.A2(n_814),
.B(n_865),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_868),
.A2(n_904),
.B1(n_780),
.B2(n_815),
.Y(n_1044)
);

OR2x4_ASAP7_75t_L g1045 ( 
.A(n_850),
.B(n_855),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_900),
.B(n_841),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_932),
.B(n_935),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_802),
.A2(n_888),
.B(n_889),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_822),
.A2(n_821),
.B(n_881),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_917),
.A2(n_790),
.B(n_920),
.C(n_916),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_893),
.A2(n_894),
.B(n_812),
.Y(n_1051)
);

O2A1O1Ixp5_ASAP7_75t_L g1052 ( 
.A1(n_883),
.A2(n_898),
.B(n_783),
.C(n_891),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_808),
.B(n_936),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_861),
.B(n_841),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_877),
.A2(n_872),
.B(n_862),
.Y(n_1055)
);

OAI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_779),
.A2(n_829),
.B1(n_806),
.B2(n_863),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_863),
.A2(n_779),
.B(n_898),
.C(n_955),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_803),
.B(n_806),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_803),
.B(n_796),
.Y(n_1059)
);

INVx5_ASAP7_75t_L g1060 ( 
.A(n_796),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_947),
.A2(n_844),
.B(n_835),
.C(n_851),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_788),
.A2(n_807),
.B(n_923),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_SL g1063 ( 
.A1(n_792),
.A2(n_885),
.B(n_836),
.C(n_843),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_928),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_796),
.B(n_829),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_930),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_796),
.Y(n_1067)
);

AO21x2_ASAP7_75t_L g1068 ( 
.A1(n_830),
.A2(n_819),
.B(n_896),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_899),
.A2(n_953),
.B1(n_933),
.B2(n_805),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_864),
.B(n_824),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_911),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_823),
.B(n_834),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_951),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_875),
.B(n_876),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_842),
.B(n_854),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_922),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_927),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_945),
.A2(n_910),
.B(n_918),
.C(n_897),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_879),
.A2(n_846),
.B(n_789),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_922),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_927),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_926),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_849),
.Y(n_1083)
);

INVx5_ASAP7_75t_L g1084 ( 
.A(n_956),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_919),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_871),
.A2(n_887),
.B(n_944),
.C(n_901),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_924),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_906),
.Y(n_1088)
);

AO21x2_ASAP7_75t_L g1089 ( 
.A1(n_905),
.A2(n_939),
.B(n_938),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_800),
.A2(n_833),
.B(n_838),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_929),
.B(n_954),
.Y(n_1091)
);

INVx4_ASAP7_75t_L g1092 ( 
.A(n_852),
.Y(n_1092)
);

INVx4_ASAP7_75t_L g1093 ( 
.A(n_857),
.Y(n_1093)
);

NAND2xp33_ASAP7_75t_SL g1094 ( 
.A(n_950),
.B(n_952),
.Y(n_1094)
);

INVx5_ASAP7_75t_L g1095 ( 
.A(n_941),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_784),
.A2(n_498),
.B(n_486),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_784),
.A2(n_498),
.B(n_486),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_794),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_L g1099 ( 
.A1(n_892),
.A2(n_949),
.B(n_867),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_878),
.A2(n_610),
.B1(n_760),
.B2(n_785),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_848),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_988),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1051),
.A2(n_1048),
.B(n_1047),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1026),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_1052),
.A2(n_1049),
.B(n_1061),
.Y(n_1105)
);

AO21x1_ASAP7_75t_L g1106 ( 
.A1(n_1003),
.A2(n_1030),
.B(n_1013),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_SL g1107 ( 
.A(n_1060),
.B(n_973),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1023),
.B(n_961),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_976),
.A2(n_1086),
.A3(n_1078),
.B(n_1003),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_SL g1110 ( 
.A1(n_1030),
.A2(n_1019),
.B(n_968),
.C(n_1100),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_965),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_980),
.A2(n_958),
.B(n_996),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_969),
.B(n_962),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1050),
.A2(n_1082),
.A3(n_1055),
.B(n_1056),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1017),
.B(n_1038),
.Y(n_1115)
);

INVx6_ASAP7_75t_L g1116 ( 
.A(n_967),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1062),
.A2(n_1097),
.B(n_1096),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1032),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1100),
.A2(n_1001),
.B1(n_981),
.B2(n_1046),
.Y(n_1119)
);

NAND2xp33_ASAP7_75t_L g1120 ( 
.A(n_1060),
.B(n_1067),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1053),
.B(n_1071),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_1067),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_964),
.A2(n_1043),
.B(n_963),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1041),
.A2(n_1057),
.B(n_1029),
.C(n_1094),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1018),
.B(n_1022),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_1027),
.B(n_1000),
.C(n_1044),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_1063),
.A2(n_993),
.B(n_1029),
.C(n_1065),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1044),
.A2(n_1019),
.B1(n_972),
.B2(n_975),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_957),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_986),
.A2(n_1040),
.B(n_1099),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1028),
.A2(n_1005),
.B(n_1020),
.C(n_994),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_990),
.A2(n_987),
.B(n_1021),
.C(n_985),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1021),
.A2(n_1035),
.B(n_1059),
.C(n_1074),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1002),
.B(n_1060),
.Y(n_1134)
);

AOI211x1_ASAP7_75t_L g1135 ( 
.A1(n_959),
.A2(n_960),
.B(n_966),
.C(n_974),
.Y(n_1135)
);

CKINVDCx8_ASAP7_75t_R g1136 ( 
.A(n_1009),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_979),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_1069),
.A2(n_1088),
.A3(n_1016),
.B(n_1092),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1045),
.A2(n_1087),
.B1(n_1060),
.B2(n_1024),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_972),
.A2(n_1034),
.B1(n_1054),
.B2(n_1033),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1016),
.A2(n_971),
.B(n_982),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_967),
.Y(n_1142)
);

NOR2xp67_ASAP7_75t_L g1143 ( 
.A(n_1017),
.B(n_1038),
.Y(n_1143)
);

NOR2x1_ASAP7_75t_L g1144 ( 
.A(n_997),
.B(n_1101),
.Y(n_1144)
);

AOI221x1_ASAP7_75t_L g1145 ( 
.A1(n_1007),
.A2(n_1012),
.B1(n_1058),
.B2(n_978),
.C(n_989),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_983),
.A2(n_992),
.B(n_1075),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1008),
.Y(n_1147)
);

INVx6_ASAP7_75t_L g1148 ( 
.A(n_967),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_991),
.A2(n_959),
.B(n_1091),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1011),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1036),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1072),
.A2(n_1075),
.B(n_1068),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_1025),
.B(n_1015),
.C(n_1083),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1068),
.A2(n_1087),
.B(n_1073),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_L g1155 ( 
.A(n_1004),
.B(n_984),
.C(n_1087),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1087),
.A2(n_995),
.B(n_1006),
.C(n_1064),
.Y(n_1156)
);

INVx3_ASAP7_75t_L g1157 ( 
.A(n_1076),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1039),
.B(n_1066),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1042),
.B(n_1070),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1077),
.B(n_1037),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_997),
.A2(n_1101),
.B1(n_998),
.B2(n_1076),
.Y(n_1161)
);

AO221x2_ASAP7_75t_L g1162 ( 
.A1(n_1014),
.A2(n_1037),
.B1(n_1070),
.B2(n_1084),
.C(n_1010),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1095),
.A2(n_1089),
.B(n_999),
.Y(n_1163)
);

AO32x2_ASAP7_75t_L g1164 ( 
.A1(n_1037),
.A2(n_1092),
.A3(n_1093),
.B1(n_1085),
.B2(n_1084),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_970),
.B(n_977),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1095),
.A2(n_1089),
.B(n_999),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1076),
.B(n_1080),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1080),
.B(n_1085),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_970),
.B(n_977),
.Y(n_1169)
);

NOR4xp25_ASAP7_75t_L g1170 ( 
.A(n_1084),
.B(n_1093),
.C(n_1085),
.D(n_1095),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_970),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1095),
.A2(n_1080),
.B(n_1081),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_977),
.A2(n_1031),
.B(n_1098),
.Y(n_1173)
);

AOI221x1_ASAP7_75t_L g1174 ( 
.A1(n_1031),
.A2(n_1098),
.B1(n_976),
.B2(n_1030),
.C(n_804),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_976),
.A2(n_1047),
.B1(n_610),
.B2(n_701),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1051),
.A2(n_498),
.B(n_486),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1051),
.A2(n_498),
.B(n_486),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_976),
.A2(n_1047),
.B1(n_610),
.B2(n_701),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1051),
.A2(n_498),
.B(n_486),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_962),
.A2(n_976),
.B(n_610),
.C(n_471),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1047),
.B(n_608),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1047),
.B(n_608),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1013),
.A2(n_1100),
.B1(n_610),
.B2(n_962),
.Y(n_1183)
);

AOI221x1_ASAP7_75t_L g1184 ( 
.A1(n_976),
.A2(n_1030),
.B1(n_804),
.B2(n_962),
.C(n_1003),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1051),
.A2(n_498),
.B(n_486),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_988),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_976),
.A2(n_1061),
.A3(n_670),
.B(n_1086),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_976),
.A2(n_1061),
.A3(n_670),
.B(n_1086),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_SL g1189 ( 
.A(n_973),
.B(n_607),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1023),
.B(n_839),
.Y(n_1190)
);

BUFx10_ASAP7_75t_L g1191 ( 
.A(n_985),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_962),
.A2(n_976),
.B(n_610),
.C(n_471),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1067),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1051),
.A2(n_498),
.B(n_486),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_969),
.B(n_674),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1030),
.A2(n_1100),
.B1(n_1003),
.B2(n_670),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_976),
.A2(n_1061),
.A3(n_670),
.B(n_1086),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1051),
.A2(n_498),
.B(n_486),
.Y(n_1198)
);

AO32x2_ASAP7_75t_L g1199 ( 
.A1(n_1100),
.A2(n_1003),
.A3(n_1030),
.B1(n_670),
.B2(n_1019),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_976),
.A2(n_674),
.B(n_471),
.C(n_962),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_976),
.A2(n_1047),
.B1(n_610),
.B2(n_701),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_SL g1202 ( 
.A1(n_990),
.A2(n_1057),
.B(n_1035),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_976),
.A2(n_980),
.B(n_610),
.Y(n_1203)
);

OAI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_1001),
.A2(n_473),
.B(n_471),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_976),
.A2(n_980),
.B(n_610),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_1060),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_1009),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_976),
.A2(n_980),
.B(n_610),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1047),
.B(n_608),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_988),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_976),
.A2(n_674),
.B(n_471),
.C(n_962),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_996),
.B(n_674),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_996),
.B(n_674),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1047),
.B(n_608),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1047),
.B(n_608),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1052),
.A2(n_1049),
.B(n_1061),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1052),
.A2(n_1049),
.B(n_1061),
.Y(n_1217)
);

O2A1O1Ixp5_ASAP7_75t_SL g1218 ( 
.A1(n_1030),
.A2(n_447),
.B(n_1019),
.C(n_670),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1051),
.A2(n_498),
.B(n_486),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1023),
.B(n_839),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_988),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1051),
.A2(n_498),
.B(n_486),
.Y(n_1222)
);

AOI221x1_ASAP7_75t_L g1223 ( 
.A1(n_976),
.A2(n_1030),
.B1(n_804),
.B2(n_962),
.C(n_1003),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_969),
.B(n_674),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1049),
.A2(n_1090),
.B(n_1079),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1013),
.A2(n_1100),
.B1(n_610),
.B2(n_962),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1047),
.B(n_608),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1049),
.A2(n_1090),
.B(n_1079),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_988),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_988),
.Y(n_1230)
);

NOR4xp25_ASAP7_75t_L g1231 ( 
.A(n_1027),
.B(n_976),
.C(n_962),
.D(n_1030),
.Y(n_1231)
);

NOR2xp67_ASAP7_75t_L g1232 ( 
.A(n_958),
.B(n_826),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_SL g1233 ( 
.A(n_1136),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_1142),
.Y(n_1234)
);

INVx2_ASAP7_75t_SL g1235 ( 
.A(n_1129),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1204),
.A2(n_1106),
.B1(n_1162),
.B2(n_1119),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1204),
.A2(n_1162),
.B1(n_1119),
.B2(n_1232),
.Y(n_1237)
);

BUFx12f_ASAP7_75t_L g1238 ( 
.A(n_1207),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1181),
.A2(n_1214),
.B1(n_1227),
.B2(n_1182),
.Y(n_1239)
);

CKINVDCx12_ASAP7_75t_R g1240 ( 
.A(n_1125),
.Y(n_1240)
);

INVx6_ASAP7_75t_L g1241 ( 
.A(n_1190),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1232),
.A2(n_1196),
.B1(n_1208),
.B2(n_1203),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1209),
.A2(n_1215),
.B1(n_1140),
.B2(n_1224),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1140),
.A2(n_1195),
.B1(n_1226),
.B2(n_1183),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1190),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1113),
.A2(n_1212),
.B1(n_1213),
.B2(n_1226),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1184),
.A2(n_1223),
.B1(n_1128),
.B2(n_1183),
.Y(n_1247)
);

CKINVDCx11_ASAP7_75t_R g1248 ( 
.A(n_1111),
.Y(n_1248)
);

OAI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1128),
.A2(n_1121),
.B1(n_1205),
.B2(n_1126),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1104),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1191),
.Y(n_1251)
);

INVx6_ASAP7_75t_L g1252 ( 
.A(n_1220),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1230),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1126),
.A2(n_1153),
.B1(n_1178),
.B2(n_1175),
.Y(n_1254)
);

INVx8_ASAP7_75t_L g1255 ( 
.A(n_1220),
.Y(n_1255)
);

BUFx12f_ASAP7_75t_L g1256 ( 
.A(n_1191),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1196),
.A2(n_1201),
.B1(n_1112),
.B2(n_1153),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1206),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_SL g1259 ( 
.A1(n_1189),
.A2(n_1202),
.B1(n_1164),
.B2(n_1160),
.Y(n_1259)
);

INVx5_ASAP7_75t_L g1260 ( 
.A(n_1206),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1116),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1118),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1108),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1108),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1169),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1200),
.A2(n_1211),
.B(n_1192),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1147),
.B(n_1150),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1115),
.B(n_1151),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1141),
.A2(n_1137),
.B1(n_1229),
.B2(n_1221),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1186),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1180),
.A2(n_1139),
.B1(n_1231),
.B2(n_1115),
.Y(n_1271)
);

BUFx4_ASAP7_75t_SL g1272 ( 
.A(n_1210),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1124),
.A2(n_1132),
.B1(n_1143),
.B2(n_1155),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_1116),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1110),
.A2(n_1159),
.B1(n_1103),
.B2(n_1155),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1174),
.A2(n_1158),
.B1(n_1143),
.B2(n_1163),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1166),
.A2(n_1135),
.B1(n_1131),
.B2(n_1134),
.Y(n_1277)
);

INVx6_ASAP7_75t_L g1278 ( 
.A(n_1148),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1148),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1157),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1144),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1171),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1167),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1165),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1107),
.A2(n_1120),
.B1(n_1161),
.B2(n_1193),
.Y(n_1285)
);

OAI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1199),
.A2(n_1164),
.B1(n_1149),
.B2(n_1152),
.Y(n_1286)
);

NAND2x1p5_ASAP7_75t_L g1287 ( 
.A(n_1144),
.B(n_1172),
.Y(n_1287)
);

BUFx8_ASAP7_75t_L g1288 ( 
.A(n_1199),
.Y(n_1288)
);

BUFx2_ASAP7_75t_SL g1289 ( 
.A(n_1122),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1156),
.A2(n_1122),
.B1(n_1168),
.B2(n_1133),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_SL g1291 ( 
.A1(n_1164),
.A2(n_1199),
.B1(n_1218),
.B2(n_1105),
.Y(n_1291)
);

BUFx8_ASAP7_75t_SL g1292 ( 
.A(n_1127),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1173),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_SL g1294 ( 
.A1(n_1170),
.A2(n_1105),
.B1(n_1216),
.B2(n_1217),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1109),
.B(n_1197),
.Y(n_1295)
);

OR2x2_ASAP7_75t_L g1296 ( 
.A(n_1187),
.B(n_1188),
.Y(n_1296)
);

BUFx4f_ASAP7_75t_SL g1297 ( 
.A(n_1170),
.Y(n_1297)
);

INVx6_ASAP7_75t_L g1298 ( 
.A(n_1154),
.Y(n_1298)
);

BUFx4f_ASAP7_75t_SL g1299 ( 
.A(n_1187),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1216),
.A2(n_1217),
.B1(n_1109),
.B2(n_1188),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1146),
.Y(n_1301)
);

CKINVDCx11_ASAP7_75t_R g1302 ( 
.A(n_1145),
.Y(n_1302)
);

CKINVDCx6p67_ASAP7_75t_R g1303 ( 
.A(n_1197),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1176),
.A2(n_1185),
.B1(n_1194),
.B2(n_1198),
.Y(n_1304)
);

INVx4_ASAP7_75t_L g1305 ( 
.A(n_1123),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1138),
.A2(n_1114),
.B1(n_1117),
.B2(n_1130),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1177),
.A2(n_1222),
.B1(n_1219),
.B2(n_1179),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1114),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1114),
.Y(n_1309)
);

CKINVDCx11_ASAP7_75t_R g1310 ( 
.A(n_1225),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1228),
.B(n_1181),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1204),
.A2(n_1106),
.B1(n_804),
.B2(n_962),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_1195),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1111),
.Y(n_1314)
);

INVx8_ASAP7_75t_L g1315 ( 
.A(n_1142),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1181),
.A2(n_1209),
.B1(n_1214),
.B2(n_1182),
.Y(n_1316)
);

INVx4_ASAP7_75t_SL g1317 ( 
.A(n_1116),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_SL g1318 ( 
.A1(n_1162),
.A2(n_417),
.B1(n_450),
.B2(n_745),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1207),
.Y(n_1319)
);

CKINVDCx11_ASAP7_75t_R g1320 ( 
.A(n_1136),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1181),
.A2(n_1209),
.B1(n_1214),
.B2(n_1182),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1204),
.A2(n_1106),
.B1(n_804),
.B2(n_962),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1125),
.B(n_981),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1109),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1107),
.B(n_1060),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1102),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1142),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1204),
.A2(n_1106),
.B1(n_804),
.B2(n_962),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1162),
.A2(n_417),
.B1(n_450),
.B2(n_745),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1204),
.A2(n_1106),
.B1(n_804),
.B2(n_962),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1181),
.A2(n_1182),
.B1(n_1214),
.B2(n_1209),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1204),
.A2(n_1106),
.B1(n_1013),
.B2(n_962),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1204),
.A2(n_818),
.B1(n_315),
.B2(n_324),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1204),
.A2(n_1106),
.B1(n_804),
.B2(n_962),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1125),
.B(n_981),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1204),
.A2(n_1106),
.B1(n_804),
.B2(n_962),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1181),
.B(n_1182),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1115),
.B(n_1108),
.Y(n_1338)
);

INVx6_ASAP7_75t_L g1339 ( 
.A(n_1142),
.Y(n_1339)
);

INVx6_ASAP7_75t_L g1340 ( 
.A(n_1142),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_1111),
.Y(n_1341)
);

BUFx4f_ASAP7_75t_SL g1342 ( 
.A(n_1111),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1265),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1304),
.A2(n_1247),
.B(n_1254),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1324),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1296),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1297),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1295),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1293),
.Y(n_1349)
);

CKINVDCx6p67_ASAP7_75t_R g1350 ( 
.A(n_1320),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1331),
.B(n_1239),
.Y(n_1351)
);

AOI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1273),
.A2(n_1311),
.B(n_1290),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1308),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1309),
.Y(n_1354)
);

BUFx10_ASAP7_75t_L g1355 ( 
.A(n_1339),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1331),
.B(n_1316),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1297),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1310),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1301),
.Y(n_1359)
);

AOI211x1_ASAP7_75t_L g1360 ( 
.A1(n_1244),
.A2(n_1249),
.B(n_1243),
.C(n_1247),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1318),
.A2(n_1329),
.B1(n_1237),
.B2(n_1302),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1303),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1277),
.A2(n_1305),
.A3(n_1291),
.B(n_1286),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1251),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1307),
.A2(n_1275),
.B(n_1266),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1283),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1294),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1281),
.A2(n_1262),
.B(n_1270),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1284),
.Y(n_1369)
);

INVx5_ASAP7_75t_L g1370 ( 
.A(n_1298),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1259),
.B(n_1242),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1307),
.A2(n_1287),
.B(n_1275),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1299),
.Y(n_1373)
);

AO21x1_ASAP7_75t_L g1374 ( 
.A1(n_1254),
.A2(n_1249),
.B(n_1286),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1306),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1321),
.B(n_1337),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1313),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1256),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1242),
.B(n_1236),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1291),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1288),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1318),
.A2(n_1329),
.B1(n_1237),
.B2(n_1236),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1323),
.B(n_1335),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1288),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1287),
.A2(n_1269),
.B(n_1257),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1300),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1300),
.Y(n_1387)
);

OAI221xp5_ASAP7_75t_L g1388 ( 
.A1(n_1332),
.A2(n_1336),
.B1(n_1328),
.B2(n_1322),
.C(n_1334),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1250),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1246),
.A2(n_1312),
.B1(n_1328),
.B2(n_1330),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1269),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1312),
.A2(n_1336),
.B1(n_1322),
.B2(n_1330),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1253),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1326),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1257),
.B(n_1334),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1268),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1271),
.B(n_1267),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1276),
.A2(n_1325),
.B(n_1260),
.Y(n_1398)
);

BUFx4f_ASAP7_75t_SL g1399 ( 
.A(n_1314),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1292),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1276),
.A2(n_1285),
.B(n_1258),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1263),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1333),
.A2(n_1313),
.B1(n_1264),
.B2(n_1342),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1282),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1289),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1338),
.A2(n_1274),
.B(n_1235),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1338),
.B(n_1245),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1280),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1240),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1245),
.B(n_1317),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1241),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1341),
.B(n_1252),
.Y(n_1412)
);

INVx5_ASAP7_75t_L g1413 ( 
.A(n_1370),
.Y(n_1413)
);

AOI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1360),
.A2(n_1234),
.B1(n_1327),
.B2(n_1315),
.C(n_1255),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1372),
.A2(n_1272),
.B(n_1317),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1388),
.A2(n_1351),
.B(n_1356),
.C(n_1376),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1361),
.A2(n_1342),
.B1(n_1241),
.B2(n_1248),
.Y(n_1417)
);

AOI211xp5_ASAP7_75t_L g1418 ( 
.A1(n_1374),
.A2(n_1279),
.B(n_1261),
.C(n_1272),
.Y(n_1418)
);

NOR2x1_ASAP7_75t_SL g1419 ( 
.A(n_1358),
.B(n_1238),
.Y(n_1419)
);

NAND4xp25_ASAP7_75t_L g1420 ( 
.A(n_1382),
.B(n_1360),
.C(n_1390),
.D(n_1392),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1399),
.B(n_1233),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1343),
.B(n_1315),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1397),
.B(n_1315),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1390),
.A2(n_1340),
.B1(n_1339),
.B2(n_1319),
.Y(n_1424)
);

AOI221xp5_ASAP7_75t_L g1425 ( 
.A1(n_1374),
.A2(n_1234),
.B1(n_1327),
.B2(n_1261),
.C(n_1279),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1368),
.Y(n_1426)
);

OR2x6_ASAP7_75t_L g1427 ( 
.A(n_1398),
.B(n_1339),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1393),
.B(n_1340),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1395),
.B(n_1340),
.Y(n_1429)
);

NOR2x1_ASAP7_75t_SL g1430 ( 
.A(n_1358),
.B(n_1233),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1392),
.A2(n_1278),
.B(n_1401),
.C(n_1395),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1386),
.B(n_1278),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1412),
.B(n_1377),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1383),
.B(n_1369),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1396),
.B(n_1366),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1409),
.B(n_1407),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1386),
.B(n_1387),
.Y(n_1437)
);

O2A1O1Ixp33_ASAP7_75t_SL g1438 ( 
.A1(n_1367),
.A2(n_1381),
.B(n_1384),
.C(n_1362),
.Y(n_1438)
);

OR2x6_ASAP7_75t_L g1439 ( 
.A(n_1385),
.B(n_1373),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1409),
.B(n_1407),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1371),
.A2(n_1379),
.B(n_1385),
.C(n_1375),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1353),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1350),
.B(n_1403),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1406),
.B(n_1402),
.Y(n_1444)
);

OAI21xp33_ASAP7_75t_L g1445 ( 
.A1(n_1371),
.A2(n_1379),
.B(n_1391),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1406),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1375),
.A2(n_1367),
.B(n_1357),
.C(n_1347),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1389),
.B(n_1394),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1389),
.B(n_1394),
.Y(n_1449)
);

NAND2xp33_ASAP7_75t_L g1450 ( 
.A(n_1358),
.B(n_1370),
.Y(n_1450)
);

OAI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1349),
.A2(n_1358),
.B1(n_1357),
.B2(n_1347),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1349),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1346),
.B(n_1363),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1350),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1411),
.B(n_1404),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_L g1456 ( 
.A(n_1358),
.B(n_1370),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1349),
.Y(n_1457)
);

NAND2xp33_ASAP7_75t_L g1458 ( 
.A(n_1358),
.B(n_1370),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1406),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1404),
.B(n_1400),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1453),
.B(n_1363),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1437),
.B(n_1380),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1442),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1453),
.B(n_1363),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1437),
.B(n_1380),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1459),
.B(n_1363),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1439),
.B(n_1363),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1426),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1418),
.A2(n_1375),
.B1(n_1365),
.B2(n_1400),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1439),
.B(n_1363),
.Y(n_1470)
);

NOR2x1_ASAP7_75t_L g1471 ( 
.A(n_1450),
.B(n_1344),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1439),
.B(n_1359),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1446),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1439),
.B(n_1354),
.Y(n_1474)
);

INVxp33_ASAP7_75t_L g1475 ( 
.A(n_1433),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1427),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1444),
.B(n_1345),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1448),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1441),
.B(n_1353),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1449),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1413),
.A2(n_1344),
.B(n_1370),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1416),
.B(n_1408),
.Y(n_1482)
);

BUFx2_ASAP7_75t_R g1483 ( 
.A(n_1454),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1441),
.B(n_1348),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1420),
.A2(n_1344),
.B1(n_1365),
.B2(n_1391),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1485),
.A2(n_1365),
.B1(n_1445),
.B2(n_1417),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1466),
.B(n_1434),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1478),
.B(n_1365),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1467),
.B(n_1415),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1473),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1473),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1467),
.B(n_1415),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1485),
.A2(n_1431),
.B1(n_1447),
.B2(n_1424),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1468),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1482),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1469),
.A2(n_1431),
.B1(n_1443),
.B2(n_1451),
.C(n_1447),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1481),
.B(n_1427),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1469),
.A2(n_1429),
.B1(n_1425),
.B2(n_1457),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1466),
.B(n_1435),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1467),
.B(n_1415),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1475),
.A2(n_1423),
.B1(n_1436),
.B2(n_1440),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1482),
.B(n_1414),
.C(n_1455),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1470),
.B(n_1461),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1466),
.B(n_1348),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1470),
.B(n_1372),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1472),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1461),
.B(n_1464),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1475),
.A2(n_1452),
.B1(n_1427),
.B2(n_1432),
.Y(n_1508)
);

OAI211xp5_ASAP7_75t_L g1509 ( 
.A1(n_1471),
.A2(n_1352),
.B(n_1438),
.C(n_1460),
.Y(n_1509)
);

INVxp67_ASAP7_75t_R g1510 ( 
.A(n_1479),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1463),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1511),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1495),
.B(n_1499),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1494),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1504),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1510),
.B(n_1464),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1510),
.B(n_1503),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1511),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1494),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1495),
.B(n_1422),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1488),
.B(n_1473),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1499),
.B(n_1478),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1488),
.B(n_1477),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1499),
.B(n_1478),
.Y(n_1524)
);

NOR2xp67_ASAP7_75t_L g1525 ( 
.A(n_1509),
.B(n_1481),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1487),
.B(n_1480),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1490),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1504),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1487),
.B(n_1480),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1510),
.B(n_1464),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1503),
.B(n_1479),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1503),
.B(n_1479),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1503),
.B(n_1474),
.Y(n_1533)
);

NAND2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1490),
.B(n_1471),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1494),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1490),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1504),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1506),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1487),
.B(n_1480),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_L g1540 ( 
.A(n_1509),
.B(n_1471),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1494),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1489),
.B(n_1474),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1527),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1515),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1513),
.B(n_1507),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1520),
.B(n_1501),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1515),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1520),
.B(n_1513),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1525),
.B(n_1501),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1525),
.B(n_1502),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1540),
.B(n_1502),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1540),
.B(n_1498),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1528),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1528),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1537),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1527),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1527),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1526),
.B(n_1498),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_L g1560 ( 
.A(n_1526),
.B(n_1454),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1523),
.B(n_1507),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1517),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1523),
.B(n_1507),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1537),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1523),
.B(n_1522),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1522),
.B(n_1484),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1541),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1541),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1512),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1529),
.B(n_1462),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1512),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1512),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1529),
.B(n_1462),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1517),
.B(n_1496),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1518),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1518),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1518),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1517),
.B(n_1489),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1539),
.B(n_1465),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1514),
.Y(n_1580)
);

INVxp67_ASAP7_75t_L g1581 ( 
.A(n_1524),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1514),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1536),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1516),
.B(n_1492),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1514),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1531),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1562),
.B(n_1516),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1552),
.B(n_1531),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1567),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1568),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1547),
.B(n_1531),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1569),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1546),
.B(n_1521),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1550),
.B(n_1532),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1583),
.B(n_1516),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1583),
.B(n_1530),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1544),
.B(n_1530),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1560),
.B(n_1483),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1557),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1546),
.B(n_1521),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1566),
.B(n_1521),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1571),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1578),
.B(n_1530),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1574),
.B(n_1532),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1553),
.B(n_1536),
.Y(n_1605)
);

AND2x2_ASAP7_75t_SL g1606 ( 
.A(n_1559),
.B(n_1496),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1574),
.B(n_1532),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1549),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1566),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1548),
.B(n_1565),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1570),
.B(n_1483),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1581),
.B(n_1533),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1572),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1575),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1576),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1579),
.B(n_1364),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1565),
.B(n_1545),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1577),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1545),
.Y(n_1620)
);

OAI31xp33_ASAP7_75t_L g1621 ( 
.A1(n_1604),
.A2(n_1493),
.A3(n_1534),
.B(n_1486),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1606),
.A2(n_1493),
.B1(n_1497),
.B2(n_1486),
.Y(n_1622)
);

AOI222xp33_ASAP7_75t_L g1623 ( 
.A1(n_1606),
.A2(n_1484),
.B1(n_1421),
.B2(n_1419),
.C1(n_1430),
.C2(n_1564),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1605),
.A2(n_1497),
.B1(n_1427),
.B2(n_1578),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1592),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1607),
.A2(n_1534),
.B(n_1544),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1592),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1595),
.B(n_1558),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1620),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1595),
.B(n_1584),
.Y(n_1630)
);

INVxp67_ASAP7_75t_SL g1631 ( 
.A(n_1599),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1611),
.A2(n_1563),
.B1(n_1561),
.B2(n_1508),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1620),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1602),
.Y(n_1634)
);

OAI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1608),
.A2(n_1497),
.B1(n_1534),
.B2(n_1561),
.Y(n_1635)
);

NOR2x1_ASAP7_75t_L g1636 ( 
.A(n_1618),
.B(n_1558),
.Y(n_1636)
);

OAI22xp33_ASAP7_75t_SL g1637 ( 
.A1(n_1586),
.A2(n_1534),
.B1(n_1563),
.B2(n_1556),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1617),
.A2(n_1497),
.B1(n_1505),
.B2(n_1476),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1613),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1594),
.A2(n_1591),
.B(n_1588),
.Y(n_1640)
);

AOI31xp33_ASAP7_75t_L g1641 ( 
.A1(n_1598),
.A2(n_1609),
.A3(n_1596),
.B(n_1610),
.Y(n_1641)
);

OAI221xp5_ASAP7_75t_L g1642 ( 
.A1(n_1610),
.A2(n_1556),
.B1(n_1554),
.B2(n_1555),
.C(n_1508),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1596),
.B(n_1584),
.Y(n_1643)
);

OAI211xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1618),
.A2(n_1585),
.B(n_1582),
.C(n_1580),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1587),
.A2(n_1505),
.B(n_1492),
.C(n_1500),
.Y(n_1645)
);

NOR4xp25_ASAP7_75t_SL g1646 ( 
.A(n_1631),
.B(n_1589),
.C(n_1590),
.D(n_1615),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1640),
.B(n_1612),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1641),
.B(n_1587),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1641),
.A2(n_1619),
.B(n_1614),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1636),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1629),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1633),
.Y(n_1652)
);

OAI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1622),
.A2(n_1497),
.B1(n_1601),
.B2(n_1593),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1625),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1627),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1634),
.B(n_1601),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1630),
.B(n_1603),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1628),
.B(n_1603),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1639),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1632),
.B(n_1593),
.Y(n_1660)
);

O2A1O1Ixp5_ASAP7_75t_L g1661 ( 
.A1(n_1626),
.A2(n_1597),
.B(n_1600),
.C(n_1555),
.Y(n_1661)
);

AOI33xp33_ASAP7_75t_L g1662 ( 
.A1(n_1635),
.A2(n_1597),
.A3(n_1554),
.B1(n_1505),
.B2(n_1492),
.B3(n_1500),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1628),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1643),
.B(n_1597),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1623),
.B(n_1621),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1656),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1656),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1657),
.B(n_1623),
.Y(n_1668)
);

AOI222xp33_ASAP7_75t_L g1669 ( 
.A1(n_1665),
.A2(n_1642),
.B1(n_1644),
.B2(n_1645),
.C1(n_1616),
.C2(n_1637),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1663),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1648),
.B(n_1600),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1649),
.A2(n_1624),
.B1(n_1638),
.B2(n_1438),
.C(n_1505),
.Y(n_1672)
);

O2A1O1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1650),
.A2(n_1378),
.B(n_1364),
.C(n_1497),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1651),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1660),
.B(n_1524),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1646),
.A2(n_1378),
.B(n_1364),
.Y(n_1676)
);

NOR2x1_ASAP7_75t_L g1677 ( 
.A(n_1666),
.B(n_1654),
.Y(n_1677)
);

NOR3xp33_ASAP7_75t_L g1678 ( 
.A(n_1671),
.B(n_1659),
.C(n_1647),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1667),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1668),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1670),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1675),
.Y(n_1682)
);

AOI222xp33_ASAP7_75t_L g1683 ( 
.A1(n_1672),
.A2(n_1653),
.B1(n_1655),
.B2(n_1652),
.C1(n_1658),
.C2(n_1657),
.Y(n_1683)
);

OAI21xp33_ASAP7_75t_L g1684 ( 
.A1(n_1669),
.A2(n_1664),
.B(n_1662),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_L g1685 ( 
.A(n_1676),
.B(n_1674),
.C(n_1673),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1682),
.Y(n_1686)
);

OAI21xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1677),
.A2(n_1669),
.B(n_1662),
.Y(n_1687)
);

NAND2xp33_ASAP7_75t_R g1688 ( 
.A(n_1679),
.B(n_1661),
.Y(n_1688)
);

O2A1O1Ixp33_ASAP7_75t_L g1689 ( 
.A1(n_1684),
.A2(n_1653),
.B(n_1378),
.C(n_1497),
.Y(n_1689)
);

NOR2x1_ASAP7_75t_L g1690 ( 
.A(n_1680),
.B(n_1538),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1687),
.B(n_1678),
.Y(n_1691)
);

NOR2xp67_ASAP7_75t_L g1692 ( 
.A(n_1686),
.B(n_1681),
.Y(n_1692)
);

NAND2xp33_ASAP7_75t_R g1693 ( 
.A(n_1688),
.B(n_1685),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1690),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1689),
.B(n_1683),
.Y(n_1695)
);

INVx1_ASAP7_75t_SL g1696 ( 
.A(n_1686),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1691),
.Y(n_1697)
);

XNOR2x1_ASAP7_75t_L g1698 ( 
.A(n_1696),
.B(n_1497),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1694),
.Y(n_1699)
);

NOR3xp33_ASAP7_75t_L g1700 ( 
.A(n_1695),
.B(n_1428),
.C(n_1456),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1692),
.B(n_1543),
.Y(n_1701)
);

OAI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1693),
.B1(n_1456),
.B2(n_1458),
.C(n_1450),
.Y(n_1702)
);

OAI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1697),
.A2(n_1538),
.B1(n_1491),
.B2(n_1514),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1700),
.A2(n_1538),
.B1(n_1492),
.B2(n_1500),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1702),
.Y(n_1705)
);

AO22x2_ASAP7_75t_L g1706 ( 
.A1(n_1705),
.A2(n_1699),
.B1(n_1698),
.B2(n_1703),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1706),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_SL g1708 ( 
.A1(n_1706),
.A2(n_1704),
.B1(n_1405),
.B2(n_1538),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1707),
.A2(n_1708),
.B1(n_1538),
.B2(n_1535),
.Y(n_1709)
);

AO21x1_ASAP7_75t_L g1710 ( 
.A1(n_1707),
.A2(n_1519),
.B(n_1535),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1709),
.A2(n_1542),
.B1(n_1535),
.B2(n_1519),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1710),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1711),
.B1(n_1355),
.B2(n_1543),
.Y(n_1713)
);

AOI21x1_ASAP7_75t_L g1714 ( 
.A1(n_1713),
.A2(n_1519),
.B(n_1542),
.Y(n_1714)
);

OA22x2_ASAP7_75t_L g1715 ( 
.A1(n_1714),
.A2(n_1519),
.B1(n_1542),
.B2(n_1535),
.Y(n_1715)
);

OAI221xp5_ASAP7_75t_R g1716 ( 
.A1(n_1715),
.A2(n_1355),
.B1(n_1542),
.B2(n_1491),
.C(n_1543),
.Y(n_1716)
);

AOI211xp5_ASAP7_75t_L g1717 ( 
.A1(n_1716),
.A2(n_1458),
.B(n_1405),
.C(n_1410),
.Y(n_1717)
);


endmodule