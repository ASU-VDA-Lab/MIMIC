module real_jpeg_4351_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_1),
.A2(n_144),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_1),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_1),
.A2(n_243),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_1),
.A2(n_95),
.B1(n_243),
.B2(n_355),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_1),
.A2(n_243),
.B1(n_377),
.B2(n_380),
.Y(n_376)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_2),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_2),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_3),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_94),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_3),
.A2(n_94),
.B1(n_189),
.B2(n_192),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_3),
.B(n_25),
.Y(n_287)
);

O2A1O1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_3),
.A2(n_343),
.B(n_345),
.C(n_349),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_3),
.B(n_367),
.C(n_369),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_3),
.B(n_159),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_3),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_3),
.B(n_79),
.Y(n_406)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_4),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_5),
.Y(n_184)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_5),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_5),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_5),
.Y(n_394)
);

INVx8_ASAP7_75t_L g402 ( 
.A(n_5),
.Y(n_402)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_6),
.Y(n_270)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_8),
.Y(n_437)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_9),
.Y(n_144)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_9),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_9),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_10),
.Y(n_440)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_11),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_12),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_12),
.A2(n_50),
.B1(n_125),
.B2(n_128),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_12),
.A2(n_50),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_12),
.A2(n_50),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_13),
.A2(n_38),
.B1(n_42),
.B2(n_45),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_13),
.A2(n_45),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_13),
.A2(n_45),
.B1(n_196),
.B2(n_200),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_13),
.A2(n_45),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_436),
.B(n_438),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_208),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_207),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_160),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_19),
.B(n_160),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_148),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_139),
.B2(n_140),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_63),
.B1(n_64),
.B2(n_138),
.Y(n_22)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_23),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_37),
.B(n_46),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_24),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_25),
.B(n_47),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_25),
.B(n_143),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_25),
.B(n_242),
.Y(n_253)
);

AO22x1_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_29),
.Y(n_274)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_31),
.Y(n_129)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_31),
.Y(n_268)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_34),
.Y(n_260)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_46),
.B(n_253),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_53),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_53),
.B(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_57),
.Y(n_276)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_98),
.B1(n_99),
.B2(n_137),
.Y(n_64)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_65),
.B(n_149),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_65),
.A2(n_137),
.B1(n_255),
.B2(n_263),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_65),
.B(n_252),
.C(n_255),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_88),
.B(n_89),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_66),
.A2(n_195),
.B(n_202),
.Y(n_194)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_67),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_67),
.B(n_90),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_67),
.B(n_354),
.Y(n_353)
);

NOR2x1_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_79),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_71),
.Y(n_201)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_71),
.Y(n_357)
);

AO22x1_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_80),
.B1(n_82),
.B2(n_86),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_78),
.Y(n_199)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_79),
.B(n_170),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_79),
.B(n_354),
.Y(n_371)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_83),
.Y(n_380)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_85),
.Y(n_235)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_87),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_87),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_88),
.B(n_89),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_88),
.A2(n_169),
.B(n_195),
.Y(n_236)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_93),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_94),
.A2(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_94),
.B(n_146),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g345 ( 
.A1(n_94),
.A2(n_346),
.B(n_348),
.Y(n_345)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_130),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_100),
.A2(n_151),
.B(n_159),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_100),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_123),
.Y(n_100)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_106),
.Y(n_347)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_122),
.Y(n_344)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_124),
.B(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_129),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_130),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_132),
.B(n_150),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_132),
.A2(n_150),
.B(n_159),
.Y(n_312)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_140),
.C(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_140),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_141),
.B(n_241),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_142),
.B(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_145),
.Y(n_272)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B(n_157),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_150),
.B(n_258),
.Y(n_285)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_152),
.Y(n_349)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_158),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_158),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_159),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_176),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_161),
.A2(n_164),
.B1(n_165),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_165),
.A2(n_166),
.B(n_175),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_167),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_169),
.B(n_371),
.Y(n_415)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_203),
.B(n_204),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_178),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_194),
.Y(n_178)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_203),
.B1(n_204),
.B2(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_179),
.A2(n_194),
.B1(n_203),
.B2(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_179),
.B(n_342),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_179),
.A2(n_203),
.B1(n_342),
.B2(n_418),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_185),
.B(n_188),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_180),
.B(n_188),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_180),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_180),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

BUFx8_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_183),
.B(n_231),
.Y(n_290)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_191),
.Y(n_379)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_194),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_198),
.Y(n_348)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_202),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_202),
.B(n_353),
.Y(n_382)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_245),
.B(n_435),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_210),
.B(n_213),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.C(n_220),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_214),
.A2(n_218),
.B1(n_219),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_214),
.Y(n_327)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_220),
.B(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_237),
.C(n_239),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_221),
.A2(n_222),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_236),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_223),
.B(n_236),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_224),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

INVx3_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_229),
.B(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_230),
.A2(n_278),
.B(n_282),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_237),
.B(n_239),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_238),
.B(n_257),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_427),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_316),
.C(n_332),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_304),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_291),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_250),
.B(n_291),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_264),
.C(n_283),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_251),
.B(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_264),
.A2(n_265),
.B1(n_283),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_277),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_266),
.B(n_277),
.Y(n_299)
);

AOI32xp33_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_269),
.A3(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_290),
.B(n_295),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.C(n_288),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_303),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_288),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_289),
.B(n_392),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_290),
.B(n_375),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_291),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_291),
.B(n_305),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.CI(n_298),
.CON(n_291),
.SN(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_296),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_297),
.B(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_304),
.A2(n_430),
.B(n_431),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_308),
.C(n_309),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_313),
.C(n_314),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_328),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_317),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_318),
.B(n_325),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.C(n_324),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_322),
.Y(n_330)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_329),
.B(n_331),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_358),
.B(n_426),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_334),
.B(n_337),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.C(n_350),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_338),
.B(n_422),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_341),
.A2(n_350),
.B1(n_351),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_341),
.Y(n_423)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_420),
.B(n_425),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_410),
.B(n_419),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_386),
.B(n_409),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_372),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_362),
.B(n_372),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_370),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_363),
.A2(n_364),
.B1(n_370),
.B2(n_389),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_370),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_381),
.Y(n_372)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_382),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_383),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_384),
.C(n_412),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_395),
.B(n_408),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_390),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_390),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_404),
.B(n_407),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_403),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

INVx4_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_406),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_413),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_416),
.C(n_417),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_424),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_421),
.B(n_424),
.Y(n_425)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_429),
.B(n_432),
.C(n_433),
.D(n_434),
.Y(n_427)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx6_ASAP7_75t_L g439 ( 
.A(n_437),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);


endmodule