module fake_jpeg_27737_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_3),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_56),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_0),
.B(n_1),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_0),
.B(n_1),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_41),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_48),
.B1(n_43),
.B2(n_39),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_47),
.B1(n_50),
.B2(n_41),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_63),
.B1(n_70),
.B2(n_8),
.Y(n_82)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_65),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_50),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_38),
.B1(n_50),
.B2(n_17),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_76),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_4),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_81),
.C(n_9),
.Y(n_93)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_7),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_7),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_8),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_22),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_89),
.A2(n_12),
.B1(n_23),
.B2(n_25),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_24),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_81),
.C(n_84),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_82),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_21),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_27),
.C(n_30),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_86),
.B(n_90),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_105),
.B(n_91),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_88),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_87),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_96),
.A3(n_101),
.B1(n_34),
.B2(n_36),
.C1(n_32),
.C2(n_33),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_66),
.B(n_101),
.C(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_66),
.Y(n_111)
);


endmodule