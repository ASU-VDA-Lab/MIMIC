module fake_netlist_1_928_n_30 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2xp67_ASAP7_75t_L g14 ( .A(n_7), .B(n_8), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_10), .Y(n_16) );
AND3x2_ASAP7_75t_L g17 ( .A(n_11), .B(n_12), .C(n_5), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
AOI22xp5_ASAP7_75t_L g19 ( .A1(n_13), .A2(n_3), .B1(n_1), .B2(n_9), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_15), .B(n_0), .Y(n_20) );
AOI21xp5_ASAP7_75t_L g21 ( .A1(n_16), .A2(n_4), .B(n_2), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_20), .B(n_18), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_17), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_18), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_24), .Y(n_26) );
INVxp67_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
NOR2x1p5_ASAP7_75t_L g28 ( .A(n_26), .B(n_23), .Y(n_28) );
OAI22xp5_ASAP7_75t_SL g29 ( .A1(n_27), .A2(n_19), .B1(n_18), .B2(n_3), .Y(n_29) );
AOI22xp33_ASAP7_75t_SL g30 ( .A1(n_29), .A2(n_28), .B1(n_14), .B2(n_2), .Y(n_30) );
endmodule