module fake_jpeg_17556_n_125 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_13),
.B(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_20),
.A3(n_22),
.B1(n_4),
.B2(n_3),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_22),
.Y(n_30)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_61),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_46),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_14),
.B1(n_23),
.B2(n_27),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_50),
.B1(n_54),
.B2(n_58),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_14),
.B1(n_27),
.B2(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_25),
.B1(n_24),
.B2(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g58 ( 
.A(n_28),
.B(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_24),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_5),
.Y(n_70)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_29),
.A2(n_21),
.B1(n_26),
.B2(n_19),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_26),
.C(n_19),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_26),
.C(n_16),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_34),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_53),
.B(n_58),
.Y(n_83)
);

XNOR2x1_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_47),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_78),
.Y(n_94)
);

AO22x2_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_49),
.B1(n_63),
.B2(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_6),
.Y(n_78)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_64),
.C(n_50),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_89),
.C(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_91),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_85),
.A2(n_88),
.B1(n_76),
.B2(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_69),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_49),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_43),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_57),
.C(n_52),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_93),
.C(n_67),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_76),
.B1(n_81),
.B2(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_100),
.Y(n_108)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_106),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_76),
.B1(n_66),
.B2(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_90),
.Y(n_114)
);

AO221x1_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_79),
.B1(n_66),
.B2(n_76),
.C(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_111),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_86),
.C(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_65),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_98),
.B1(n_86),
.B2(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_115),
.B(n_117),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_116),
.A2(n_118),
.A3(n_109),
.B1(n_112),
.B2(n_111),
.C1(n_96),
.C2(n_79),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_104),
.A3(n_100),
.B1(n_101),
.B2(n_97),
.C1(n_102),
.C2(n_105),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_10),
.A3(n_11),
.B1(n_68),
.B2(n_80),
.C1(n_117),
.C2(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_124),
.A2(n_68),
.B(n_122),
.C(n_123),
.Y(n_125)
);


endmodule