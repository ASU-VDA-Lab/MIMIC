module fake_jpeg_7079_n_174 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx2_ASAP7_75t_SL g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_15),
.B1(n_17),
.B2(n_20),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_14),
.B1(n_18),
.B2(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_15),
.B1(n_25),
.B2(n_22),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_14),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_23),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_15),
.B1(n_30),
.B2(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_65),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_44),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_13),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_50),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_80),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_59),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_62),
.B1(n_60),
.B2(n_66),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_74),
.B(n_18),
.Y(n_114)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_93),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_64),
.B1(n_42),
.B2(n_52),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_98),
.B1(n_80),
.B2(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_99),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_42),
.B1(n_54),
.B2(n_30),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_32),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_61),
.B1(n_54),
.B2(n_37),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_70),
.B1(n_76),
.B2(n_72),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_103),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_71),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_75),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_116),
.B(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_83),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_111),
.Y(n_125)
);

AOI221xp5_ASAP7_75t_L g119 ( 
.A1(n_112),
.A2(n_114),
.B1(n_115),
.B2(n_26),
.C(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_116),
.B1(n_61),
.B2(n_24),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_74),
.B(n_19),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

OAI322xp33_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_97),
.A3(n_99),
.B1(n_90),
.B2(n_93),
.C1(n_87),
.C2(n_85),
.Y(n_118)
);

AOI321xp33_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_124),
.A3(n_35),
.B1(n_29),
.B2(n_28),
.C(n_16),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_121),
.B(n_16),
.Y(n_141)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_32),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_40),
.C(n_53),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_126),
.C(n_16),
.Y(n_140)
);

OAI321xp33_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_26),
.A3(n_24),
.B1(n_19),
.B2(n_13),
.C(n_47),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g133 ( 
.A(n_123),
.B(n_16),
.C(n_13),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_35),
.C(n_40),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_104),
.B(n_101),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_127),
.B(n_133),
.C(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_128),
.B(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_136),
.Y(n_149)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_40),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_139),
.Y(n_146)
);

NOR4xp25_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_29),
.C(n_28),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_151),
.B(n_142),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_131),
.B(n_127),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_3),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_134),
.A2(n_130),
.B1(n_49),
.B2(n_13),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_140),
.B1(n_49),
.B2(n_27),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_29),
.C(n_16),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_27),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_157),
.B(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_160),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_155),
.B(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_159),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_9),
.B(n_12),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_8),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_11),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_10),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_49),
.B1(n_4),
.B2(n_5),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_167),
.A2(n_168),
.B(n_169),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_5),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_6),
.B(n_7),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_SL g171 ( 
.A(n_166),
.B(n_165),
.C(n_6),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_6),
.B(n_27),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

NAND2x1_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_27),
.Y(n_173)
);


endmodule