module fake_jpeg_27747_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_2),
.Y(n_7)
);

BUFx12_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_12),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_11),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_15),
.A2(n_13),
.B1(n_6),
.B2(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_17),
.B(n_20),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_10),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

MAJx2_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_8),
.C(n_1),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_27),
.C(n_18),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

AOI211xp5_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_35),
.B(n_16),
.C(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_33),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_36),
.C(n_40),
.Y(n_42)
);

AOI321xp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_37),
.A3(n_29),
.B1(n_14),
.B2(n_32),
.C(n_19),
.Y(n_43)
);


endmodule