module fake_jpeg_26760_n_195 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_195);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_41),
.Y(n_47)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_2),
.C(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_16),
.B(n_4),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_50),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_57),
.B1(n_59),
.B2(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_22),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_43),
.B1(n_38),
.B2(n_44),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_61),
.B1(n_31),
.B2(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_29),
.B1(n_28),
.B2(n_32),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_32),
.B1(n_21),
.B2(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_18),
.B1(n_19),
.B2(n_17),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_37),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_71),
.Y(n_91)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_33),
.B(n_31),
.C(n_17),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_83),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_43),
.C(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_80),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_45),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_47),
.B1(n_63),
.B2(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_33),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_25),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_28),
.B(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_39),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_90),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_57),
.B1(n_49),
.B2(n_53),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_99),
.B1(n_75),
.B2(n_76),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_73),
.B1(n_70),
.B2(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_6),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_39),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_102),
.B(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_56),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_106),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_28),
.B1(n_56),
.B2(n_7),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_5),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_5),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_5),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_108),
.B1(n_122),
.B2(n_99),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_104),
.A2(n_70),
.B1(n_77),
.B2(n_82),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_111),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_71),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_114),
.C(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_125),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_77),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_119),
.B1(n_89),
.B2(n_94),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_95),
.A2(n_72),
.B1(n_74),
.B2(n_69),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_102),
.B(n_101),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_74),
.B1(n_69),
.B2(n_66),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_91),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_103),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_135),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_129),
.B(n_138),
.CI(n_8),
.CON(n_153),
.SN(n_153)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_134),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_95),
.C(n_121),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_90),
.C(n_98),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_87),
.B1(n_105),
.B2(n_89),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_139),
.B1(n_120),
.B2(n_118),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_92),
.B1(n_116),
.B2(n_100),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_89),
.B1(n_92),
.B2(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_149),
.B1(n_128),
.B2(n_136),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_137),
.A2(n_125),
.B1(n_115),
.B2(n_114),
.Y(n_146)
);

OAI211xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_138),
.B(n_126),
.C(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_153),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_116),
.B1(n_92),
.B2(n_100),
.Y(n_149)
);

AO221x1_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_150)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_SL g152 ( 
.A(n_142),
.B(n_13),
.C(n_15),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_156),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_162),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_134),
.C(n_129),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_160),
.C(n_161),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_133),
.C(n_140),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_127),
.C(n_141),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_154),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_132),
.B(n_10),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_157),
.C(n_163),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_174),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_153),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_152),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

AOI31xp67_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_153),
.A3(n_155),
.B(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_166),
.B1(n_147),
.B2(n_149),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_177),
.C(n_178),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_148),
.B(n_144),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_9),
.B(n_10),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_11),
.B(n_12),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_10),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_171),
.C(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_185),
.B(n_187),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_11),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_182),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_11),
.B(n_180),
.C(n_178),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_190),
.B(n_191),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_188),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_192),
.Y(n_195)
);


endmodule