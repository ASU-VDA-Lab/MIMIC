module fake_jpeg_31177_n_60 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_60);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_60;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_0),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_31),
.C(n_32),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_8),
.C(n_16),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_7),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_22),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_35),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_38),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_27),
.B(n_24),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_5),
.C(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_25),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_6),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_5),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_50),
.B(n_13),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_12),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_11),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_55),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_47),
.C(n_51),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_53),
.C(n_39),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_58),
.B1(n_14),
.B2(n_18),
.Y(n_60)
);


endmodule