module fake_jpeg_15032_n_118 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_118);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_6),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_28),
.Y(n_35)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_22),
.B1(n_15),
.B2(n_21),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_22),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_15),
.B1(n_16),
.B2(n_12),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_22),
.B1(n_12),
.B2(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_21),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_45),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_52),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_0),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_13),
.B1(n_20),
.B2(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_50),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_51),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_49),
.B(n_52),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_40),
.B1(n_36),
.B2(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_20),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_70),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_72),
.B(n_62),
.Y(n_79)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_60),
.B(n_54),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_51),
.C(n_24),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_74),
.C(n_57),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_44),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_81),
.C(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_80),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_82),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_55),
.C(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_58),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_14),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_66),
.B1(n_75),
.B2(n_31),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_51),
.C(n_53),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_71),
.C(n_75),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_74),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_91),
.C(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_92),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_71),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_65),
.B1(n_34),
.B2(n_39),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_41),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_13),
.B1(n_40),
.B2(n_37),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_98),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_7),
.B(n_10),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_15),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_9),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_6),
.Y(n_104)
);

AOI211xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_107),
.B(n_101),
.C(n_9),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_93),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_5),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_95),
.B(n_3),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_111),
.B(n_4),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_1),
.B(n_4),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_112),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_103),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_113),
.A2(n_114),
.B1(n_37),
.B2(n_18),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_18),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_116),
.Y(n_118)
);


endmodule