module real_jpeg_23169_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_2),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_41),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_41),
.B1(n_53),
.B2(n_55),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_6),
.A2(n_25),
.B1(n_39),
.B2(n_42),
.Y(n_123)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_9),
.B1(n_32),
.B2(n_62),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_9),
.A2(n_32),
.B1(n_39),
.B2(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_32),
.B1(n_53),
.B2(n_55),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_9),
.B(n_52),
.C(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_9),
.B(n_51),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_9),
.B(n_39),
.C(n_72),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_9),
.B(n_24),
.C(n_36),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_9),
.B(n_11),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_9),
.B(n_87),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_9),
.B(n_103),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_11),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_96)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_126),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_125),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_104),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_16),
.B(n_104),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_78),
.C(n_88),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_17),
.A2(n_18),
.B1(n_78),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_47),
.B2(n_48),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_19),
.B(n_49),
.C(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_21),
.A2(n_33),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_21),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_27),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_22),
.A2(n_29),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_24),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_24),
.B(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_26),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_28),
.A2(n_98),
.B(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_29),
.B(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_33),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_33),
.A2(n_132),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_33),
.B(n_182),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_33),
.A2(n_110),
.B1(n_112),
.B2(n_132),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_33),
.B(n_110),
.C(n_203),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B(n_43),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_34),
.A2(n_43),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_34),
.B(n_137),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_38),
.A2(n_44),
.B1(n_45),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

OA22x2_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_42),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_39),
.B(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_44),
.B(n_136),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_45),
.Y(n_137)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_67),
.B1(n_68),
.B2(n_77),
.Y(n_48)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_49),
.A2(n_77),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_57),
.B(n_60),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_61),
.B1(n_64),
.B2(n_90),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_56),
.B1(n_58),
.B2(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_55),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_55),
.B(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_74),
.B(n_75),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_76),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_70),
.B(n_76),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_102),
.B(n_111),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_77),
.B(n_112),
.C(n_135),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_78),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_85),
.Y(n_108)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_85),
.A2(n_86),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_85),
.A2(n_86),
.B1(n_165),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_86),
.B(n_159),
.C(n_165),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_86),
.B(n_96),
.C(n_196),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_88),
.B(n_217),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.C(n_100),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_89),
.A2(n_100),
.B1(n_113),
.B2(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_95),
.A2(n_96),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_96),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_96),
.B(n_188),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_99),
.B(n_117),
.Y(n_170)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_152),
.C(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_100),
.A2(n_142),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_112),
.B1(n_135),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_155),
.B(n_214),
.C(n_219),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_144),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_128),
.B(n_144),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_140),
.B2(n_143),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_138),
.B2(n_139),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_131),
.B(n_139),
.C(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.C(n_151),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_145),
.A2(n_146),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_151),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_154),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_213),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_174),
.B(n_212),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_171),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_158),
.B(n_171),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_160),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_164),
.B(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_205),
.B(n_211),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_199),
.B(n_204),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_191),
.B(n_198),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_183),
.B(n_190),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B(n_189),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_192),
.B(n_193),
.Y(n_198)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_200),
.B(n_201),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_206),
.B(n_207),
.Y(n_211)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_216),
.Y(n_219)
);


endmodule