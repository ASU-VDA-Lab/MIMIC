module fake_netlist_6_4849_n_177 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_29, n_25, n_177);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_177;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_30;
wire n_79;
wire n_43;
wire n_171;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_R g37 ( 
.A(n_28),
.B(n_25),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_46),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_31),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_2),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_3),
.Y(n_60)
);

OR2x6_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_5),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_7),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_11),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_34),
.B1(n_32),
.B2(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_41),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

O2A1O1Ixp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_37),
.B(n_36),
.C(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_12),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_15),
.B(n_17),
.C(n_18),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_20),
.B(n_21),
.C(n_24),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_64),
.B1(n_61),
.B2(n_59),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_61),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_52),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_83),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_61),
.B(n_69),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_57),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_85),
.Y(n_92)
);

AND2x4_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_62),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_53),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_75),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_84),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_60),
.B(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

OR2x6_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_91),
.B(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_92),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_SL g108 ( 
.A(n_105),
.B(n_89),
.C(n_97),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_74),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_89),
.C(n_80),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_97),
.C(n_88),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_87),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_101),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

AO21x2_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_108),
.B(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_110),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_90),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_118),
.B(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_92),
.B1(n_100),
.B2(n_93),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_86),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_92),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_127),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_119),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_SL g143 ( 
.A(n_131),
.B(n_129),
.C(n_125),
.Y(n_143)
);

NOR4xp25_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_84),
.C(n_129),
.D(n_63),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_121),
.C(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_124),
.B1(n_92),
.B2(n_100),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_121),
.B1(n_100),
.B2(n_86),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_121),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_119),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_148),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_63),
.C(n_106),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_121),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_144),
.B1(n_92),
.B2(n_103),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_92),
.B1(n_164),
.B2(n_163),
.Y(n_167)
);

OR3x1_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_153),
.C(n_92),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_165),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_93),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_166),
.A2(n_93),
.B1(n_104),
.B2(n_71),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_26),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_172),
.B(n_157),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_173),
.B(n_168),
.Y(n_175)
);

OAI21x1_ASAP7_75t_SL g176 ( 
.A1(n_174),
.A2(n_167),
.B(n_171),
.Y(n_176)
);

OAI221xp5_ASAP7_75t_R g177 ( 
.A1(n_175),
.A2(n_176),
.B1(n_170),
.B2(n_166),
.C(n_71),
.Y(n_177)
);


endmodule