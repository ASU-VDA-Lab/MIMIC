module real_aes_6365_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_507, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_507;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_330;
wire n_388;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_297;
wire n_383;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_502;
wire n_434;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_484;
wire n_326;
wire n_492;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_SL g240 ( .A1(n_0), .A2(n_241), .B(n_242), .C(n_246), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_1), .B(n_235), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_2), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_3), .B(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_4), .A2(n_229), .B(n_331), .Y(n_330) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_5), .A2(n_202), .B(n_288), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_6), .A2(n_44), .B1(n_146), .B2(n_149), .Y(n_145) );
INVx1_ASAP7_75t_L g83 ( .A(n_7), .Y(n_83) );
INVx1_ASAP7_75t_L g192 ( .A(n_8), .Y(n_192) );
AND2x6_ASAP7_75t_L g227 ( .A(n_8), .B(n_190), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_8), .B(n_495), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_9), .A2(n_210), .B(n_227), .C(n_306), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_10), .A2(n_61), .B1(n_113), .B2(n_118), .Y(n_112) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_11), .A2(n_24), .B1(n_90), .B2(n_91), .Y(n_89) );
INVx1_ASAP7_75t_L g207 ( .A(n_12), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_13), .A2(n_39), .B1(n_162), .B2(n_166), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_14), .B(n_221), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_15), .A2(n_52), .B1(n_177), .B2(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_15), .Y(n_177) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_16), .A2(n_26), .B1(n_90), .B2(n_94), .Y(n_93) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_17), .A2(n_210), .B(n_272), .C(n_277), .Y(n_271) );
OAI22xp5_ASAP7_75t_SL g173 ( .A1(n_18), .A2(n_56), .B1(n_174), .B2(n_175), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_18), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_19), .A2(n_210), .B(n_277), .C(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_20), .Y(n_214) );
AOI22xp33_ASAP7_75t_SL g154 ( .A1(n_21), .A2(n_68), .B1(n_155), .B2(n_158), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_22), .A2(n_229), .B(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g212 ( .A(n_23), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_25), .A2(n_225), .B(n_256), .C(n_257), .Y(n_255) );
OAI221xp5_ASAP7_75t_L g183 ( .A1(n_26), .A2(n_38), .B1(n_50), .B2(n_184), .C(n_185), .Y(n_183) );
INVxp67_ASAP7_75t_L g186 ( .A(n_26), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_27), .B(n_293), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_28), .A2(n_80), .B1(n_169), .B2(n_170), .Y(n_79) );
CKINVDCx14_ASAP7_75t_R g169 ( .A(n_28), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_29), .B(n_270), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_30), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_31), .B(n_221), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_32), .B(n_229), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g316 ( .A1(n_33), .A2(n_225), .B(n_256), .C(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g243 ( .A(n_34), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_34), .A2(n_80), .B1(n_170), .B2(n_243), .Y(n_491) );
INVx1_ASAP7_75t_L g318 ( .A(n_35), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_36), .B(n_229), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_37), .Y(n_281) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_38), .A2(n_59), .B1(n_90), .B2(n_94), .Y(n_99) );
INVxp67_ASAP7_75t_L g187 ( .A(n_38), .Y(n_187) );
INVx1_ASAP7_75t_L g190 ( .A(n_40), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_41), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_42), .B(n_235), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g333 ( .A1(n_43), .A2(n_217), .B(n_276), .C(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g206 ( .A(n_45), .Y(n_206) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_46), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_47), .B(n_221), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_48), .B(n_222), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_49), .Y(n_129) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_50), .A2(n_66), .B1(n_90), .B2(n_91), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_51), .Y(n_238) );
INVx1_ASAP7_75t_L g178 ( .A(n_52), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_53), .B(n_260), .Y(n_273) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_54), .A2(n_210), .B(n_215), .C(n_225), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g332 ( .A(n_55), .Y(n_332) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_56), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_56), .B(n_259), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_57), .A2(n_72), .B1(n_136), .B2(n_141), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_58), .Y(n_265) );
INVx2_ASAP7_75t_L g204 ( .A(n_60), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_62), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_63), .B(n_245), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_64), .A2(n_80), .B1(n_170), .B2(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_64), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_65), .B(n_229), .Y(n_254) );
INVx1_ASAP7_75t_L g258 ( .A(n_67), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_69), .Y(n_105) );
INVxp67_ASAP7_75t_L g335 ( .A(n_70), .Y(n_335) );
INVx1_ASAP7_75t_L g90 ( .A(n_71), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_71), .Y(n_92) );
INVx1_ASAP7_75t_L g100 ( .A(n_73), .Y(n_100) );
INVx1_ASAP7_75t_L g216 ( .A(n_74), .Y(n_216) );
INVx1_ASAP7_75t_L g303 ( .A(n_75), .Y(n_303) );
AND2x2_ASAP7_75t_L g320 ( .A(n_76), .B(n_263), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_180), .B1(n_193), .B2(n_485), .C(n_490), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_171), .Y(n_78) );
INVx1_ASAP7_75t_L g170 ( .A(n_80), .Y(n_170) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_133), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_104), .C(n_122), .Y(n_81) );
OAI22xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_84), .B1(n_100), .B2(n_101), .Y(n_82) );
INVx1_ASAP7_75t_SL g84 ( .A(n_85), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
OR2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
INVx2_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
OR2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
AND2x2_ASAP7_75t_L g103 ( .A(n_88), .B(n_93), .Y(n_103) );
AND2x2_ASAP7_75t_L g140 ( .A(n_88), .B(n_128), .Y(n_140) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g109 ( .A(n_89), .B(n_93), .Y(n_109) );
AND2x2_ASAP7_75t_L g117 ( .A(n_89), .B(n_99), .Y(n_117) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_92), .Y(n_94) );
INVx2_ASAP7_75t_L g128 ( .A(n_93), .Y(n_128) );
INVx1_ASAP7_75t_L g168 ( .A(n_93), .Y(n_168) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NAND2x1p5_ASAP7_75t_L g102 ( .A(n_96), .B(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g165 ( .A(n_96), .B(n_140), .Y(n_165) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_98), .Y(n_96) );
INVx1_ASAP7_75t_L g111 ( .A(n_97), .Y(n_111) );
INVx1_ASAP7_75t_L g116 ( .A(n_97), .Y(n_116) );
INVx1_ASAP7_75t_L g121 ( .A(n_97), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_97), .B(n_99), .Y(n_144) );
AND2x2_ASAP7_75t_L g110 ( .A(n_98), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g139 ( .A(n_99), .B(n_121), .Y(n_139) );
BUFx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x4_ASAP7_75t_L g157 ( .A(n_103), .B(n_110), .Y(n_157) );
AND2x2_ASAP7_75t_L g160 ( .A(n_103), .B(n_139), .Y(n_160) );
OAI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_106), .B(n_112), .Y(n_104) );
INVx2_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x6_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x4_ASAP7_75t_L g119 ( .A(n_109), .B(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g148 ( .A(n_110), .B(n_140), .Y(n_148) );
AND2x6_ASAP7_75t_L g151 ( .A(n_110), .B(n_152), .Y(n_151) );
BUFx12f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g127 ( .A(n_116), .B(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g126 ( .A(n_117), .B(n_127), .Y(n_126) );
NAND2x1p5_ASAP7_75t_L g131 ( .A(n_117), .B(n_132), .Y(n_131) );
BUFx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_129), .B2(n_130), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx4f_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g132 ( .A(n_128), .Y(n_132) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_153), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_145), .Y(n_134) );
BUFx4f_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g142 ( .A(n_140), .B(n_143), .Y(n_142) );
BUFx2_ASAP7_75t_SL g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
OR2x6_ASAP7_75t_L g167 ( .A(n_144), .B(n_168), .Y(n_167) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx11_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_161), .Y(n_153) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx6_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx8_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx6_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B1(n_176), .B2(n_179), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_176), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_181), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
AND3x1_ASAP7_75t_SL g182 ( .A(n_183), .B(n_188), .C(n_191), .Y(n_182) );
INVxp67_ASAP7_75t_L g495 ( .A(n_183), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_188), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_188), .A2(n_499), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g505 ( .A(n_188), .Y(n_505) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_189), .B(n_192), .Y(n_501) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_SL g504 ( .A(n_191), .B(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_196), .B(n_428), .Y(n_195) );
AND4x1_ASAP7_75t_L g196 ( .A(n_197), .B(n_368), .C(n_383), .D(n_408), .Y(n_196) );
NOR2xp33_ASAP7_75t_SL g197 ( .A(n_198), .B(n_341), .Y(n_197) );
OAI21xp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_249), .B(n_321), .Y(n_198) );
AND2x2_ASAP7_75t_L g371 ( .A(n_199), .B(n_267), .Y(n_371) );
AND2x2_ASAP7_75t_L g384 ( .A(n_199), .B(n_266), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_199), .B(n_250), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_199), .Y(n_438) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_234), .Y(n_199) );
INVx2_ASAP7_75t_L g355 ( .A(n_200), .Y(n_355) );
BUFx2_ASAP7_75t_L g382 ( .A(n_200), .Y(n_382) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_208), .B(n_232), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_201), .B(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g235 ( .A(n_201), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_201), .B(n_265), .Y(n_264) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_201), .A2(n_302), .B(n_309), .Y(n_301) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_202), .A2(n_289), .B(n_290), .Y(n_288) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_202), .Y(n_329) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g311 ( .A(n_203), .Y(n_311) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
AND2x2_ASAP7_75t_SL g263 ( .A(n_204), .B(n_205), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_228), .Y(n_208) );
INVx5_ASAP7_75t_L g239 ( .A(n_210), .Y(n_239) );
AND2x6_ASAP7_75t_L g210 ( .A(n_211), .B(n_213), .Y(n_210) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_211), .Y(n_224) );
BUFx3_ASAP7_75t_L g247 ( .A(n_211), .Y(n_247) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g231 ( .A(n_212), .Y(n_231) );
INVx1_ASAP7_75t_L g297 ( .A(n_212), .Y(n_297) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_214), .Y(n_219) );
INVx3_ASAP7_75t_L g222 ( .A(n_214), .Y(n_222) );
AND2x2_ASAP7_75t_L g230 ( .A(n_214), .B(n_231), .Y(n_230) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_214), .Y(n_245) );
INVx1_ASAP7_75t_L g293 ( .A(n_214), .Y(n_293) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_220), .C(n_223), .Y(n_215) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g260 ( .A(n_219), .Y(n_260) );
INVx2_ASAP7_75t_L g241 ( .A(n_221), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_221), .B(n_335), .Y(n_334) );
INVx5_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_SL g237 ( .A1(n_226), .A2(n_238), .B(n_239), .C(n_240), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_226), .A2(n_239), .B(n_332), .C(n_333), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_226), .B(n_275), .Y(n_489) );
INVx4_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
AND2x4_ASAP7_75t_L g229 ( .A(n_227), .B(n_230), .Y(n_229) );
BUFx3_ASAP7_75t_L g277 ( .A(n_227), .Y(n_277) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_227), .B(n_230), .Y(n_304) );
BUFx2_ASAP7_75t_L g270 ( .A(n_229), .Y(n_270) );
INVx1_ASAP7_75t_L g276 ( .A(n_231), .Y(n_276) );
AND2x2_ASAP7_75t_L g322 ( .A(n_234), .B(n_267), .Y(n_322) );
INVx2_ASAP7_75t_L g338 ( .A(n_234), .Y(n_338) );
AND2x2_ASAP7_75t_L g347 ( .A(n_234), .B(n_266), .Y(n_347) );
AND2x2_ASAP7_75t_L g426 ( .A(n_234), .B(n_355), .Y(n_426) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_236), .B(n_248), .Y(n_234) );
INVx2_ASAP7_75t_L g256 ( .A(n_239), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
OAI322xp33_ASAP7_75t_L g490 ( .A1(n_243), .A2(n_491), .A3(n_492), .B1(n_496), .B2(n_497), .C1(n_502), .C2(n_504), .Y(n_490) );
INVx4_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_247), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_283), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_250), .B(n_353), .Y(n_391) );
INVx1_ASAP7_75t_L g479 ( .A(n_250), .Y(n_479) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_266), .Y(n_250) );
AND2x2_ASAP7_75t_L g337 ( .A(n_251), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g351 ( .A(n_251), .B(n_352), .Y(n_351) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_251), .Y(n_380) );
OR2x2_ASAP7_75t_L g412 ( .A(n_251), .B(n_354), .Y(n_412) );
AND2x2_ASAP7_75t_L g420 ( .A(n_251), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g453 ( .A(n_251), .B(n_422), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_251), .B(n_322), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_251), .B(n_382), .Y(n_478) );
AND2x2_ASAP7_75t_L g484 ( .A(n_251), .B(n_371), .Y(n_484) );
INVx5_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_L g344 ( .A(n_252), .Y(n_344) );
AND2x2_ASAP7_75t_L g374 ( .A(n_252), .B(n_354), .Y(n_374) );
AND2x2_ASAP7_75t_L g407 ( .A(n_252), .B(n_367), .Y(n_407) );
AND2x2_ASAP7_75t_L g427 ( .A(n_252), .B(n_267), .Y(n_427) );
AND2x2_ASAP7_75t_L g461 ( .A(n_252), .B(n_327), .Y(n_461) );
OR2x6_ASAP7_75t_L g252 ( .A(n_253), .B(n_264), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_263), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B(n_261), .C(n_262), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_259), .A2(n_262), .B(n_318), .C(n_319), .Y(n_317) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_259), .Y(n_488) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g279 ( .A(n_263), .Y(n_279) );
INVx1_ASAP7_75t_L g282 ( .A(n_263), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_263), .A2(n_315), .B(n_316), .Y(n_314) );
AND2x4_ASAP7_75t_L g367 ( .A(n_266), .B(n_338), .Y(n_367) );
AND2x2_ASAP7_75t_L g378 ( .A(n_266), .B(n_374), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_266), .B(n_354), .Y(n_417) );
INVx2_ASAP7_75t_L g432 ( .A(n_266), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_266), .B(n_366), .Y(n_455) );
AND2x2_ASAP7_75t_L g474 ( .A(n_266), .B(n_426), .Y(n_474) );
INVx5_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_267), .Y(n_373) );
AND2x2_ASAP7_75t_L g381 ( .A(n_267), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g422 ( .A(n_267), .B(n_338), .Y(n_422) );
OR2x6_ASAP7_75t_L g267 ( .A(n_268), .B(n_280), .Y(n_267) );
AOI21xp5_ASAP7_75t_SL g268 ( .A1(n_269), .A2(n_271), .B(n_278), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B(n_275), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_275), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_298), .Y(n_284) );
AND2x2_ASAP7_75t_L g345 ( .A(n_285), .B(n_328), .Y(n_345) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_286), .B(n_301), .Y(n_325) );
OR2x2_ASAP7_75t_L g358 ( .A(n_286), .B(n_328), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_286), .B(n_328), .Y(n_363) );
AND2x2_ASAP7_75t_L g390 ( .A(n_286), .B(n_327), .Y(n_390) );
AND2x2_ASAP7_75t_L g442 ( .A(n_286), .B(n_300), .Y(n_442) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_287), .B(n_312), .Y(n_350) );
AND2x2_ASAP7_75t_L g386 ( .A(n_287), .B(n_301), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .B(n_295), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_295), .A2(n_307), .B(n_308), .Y(n_306) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_298), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g376 ( .A(n_299), .B(n_358), .Y(n_376) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_312), .Y(n_299) );
OAI322xp33_ASAP7_75t_L g341 ( .A1(n_300), .A2(n_342), .A3(n_346), .B1(n_348), .B2(n_351), .C1(n_356), .C2(n_364), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_300), .B(n_327), .Y(n_349) );
OR2x2_ASAP7_75t_L g359 ( .A(n_300), .B(n_313), .Y(n_359) );
AND2x2_ASAP7_75t_L g361 ( .A(n_300), .B(n_313), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_300), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_300), .B(n_328), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_300), .B(n_457), .Y(n_456) );
INVx5_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_301), .B(n_345), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_305), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_312), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g339 ( .A(n_312), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_312), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g401 ( .A(n_312), .B(n_328), .Y(n_401) );
AOI211xp5_ASAP7_75t_SL g429 ( .A1(n_312), .A2(n_430), .B(n_433), .C(n_445), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_312), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g467 ( .A(n_312), .B(n_442), .Y(n_467) );
INVx5_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g395 ( .A(n_313), .B(n_328), .Y(n_395) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_313), .Y(n_404) );
AND2x2_ASAP7_75t_L g444 ( .A(n_313), .B(n_442), .Y(n_444) );
AND2x2_ASAP7_75t_SL g475 ( .A(n_313), .B(n_345), .Y(n_475) );
AND2x2_ASAP7_75t_L g482 ( .A(n_313), .B(n_441), .Y(n_482) );
OR2x6_ASAP7_75t_L g313 ( .A(n_314), .B(n_320), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B1(n_337), .B2(n_339), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_322), .B(n_344), .Y(n_392) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g340 ( .A(n_325), .Y(n_340) );
OR2x2_ASAP7_75t_L g400 ( .A(n_325), .B(n_401), .Y(n_400) );
OAI221xp5_ASAP7_75t_SL g448 ( .A1(n_325), .A2(n_449), .B1(n_451), .B2(n_452), .C(n_454), .Y(n_448) );
INVx2_ASAP7_75t_L g387 ( .A(n_326), .Y(n_387) );
AND2x2_ASAP7_75t_L g360 ( .A(n_327), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g450 ( .A(n_327), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_327), .B(n_442), .Y(n_463) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVxp67_ASAP7_75t_L g405 ( .A(n_328), .Y(n_405) );
AND2x2_ASAP7_75t_L g441 ( .A(n_328), .B(n_442), .Y(n_441) );
OA21x2_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B(n_336), .Y(n_328) );
AND2x2_ASAP7_75t_L g443 ( .A(n_337), .B(n_382), .Y(n_443) );
AND2x2_ASAP7_75t_L g353 ( .A(n_338), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_338), .B(n_411), .Y(n_410) );
NOR2xp33_ASAP7_75t_SL g424 ( .A(n_340), .B(n_387), .Y(n_424) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g430 ( .A(n_343), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
OR2x2_ASAP7_75t_L g416 ( .A(n_344), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g481 ( .A(n_344), .B(n_426), .Y(n_481) );
INVx2_ASAP7_75t_L g414 ( .A(n_345), .Y(n_414) );
NAND4xp25_ASAP7_75t_SL g477 ( .A(n_346), .B(n_478), .C(n_479), .D(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_347), .B(n_411), .Y(n_446) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_SL g483 ( .A(n_350), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g445 ( .A1(n_351), .A2(n_414), .B(n_418), .C(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g440 ( .A(n_353), .B(n_432), .Y(n_440) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_354), .Y(n_366) );
INVx1_ASAP7_75t_L g421 ( .A(n_354), .Y(n_421) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_355), .Y(n_398) );
AOI211xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B(n_360), .C(n_362), .Y(n_356) );
AND2x2_ASAP7_75t_L g377 ( .A(n_357), .B(n_361), .Y(n_377) );
OAI322xp33_ASAP7_75t_SL g415 ( .A1(n_357), .A2(n_416), .A3(n_418), .B1(n_419), .B2(n_423), .C1(n_424), .C2(n_425), .Y(n_415) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g437 ( .A(n_359), .B(n_363), .Y(n_437) );
INVx1_ASAP7_75t_L g418 ( .A(n_361), .Y(n_418) );
INVx1_ASAP7_75t_SL g436 ( .A(n_363), .Y(n_436) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_375), .B1(n_377), .B2(n_378), .C1(n_379), .C2(n_507), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_372), .Y(n_369) );
OAI322xp33_ASAP7_75t_L g458 ( .A1(n_370), .A2(n_432), .A3(n_437), .B1(n_459), .B2(n_460), .C1(n_462), .C2(n_463), .Y(n_458) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_371), .A2(n_385), .B1(n_409), .B2(n_413), .C(n_415), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
OAI222xp33_ASAP7_75t_L g388 ( .A1(n_376), .A2(n_389), .B1(n_391), .B2(n_392), .C1(n_393), .C2(n_396), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_378), .A2(n_385), .B1(n_455), .B2(n_456), .Y(n_454) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AOI211xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_388), .C(n_399), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g464 ( .A1(n_385), .A2(n_422), .B(n_465), .C(n_468), .Y(n_464) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g394 ( .A(n_386), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g457 ( .A(n_390), .Y(n_457) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_397), .B(n_422), .Y(n_451) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B(n_406), .Y(n_399) );
OAI221xp5_ASAP7_75t_SL g468 ( .A1(n_400), .A2(n_469), .B1(n_470), .B2(n_471), .C(n_472), .Y(n_468) );
INVxp33_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_404), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_411), .B(n_422), .Y(n_462) );
INVx2_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AND2x2_ASAP7_75t_L g473 ( .A(n_426), .B(n_432), .Y(n_473) );
AND4x1_ASAP7_75t_L g428 ( .A(n_429), .B(n_447), .C(n_464), .D(n_476), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI221xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_435), .B1(n_437), .B2(n_438), .C(n_439), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B1(n_443), .B2(n_444), .Y(n_439) );
INVx1_ASAP7_75t_L g469 ( .A(n_440), .Y(n_469) );
INVx1_ASAP7_75t_SL g459 ( .A(n_444), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g447 ( .A(n_448), .B(n_458), .Y(n_447) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_460), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_467), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_482), .B1(n_483), .B2(n_484), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g500 ( .A(n_488), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_498), .Y(n_497) );
endmodule