module fake_jpeg_7790_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_25),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_23),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_65),
.Y(n_75)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_70),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_0),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_49),
.B(n_55),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_52),
.C(n_9),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_53),
.B1(n_46),
.B2(n_40),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_81),
.B1(n_88),
.B2(n_8),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_57),
.B1(n_56),
.B2(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_1),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_6),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_47),
.B1(n_43),
.B2(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_59),
.B1(n_58),
.B2(n_48),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_95),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_2),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_3),
.B1(n_4),
.B2(n_51),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_3),
.C(n_4),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_113),
.B1(n_103),
.B2(n_102),
.Y(n_114)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_108),
.B1(n_100),
.B2(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_105),
.C(n_110),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_93),
.B1(n_76),
.B2(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_104),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_101),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_101),
.C(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_122),
.B(n_10),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_11),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_13),
.C(n_15),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_16),
.B(n_19),
.Y(n_126)
);

OAI31xp33_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_20),
.A3(n_21),
.B(n_26),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_127),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_129)
);


endmodule