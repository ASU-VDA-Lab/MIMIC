module real_jpeg_19993_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_270, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_270;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_197;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_0),
.A2(n_3),
.B1(n_37),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_49),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_49),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_0),
.A2(n_5),
.B1(n_49),
.B2(n_62),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_1),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_1),
.A2(n_5),
.B1(n_19),
.B2(n_62),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_2),
.A2(n_3),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_20),
.B1(n_21),
.B2(n_42),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_42),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_5),
.B1(n_42),
.B2(n_62),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_2),
.A2(n_20),
.B(n_45),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_2),
.B(n_52),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_2),
.A2(n_5),
.B(n_10),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_2),
.B(n_24),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_2),
.A2(n_27),
.B(n_28),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_3),
.A2(n_7),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_3),
.A2(n_35),
.B(n_42),
.C(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_4),
.Y(n_99)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_4),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_5),
.A2(n_10),
.B1(n_60),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_7),
.B1(n_38),
.B2(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_5),
.B(n_106),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_7),
.A2(n_20),
.B1(n_21),
.B2(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_227)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_35),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_34),
.B(n_37),
.C(n_44),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_82),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_81),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_64),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_16),
.B(n_64),
.Y(n_81)
);

BUFx24_ASAP7_75t_SL g268 ( 
.A(n_16),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_33),
.CI(n_46),
.CON(n_16),
.SN(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_22),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_18),
.A2(n_24),
.B1(n_30),
.B2(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_20),
.A2(n_29),
.B(n_42),
.C(n_172),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_21),
.A2(n_25),
.B(n_28),
.C(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_28),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_23),
.B(n_80),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_24),
.A2(n_79),
.B(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_25),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_25),
.A2(n_31),
.B1(n_80),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_27),
.A2(n_42),
.B(n_60),
.C(n_148),
.Y(n_147)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_31),
.B(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_36),
.B(n_39),
.Y(n_33)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_34),
.B(n_43),
.Y(n_246)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_45),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_48),
.B(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_43),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_42),
.B(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_42),
.B(n_61),
.Y(n_154)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.C(n_55),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_47),
.A2(n_67),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_47),
.B(n_116),
.C(n_117),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_47),
.A2(n_67),
.B1(n_108),
.B2(n_127),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_47),
.B(n_108),
.C(n_222),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_51),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_55),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_58),
.A2(n_61),
.B1(n_93),
.B2(n_96),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_58),
.A2(n_61),
.B1(n_63),
.B2(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_61),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_62),
.B(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_72),
.C(n_74),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_260)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.C(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_72),
.A2(n_73),
.B1(n_125),
.B2(n_128),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_72),
.A2(n_73),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_72),
.A2(n_73),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_108),
.C(n_110),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_73),
.B(n_209),
.C(n_211),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_74),
.B(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_252),
.A3(n_261),
.B1(n_266),
.B2(n_267),
.C(n_270),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_235),
.B(n_251),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_216),
.B(n_234),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_137),
.B(n_197),
.C(n_215),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_123),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_87),
.B(n_123),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_112),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_107),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_89),
.B(n_107),
.C(n_112),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_97),
.B2(n_98),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_90),
.A2(n_91),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_90),
.A2(n_91),
.B1(n_108),
.B2(n_127),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_90),
.B(n_98),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_91),
.B(n_147),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_91),
.B(n_108),
.C(n_170),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B(n_95),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_95),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_99),
.B(n_105),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_99),
.A2(n_100),
.B1(n_105),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_122),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_102),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_105),
.B1(n_106),
.B2(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_110),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_114),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_132),
.C(n_134),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_114),
.A2(n_116),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_114),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_114),
.B(n_241),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_154),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_130),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_121),
.B(n_162),
.C(n_165),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.C(n_131),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_124),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_125),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_129),
.B(n_131),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_144),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_196),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_191),
.B(n_195),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_179),
.B(n_190),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_167),
.B(n_178),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_157),
.B(n_166),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_149),
.B(n_156),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_145),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_153),
.B(n_155),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_159),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_165),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_165),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_182),
.C(n_189),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_165),
.B(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_177),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_171),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_176),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_181),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_188),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_199),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_213),
.B2(n_214),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_208),
.C(n_214),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_213),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_217),
.B(n_218),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_233),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_225),
.C(n_233),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_229),
.B1(n_230),
.B2(n_232),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_226),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_230),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_230),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_245),
.B(n_248),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_237),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_249),
.B2(n_250),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_243),
.C(n_250),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_254),
.C(n_257),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_254),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_257),
.A2(n_258),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_262),
.B(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);


endmodule