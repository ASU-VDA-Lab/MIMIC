module real_jpeg_13129_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_0),
.A2(n_19),
.B1(n_20),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_0),
.A2(n_29),
.B1(n_52),
.B2(n_54),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_0),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_24),
.C(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_0),
.B(n_87),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_0),
.A2(n_8),
.B(n_23),
.C(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_0),
.B(n_37),
.C(n_40),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_0),
.B(n_18),
.Y(n_136)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

AO22x1_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_10),
.A2(n_26),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_10),
.A2(n_19),
.B1(n_20),
.B2(n_26),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_10),
.A2(n_26),
.B1(n_39),
.B2(n_40),
.Y(n_82)
);

XNOR2x2_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_106),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_104),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_92),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_92),
.Y(n_105)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_14),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_59),
.CI(n_76),
.CON(n_14),
.SN(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_32),
.C(n_46),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_16),
.A2(n_32),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_16),
.A2(n_70),
.B1(n_75),
.B2(n_97),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_22),
.B(n_27),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_17),
.A2(n_22),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

O2A1O1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_21),
.B(n_24),
.C(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_19),
.A2(n_20),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_19),
.A2(n_21),
.B(n_29),
.Y(n_113)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_20),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_24),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_23),
.A2(n_24),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_29),
.B(n_63),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_29),
.B(n_43),
.Y(n_148)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_43),
.B(n_44),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_45),
.Y(n_73)
);

AO22x1_ASAP7_75t_SL g125 ( 
.A1(n_34),
.A2(n_38),
.B1(n_45),
.B2(n_72),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

AO22x1_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_39),
.B(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_63),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OA21x2_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_71),
.B(n_73),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_47),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OA21x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_55),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_56),
.A2(n_57),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_63),
.B(n_65),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_67),
.B1(n_69),
.B2(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_65),
.B(n_82),
.Y(n_101)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_97),
.C(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_70),
.B(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_70),
.A2(n_75),
.B1(n_132),
.B2(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_83),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_81),
.A2(n_99),
.B1(n_135),
.B2(n_138),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_81),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_81),
.B(n_148),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_81),
.B(n_125),
.C(n_137),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_89),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_101),
.C(n_102),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.C(n_100),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_93),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_98),
.B(n_100),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_101),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_159),
.B(n_163),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_128),
.B(n_158),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_116),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_109),
.B(n_116),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_110),
.A2(n_111),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_122),
.B2(n_123),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_125),
.C(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_119),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_127),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_152),
.B(n_157),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_139),
.B(n_151),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_136),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_143),
.B(n_150),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_147),
.B(n_149),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_153),
.B(n_154),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_160),
.B(n_161),
.Y(n_163)
);


endmodule