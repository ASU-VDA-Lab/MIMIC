module fake_jpeg_10620_n_126 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_126);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_35),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_19),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_35),
.B1(n_25),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_21),
.B1(n_18),
.B2(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_16),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_30),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_64),
.Y(n_82)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_57),
.B1(n_17),
.B2(n_3),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_14),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_32),
.B1(n_16),
.B2(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_63),
.Y(n_83)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_24),
.Y(n_64)
);

OA22x2_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_36),
.B1(n_34),
.B2(n_22),
.Y(n_65)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_17),
.B(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_36),
.B(n_34),
.C(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_22),
.Y(n_71)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_1),
.B(n_4),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_84),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_50),
.B1(n_65),
.B2(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_92),
.B1(n_68),
.B2(n_78),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_61),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_91),
.C(n_93),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_64),
.C(n_59),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_50),
.C(n_65),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_77),
.B(n_1),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_84),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_70),
.C(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_63),
.Y(n_96)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_81),
.B(n_71),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_101),
.C(n_91),
.Y(n_110)
);

OAI322xp33_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_72),
.A3(n_78),
.B1(n_76),
.B2(n_77),
.C1(n_75),
.C2(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_4),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_105),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_93),
.B1(n_85),
.B2(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_112),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_103),
.B1(n_99),
.B2(n_73),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_116),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_107),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_108),
.B1(n_110),
.B2(n_97),
.Y(n_120)
);

AOI31xp67_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_111),
.A3(n_106),
.B(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_119),
.B(n_120),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_73),
.B1(n_116),
.B2(n_88),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_121),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_123),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_122),
.B(n_11),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_125),
.Y(n_126)
);


endmodule