module fake_jpeg_2981_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_0),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_56),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_58),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_63),
.B1(n_57),
.B2(n_55),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_37),
.B1(n_51),
.B2(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_48),
.B1(n_43),
.B2(n_46),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_52),
.B1(n_56),
.B2(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_38),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_72),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_68),
.A2(n_54),
.B1(n_53),
.B2(n_58),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_60),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_56),
.B1(n_57),
.B2(n_55),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_61),
.B1(n_39),
.B2(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_76),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_65),
.B1(n_57),
.B2(n_55),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_35),
.B1(n_14),
.B2(n_22),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_49),
.B(n_42),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_2),
.B(n_3),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_97),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_0),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_101),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_99),
.A2(n_112),
.B(n_95),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_72),
.B1(n_71),
.B2(n_76),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_104),
.B1(n_107),
.B2(n_110),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_2),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_39),
.B1(n_15),
.B2(n_20),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_96),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_109),
.B(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_108),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_4),
.B(n_5),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_4),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_107),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_95),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_125),
.C(n_104),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_83),
.B(n_24),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_119),
.A2(n_120),
.B(n_104),
.Y(n_127)
);

FAx1_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_83),
.CI(n_27),
.CON(n_120),
.SN(n_120)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_125),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_28),
.C(n_31),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_127),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_130),
.C(n_117),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_131),
.B1(n_116),
.B2(n_124),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_13),
.C(n_30),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_134),
.C(n_120),
.Y(n_136)
);

AOI31xp33_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_120),
.A3(n_118),
.B(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_29),
.B(n_33),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_8),
.B(n_10),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_10),
.C(n_11),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_11),
.C(n_12),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_12),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_142),
.Y(n_143)
);


endmodule