module fake_jpeg_27040_n_121 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx11_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_17),
.Y(n_38)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx12_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_23),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_28),
.B1(n_13),
.B2(n_24),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_28),
.B1(n_36),
.B2(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_43),
.Y(n_60)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_13),
.B1(n_11),
.B2(n_25),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_37),
.A3(n_31),
.B1(n_33),
.B2(n_26),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_39),
.C(n_32),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_31),
.C(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_40),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_63),
.B(n_72),
.Y(n_78)
);

AND2x6_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_9),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_72),
.C(n_2),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_53),
.B(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_71),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_9),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_53),
.B(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_75),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_78),
.B(n_82),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_69),
.A2(n_18),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_15),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_44),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_87),
.Y(n_93)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_52),
.C(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_91),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_75),
.B(n_79),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_49),
.C(n_22),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_2),
.B(n_3),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_79),
.B(n_49),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_88),
.B1(n_85),
.B2(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_99),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_85),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_103),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_49),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_105),
.C(n_101),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_94),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_105),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_111),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_108),
.B(n_107),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_109),
.B(n_50),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_113),
.A2(n_26),
.B1(n_50),
.B2(n_14),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_116),
.B(n_29),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_118),
.B(n_5),
.C(n_6),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_22),
.C(n_27),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_6),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_7),
.Y(n_121)
);


endmodule