module fake_jpeg_13527_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_47),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_28),
.A2(n_24),
.B1(n_27),
.B2(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_25),
.B1(n_21),
.B2(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_46),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_28),
.B(n_0),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_27),
.B1(n_33),
.B2(n_28),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_59),
.B1(n_41),
.B2(n_30),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_56),
.B(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_27),
.B1(n_20),
.B2(n_25),
.Y(n_59)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_23),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_29),
.B1(n_21),
.B2(n_17),
.Y(n_100)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_18),
.CON(n_67),
.SN(n_67)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_71),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_70),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_74),
.B(n_76),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_25),
.B1(n_32),
.B2(n_19),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_25),
.B1(n_32),
.B2(n_19),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

FAx1_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_18),
.CI(n_40),
.CON(n_84),
.SN(n_84)
);

NAND2xp33_ASAP7_75t_SL g127 ( 
.A(n_84),
.B(n_72),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_32),
.B1(n_19),
.B2(n_18),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_48),
.B1(n_42),
.B2(n_17),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_57),
.Y(n_122)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_45),
.B1(n_46),
.B2(n_27),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_93),
.B1(n_52),
.B2(n_17),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_48),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_66),
.A2(n_21),
.B1(n_29),
.B2(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_31),
.C(n_40),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_99),
.C(n_52),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_98),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_53),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_101),
.B1(n_78),
.B2(n_50),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_29),
.B1(n_20),
.B2(n_42),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_71),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_120),
.C(n_128),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_61),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_112),
.Y(n_136)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_61),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_117),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_122),
.B1(n_78),
.B2(n_100),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_80),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_58),
.C(n_69),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_17),
.A3(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_84),
.B(n_16),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_74),
.B(n_75),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_81),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_81),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_86),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_86),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_50),
.Y(n_128)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_133),
.B(n_143),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_141),
.C(n_111),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_142),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_116),
.B(n_108),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_106),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_120),
.C(n_69),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_73),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_149),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_152),
.B(n_156),
.Y(n_162)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_102),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_90),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_88),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_128),
.Y(n_159)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_185),
.C(n_187),
.Y(n_209)
);

INVxp33_ASAP7_75t_SL g165 ( 
.A(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_165),
.B(n_180),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_181),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_110),
.B(n_109),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_189),
.B(n_191),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_110),
.B1(n_126),
.B2(n_109),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_179),
.B1(n_149),
.B2(n_150),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_151),
.B1(n_122),
.B2(n_136),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_193),
.B1(n_138),
.B2(n_154),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_128),
.B(n_84),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_122),
.B1(n_84),
.B2(n_89),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_132),
.A2(n_130),
.B1(n_91),
.B2(n_97),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_182),
.A2(n_193),
.B(n_173),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_190),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_108),
.C(n_97),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_50),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_187),
.B(n_145),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_153),
.A2(n_72),
.B(n_97),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_135),
.B(n_11),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_155),
.B(n_142),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_137),
.A2(n_57),
.B1(n_91),
.B2(n_72),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_208),
.B1(n_172),
.B2(n_188),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_204),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_191),
.A2(n_133),
.B(n_146),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_175),
.A2(n_134),
.B1(n_156),
.B2(n_157),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_213),
.C(n_218),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_158),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_192),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_145),
.C(n_147),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_215),
.B(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_57),
.C(n_160),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_222),
.Y(n_228)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_164),
.B(n_148),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_199),
.C(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_160),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_168),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_242),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_34),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_210),
.B(n_162),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_235),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_249),
.B1(n_250),
.B2(n_198),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_179),
.B(n_188),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_241),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_181),
.A3(n_171),
.B1(n_190),
.B2(n_194),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_198),
.A2(n_189),
.B(n_182),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_9),
.B(n_16),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_201),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_248),
.B(n_208),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_197),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_63),
.B1(n_9),
.B2(n_10),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_213),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_240),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_258),
.B1(n_240),
.B2(n_246),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_254),
.A2(n_243),
.B1(n_229),
.B2(n_225),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_218),
.C(n_221),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_257),
.C(n_259),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_200),
.C(n_196),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_212),
.B1(n_238),
.B2(n_249),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_196),
.C(n_220),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_223),
.C(n_216),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_214),
.C(n_207),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_205),
.C(n_202),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_230),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_250),
.B(n_238),
.Y(n_277)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_34),
.C(n_8),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_272),
.C(n_232),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_34),
.C(n_9),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_256),
.C(n_263),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_260),
.B1(n_262),
.B2(n_272),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_277),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_285),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_259),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_241),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_247),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_245),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_287),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_244),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_7),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_264),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_293),
.B(n_0),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_270),
.B(n_265),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_298),
.B(n_302),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_275),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_284),
.B1(n_287),
.B2(n_278),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_224),
.B(n_239),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_283),
.A2(n_239),
.B(n_10),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_279),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_13),
.Y(n_314)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_304),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_306),
.B(n_309),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_296),
.A2(n_286),
.B1(n_275),
.B2(n_11),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_307),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_290),
.B(n_15),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_312),
.Y(n_318)
);

NOR2x1_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_14),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_314),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_292),
.B(n_14),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_34),
.C(n_13),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_299),
.C(n_1),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_7),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_315),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_304),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_323),
.Y(n_330)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_305),
.A2(n_291),
.A3(n_297),
.B1(n_301),
.B2(n_302),
.C1(n_298),
.C2(n_294),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_320),
.A2(n_322),
.B1(n_324),
.B2(n_1),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_291),
.A3(n_308),
.B1(n_311),
.B2(n_299),
.C1(n_309),
.C2(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_308),
.C(n_34),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_327),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_323),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_329),
.C(n_331),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_321),
.B(n_2),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_2),
.C(n_3),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_3),
.Y(n_332)
);

OAI31xp33_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_325),
.A3(n_324),
.B(n_5),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_334),
.Y(n_336)
);

OAI321xp33_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_330),
.A3(n_333),
.B1(n_335),
.B2(n_327),
.C(n_5),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_4),
.B(n_5),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_4),
.B(n_5),
.Y(n_339)
);


endmodule