module fake_ariane_2192_n_921 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_921);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_921;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_919;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_352;
wire n_206;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_872;
wire n_774;
wire n_916;
wire n_254;
wire n_596;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_203;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_852;
wire n_793;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_170),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_33),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_71),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_64),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_103),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_23),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_16),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_51),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_16),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_169),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_36),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_40),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_81),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_133),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_165),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_67),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_41),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_72),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_77),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_126),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_124),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_135),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_118),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_89),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_148),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_144),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_37),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_7),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_177),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_19),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_99),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_17),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_59),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_20),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_123),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_142),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_117),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_23),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_146),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_5),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_35),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_49),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_44),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_66),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_38),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_122),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_13),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_86),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_17),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_140),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_24),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_32),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_84),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_171),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_172),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_141),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_25),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_107),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_115),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_62),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_200),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_192),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_192),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_192),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_192),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_197),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_200),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_200),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_208),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_L g271 ( 
.A(n_195),
.B(n_0),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_183),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_208),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_187),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_L g279 ( 
.A(n_224),
.B(n_0),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_188),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_184),
.B(n_1),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_R g282 ( 
.A(n_185),
.B(n_30),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_194),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_189),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_187),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_228),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_229),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_199),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_232),
.B(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_211),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_215),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_244),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_231),
.B(n_1),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_233),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_249),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_240),
.B(n_2),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_191),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_191),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_245),
.B(n_2),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_260),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_269),
.B(n_251),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_285),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_284),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_261),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_256),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_263),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_263),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_R g322 ( 
.A(n_264),
.B(n_186),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_266),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_265),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_269),
.B(n_253),
.Y(n_325)
);

AND3x2_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_248),
.C(n_252),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_284),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_275),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_273),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_288),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_296),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_296),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_280),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_267),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_264),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_269),
.B(n_202),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_278),
.B(n_209),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_270),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_303),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_270),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_304),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_301),
.Y(n_349)
);

CKINVDCx8_ASAP7_75t_R g350 ( 
.A(n_268),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_R g351 ( 
.A(n_282),
.B(n_247),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_262),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_274),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_262),
.Y(n_355)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_285),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_299),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_294),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_294),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_276),
.B(n_213),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_346),
.B(n_259),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_315),
.B(n_283),
.Y(n_363)
);

AND3x2_ASAP7_75t_L g364 ( 
.A(n_310),
.B(n_297),
.C(n_281),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_344),
.Y(n_365)
);

BUFx6f_ASAP7_75t_SL g366 ( 
.A(n_343),
.Y(n_366)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_221),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_289),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_311),
.B(n_291),
.Y(n_369)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_331),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_300),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_340),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_344),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_311),
.B(n_292),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_351),
.B(n_322),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_359),
.B(n_293),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_353),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_341),
.B(n_290),
.Y(n_383)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_325),
.B(n_221),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_311),
.Y(n_385)
);

OR2x6_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_271),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_329),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_323),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

BUFx4f_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

OR2x2_ASAP7_75t_SL g393 ( 
.A(n_319),
.B(n_305),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_309),
.B(n_295),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_323),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_356),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_324),
.A2(n_332),
.B1(n_335),
.B2(n_325),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_352),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_306),
.B(n_298),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_356),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

OR2x6_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_279),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_352),
.B(n_302),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_356),
.Y(n_407)
);

BUFx8_ASAP7_75t_SL g408 ( 
.A(n_328),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g409 ( 
.A(n_320),
.B(n_221),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_307),
.B(n_246),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_345),
.B(n_190),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_321),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_347),
.A2(n_242),
.B1(n_237),
.B2(n_236),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_316),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_313),
.B(n_221),
.Y(n_417)
);

BUFx10_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_321),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_340),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_318),
.B(n_196),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_308),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_338),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_354),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_314),
.B(n_198),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_354),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_357),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_316),
.B(n_356),
.Y(n_433)
);

OR2x6_ASAP7_75t_L g434 ( 
.A(n_339),
.B(n_3),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_429),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_429),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_391),
.B(n_317),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_389),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_391),
.B(n_316),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_374),
.B(n_326),
.Y(n_440)
);

NAND2x1p5_ASAP7_75t_L g441 ( 
.A(n_378),
.B(n_317),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_408),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_403),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_403),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_374),
.B(n_201),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_380),
.B(n_334),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_368),
.B(n_334),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_375),
.B(n_203),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_392),
.B(n_204),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_3),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_397),
.B(n_205),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_363),
.B(n_206),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_395),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_348),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_421),
.A2(n_212),
.B(n_210),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_434),
.A2(n_328),
.B1(n_348),
.B2(n_235),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_400),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_368),
.B(n_4),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_398),
.B(n_214),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_363),
.B(n_216),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_414),
.B(n_217),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_423),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_420),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_412),
.B(n_4),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_371),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_362),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_399),
.A2(n_234),
.B1(n_227),
.B2(n_226),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_421),
.B(n_5),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_399),
.B(n_219),
.Y(n_472)
);

O2A1O1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_369),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_416),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_418),
.B(n_225),
.Y(n_475)
);

NOR3xp33_ASAP7_75t_L g476 ( 
.A(n_431),
.B(n_6),
.C(n_8),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_428),
.B(n_9),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_404),
.B(n_369),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_428),
.B(n_9),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_411),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_377),
.B(n_10),
.Y(n_482)
);

AO22x1_ASAP7_75t_L g483 ( 
.A1(n_422),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_418),
.B(n_11),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_392),
.B(n_13),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_392),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_410),
.B(n_14),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_425),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_377),
.B(n_14),
.Y(n_489)
);

NOR3xp33_ASAP7_75t_L g490 ( 
.A(n_422),
.B(n_15),
.C(n_18),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_404),
.B(n_372),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_382),
.B(n_15),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_430),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_404),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_390),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_410),
.B(n_18),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_387),
.B(n_19),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_366),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_381),
.B(n_20),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_366),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_394),
.B(n_182),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_402),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_367),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_394),
.B(n_26),
.Y(n_504)
);

A2O1A1Ixp33_ASAP7_75t_L g505 ( 
.A1(n_406),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_424),
.B(n_426),
.Y(n_506)
);

AOI221xp5_ASAP7_75t_L g507 ( 
.A1(n_383),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C(n_31),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_SL g509 ( 
.A(n_415),
.B(n_29),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_432),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_367),
.B(n_181),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_367),
.B(n_34),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_434),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_419),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_367),
.B(n_45),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_367),
.B(n_179),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_415),
.B(n_365),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_449),
.A2(n_427),
.B(n_433),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_486),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_447),
.A2(n_433),
.B(n_417),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_443),
.A2(n_417),
.B(n_415),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_442),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_438),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_451),
.A2(n_386),
.B1(n_434),
.B2(n_393),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_517),
.A2(n_373),
.B(n_376),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_L g526 ( 
.A1(n_451),
.A2(n_379),
.B(n_364),
.C(n_384),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_493),
.B(n_370),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_465),
.Y(n_528)
);

AOI21x1_ASAP7_75t_L g529 ( 
.A1(n_517),
.A2(n_386),
.B(n_384),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_506),
.A2(n_384),
.B(n_407),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_469),
.B(n_386),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_445),
.A2(n_407),
.B(n_401),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_460),
.B(n_364),
.Y(n_533)
);

O2A1O1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_487),
.A2(n_384),
.B(n_409),
.C(n_396),
.Y(n_534)
);

O2A1O1Ixp33_ASAP7_75t_L g535 ( 
.A1(n_496),
.A2(n_384),
.B(n_409),
.C(n_396),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_471),
.A2(n_401),
.B(n_370),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_471),
.A2(n_409),
.B(n_47),
.Y(n_537)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_467),
.B(n_409),
.C(n_48),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_482),
.A2(n_409),
.B(n_50),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_455),
.A2(n_46),
.B(n_52),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_466),
.A2(n_53),
.B(n_54),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_478),
.B(n_55),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_478),
.B(n_56),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_489),
.A2(n_57),
.B(n_58),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_472),
.B(n_60),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_468),
.B(n_61),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_444),
.A2(n_63),
.B(n_65),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_444),
.A2(n_439),
.B(n_477),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_439),
.A2(n_68),
.B(n_69),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_480),
.A2(n_70),
.B(n_73),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_446),
.B(n_74),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_435),
.A2(n_75),
.B(n_76),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_448),
.B(n_78),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_467),
.B(n_79),
.C(n_80),
.Y(n_554)
);

AO21x1_ASAP7_75t_L g555 ( 
.A1(n_485),
.A2(n_175),
.B(n_83),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_448),
.B(n_82),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_504),
.A2(n_497),
.B(n_492),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_446),
.B(n_85),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_479),
.B(n_174),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_436),
.A2(n_514),
.B(n_510),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_457),
.A2(n_87),
.B(n_88),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_450),
.A2(n_90),
.B(n_91),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_450),
.A2(n_92),
.B(n_93),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_462),
.A2(n_94),
.B(n_95),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_437),
.A2(n_96),
.B(n_97),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_495),
.A2(n_98),
.B(n_100),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_454),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_461),
.B(n_101),
.Y(n_568)
);

O2A1O1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_499),
.A2(n_102),
.B(n_104),
.C(n_105),
.Y(n_569)
);

O2A1O1Ixp33_ASAP7_75t_L g570 ( 
.A1(n_479),
.A2(n_106),
.B(n_108),
.C(n_109),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_456),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_459),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_486),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_508),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_498),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_453),
.A2(n_110),
.B(n_112),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_461),
.B(n_113),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_474),
.Y(n_578)
);

OAI21x1_ASAP7_75t_L g579 ( 
.A1(n_530),
.A2(n_488),
.B(n_515),
.Y(n_579)
);

OAI21x1_ASAP7_75t_L g580 ( 
.A1(n_521),
.A2(n_516),
.B(n_512),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_548),
.A2(n_511),
.B(n_485),
.Y(n_581)
);

AO31x2_ASAP7_75t_L g582 ( 
.A1(n_536),
.A2(n_491),
.A3(n_505),
.B(n_440),
.Y(n_582)
);

NOR2x1_ASAP7_75t_L g583 ( 
.A(n_531),
.B(n_475),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_571),
.Y(n_584)
);

A2O1A1Ixp33_ASAP7_75t_L g585 ( 
.A1(n_551),
.A2(n_558),
.B(n_559),
.C(n_537),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_520),
.A2(n_501),
.B(n_473),
.Y(n_586)
);

AOI21x1_ASAP7_75t_L g587 ( 
.A1(n_545),
.A2(n_509),
.B(n_464),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_528),
.B(n_481),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_524),
.B(n_441),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_557),
.A2(n_491),
.B(n_486),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_573),
.Y(n_591)
);

AOI21x1_ASAP7_75t_SL g592 ( 
.A1(n_568),
.A2(n_481),
.B(n_463),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_574),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_525),
.A2(n_502),
.B(n_503),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_522),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_578),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_575),
.B(n_441),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_532),
.A2(n_486),
.B(n_452),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_518),
.A2(n_502),
.B(n_507),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_546),
.A2(n_484),
.B(n_470),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_533),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_557),
.A2(n_577),
.B(n_543),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_542),
.A2(n_544),
.B(n_537),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_560),
.B(n_494),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_529),
.A2(n_500),
.B(n_498),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_539),
.A2(n_500),
.B(n_513),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_544),
.A2(n_483),
.B(n_490),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_523),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_567),
.B(n_458),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_572),
.Y(n_610)
);

AOI21x1_ASAP7_75t_L g611 ( 
.A1(n_539),
.A2(n_476),
.B(n_116),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_550),
.A2(n_114),
.B(n_119),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_526),
.B(n_120),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_519),
.B(n_121),
.Y(n_614)
);

OAI21x1_ASAP7_75t_L g615 ( 
.A1(n_561),
.A2(n_125),
.B(n_127),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_553),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_556),
.A2(n_136),
.B1(n_138),
.B2(n_143),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_527),
.B(n_173),
.Y(n_618)
);

NOR2x1_ASAP7_75t_SL g619 ( 
.A(n_573),
.B(n_145),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_519),
.B(n_147),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_576),
.A2(n_149),
.B(n_151),
.Y(n_621)
);

AOI21x1_ASAP7_75t_SL g622 ( 
.A1(n_570),
.A2(n_555),
.B(n_565),
.Y(n_622)
);

AOI21xp33_ASAP7_75t_L g623 ( 
.A1(n_554),
.A2(n_152),
.B(n_153),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_527),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_549),
.A2(n_154),
.B(n_155),
.Y(n_625)
);

OAI21x1_ASAP7_75t_SL g626 ( 
.A1(n_569),
.A2(n_156),
.B(n_157),
.Y(n_626)
);

OAI21x1_ASAP7_75t_L g627 ( 
.A1(n_547),
.A2(n_158),
.B(n_159),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_573),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_534),
.B(n_160),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_588),
.B(n_564),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_588),
.B(n_563),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_584),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_591),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_591),
.Y(n_634)
);

A2O1A1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_607),
.A2(n_562),
.B(n_538),
.C(n_535),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_593),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_595),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_589),
.B(n_601),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_608),
.Y(n_639)
);

CKINVDCx8_ASAP7_75t_R g640 ( 
.A(n_591),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_609),
.B(n_541),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_624),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_596),
.B(n_610),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_628),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_585),
.A2(n_540),
.B(n_566),
.C(n_552),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_603),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_646)
);

INVxp67_ASAP7_75t_SL g647 ( 
.A(n_628),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_597),
.B(n_164),
.Y(n_648)
);

O2A1O1Ixp5_ASAP7_75t_L g649 ( 
.A1(n_602),
.A2(n_166),
.B(n_167),
.C(n_168),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_590),
.B(n_604),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_602),
.A2(n_586),
.B(n_598),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_590),
.B(n_604),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_583),
.B(n_628),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_606),
.A2(n_600),
.B(n_599),
.C(n_613),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_618),
.B(n_605),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_582),
.B(n_613),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_582),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_579),
.A2(n_580),
.B(n_581),
.Y(n_658)
);

O2A1O1Ixp5_ASAP7_75t_SL g659 ( 
.A1(n_623),
.A2(n_629),
.B(n_617),
.C(n_616),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_582),
.B(n_619),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_611),
.A2(n_617),
.B1(n_616),
.B2(n_629),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_625),
.A2(n_587),
.B1(n_621),
.B2(n_620),
.Y(n_662)
);

OR2x2_ASAP7_75t_SL g663 ( 
.A(n_614),
.B(n_620),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_594),
.B(n_614),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_623),
.A2(n_621),
.B1(n_615),
.B2(n_612),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_627),
.Y(n_666)
);

AOI21xp33_ASAP7_75t_L g667 ( 
.A1(n_626),
.A2(n_592),
.B(n_622),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_593),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_588),
.B(n_388),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_601),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_590),
.B(n_588),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_588),
.B(n_456),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_593),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_593),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_589),
.B(n_575),
.Y(n_675)
);

NOR2xp67_ASAP7_75t_SL g676 ( 
.A(n_595),
.B(n_442),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_595),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_595),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_589),
.B(n_624),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_591),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_SL g681 ( 
.A1(n_638),
.A2(n_670),
.B1(n_669),
.B2(n_637),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_644),
.Y(n_682)
);

OAI22xp33_ASAP7_75t_L g683 ( 
.A1(n_672),
.A2(n_641),
.B1(n_675),
.B2(n_661),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_632),
.B(n_668),
.Y(n_684)
);

NAND2x1p5_ASAP7_75t_L g685 ( 
.A(n_632),
.B(n_679),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_636),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_673),
.B(n_674),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_SL g688 ( 
.A1(n_661),
.A2(n_656),
.B1(n_660),
.B2(n_675),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_633),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_643),
.Y(n_690)
);

AOI21x1_ASAP7_75t_L g691 ( 
.A1(n_662),
.A2(n_651),
.B(n_666),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_656),
.A2(n_675),
.B1(n_639),
.B2(n_671),
.Y(n_692)
);

AO21x1_ASAP7_75t_L g693 ( 
.A1(n_671),
.A2(n_630),
.B(n_631),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_677),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_652),
.Y(n_695)
);

AOI21x1_ASAP7_75t_L g696 ( 
.A1(n_662),
.A2(n_664),
.B(n_658),
.Y(n_696)
);

AO21x2_ASAP7_75t_L g697 ( 
.A1(n_665),
.A2(n_654),
.B(n_667),
.Y(n_697)
);

OAI21xp33_ASAP7_75t_L g698 ( 
.A1(n_659),
.A2(n_667),
.B(n_645),
.Y(n_698)
);

BUFx4f_ASAP7_75t_SL g699 ( 
.A(n_678),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_642),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_657),
.A2(n_648),
.B1(n_653),
.B2(n_655),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_647),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_SL g703 ( 
.A1(n_657),
.A2(n_655),
.B1(n_663),
.B2(n_678),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_633),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_640),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_634),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_633),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_635),
.A2(n_646),
.B(n_649),
.Y(n_708)
);

NAND2x1p5_ASAP7_75t_L g709 ( 
.A(n_680),
.B(n_676),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_680),
.A2(n_458),
.B1(n_524),
.B2(n_434),
.Y(n_710)
);

AOI21x1_ASAP7_75t_L g711 ( 
.A1(n_661),
.A2(n_662),
.B(n_651),
.Y(n_711)
);

BUFx12f_ASAP7_75t_L g712 ( 
.A(n_637),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_638),
.A2(n_334),
.B1(n_317),
.B2(n_333),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_633),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_672),
.B(n_670),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_668),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_668),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_640),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_640),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_669),
.B(n_672),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_L g721 ( 
.A1(n_659),
.A2(n_585),
.B(n_607),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_650),
.Y(n_722)
);

INVxp33_ASAP7_75t_L g723 ( 
.A(n_638),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_668),
.Y(n_724)
);

BUFx2_ASAP7_75t_R g725 ( 
.A(n_637),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_640),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_668),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_650),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_638),
.A2(n_334),
.B1(n_317),
.B2(n_333),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_668),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_670),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_722),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_685),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_711),
.A2(n_691),
.B(n_696),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_722),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_728),
.Y(n_736)
);

AO21x2_ASAP7_75t_L g737 ( 
.A1(n_721),
.A2(n_683),
.B(n_693),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_685),
.Y(n_738)
);

INVx8_ASAP7_75t_L g739 ( 
.A(n_705),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_695),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_686),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_697),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_716),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_717),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_700),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_683),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_692),
.B(n_720),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_687),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_684),
.B(n_692),
.Y(n_749)
);

HB1xp67_ASAP7_75t_L g750 ( 
.A(n_702),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_688),
.B(n_715),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_688),
.B(n_723),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_R g753 ( 
.A(n_705),
.B(n_718),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_714),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_714),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_724),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_723),
.B(n_730),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_727),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_690),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_SL g760 ( 
.A1(n_708),
.A2(n_698),
.B(n_709),
.Y(n_760)
);

OAI22xp33_ASAP7_75t_L g761 ( 
.A1(n_713),
.A2(n_729),
.B1(n_726),
.B2(n_719),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_689),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_703),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_706),
.Y(n_764)
);

AO31x2_ASAP7_75t_L g765 ( 
.A1(n_707),
.A2(n_704),
.A3(n_703),
.B(n_682),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_681),
.B(n_714),
.Y(n_766)
);

OAI21x1_ASAP7_75t_SL g767 ( 
.A1(n_701),
.A2(n_710),
.B(n_709),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_731),
.B(n_694),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_726),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_718),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_719),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_712),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_751),
.B(n_710),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_754),
.Y(n_774)
);

AO21x1_ASAP7_75t_SL g775 ( 
.A1(n_763),
.A2(n_732),
.B(n_741),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_751),
.B(n_725),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_735),
.B(n_712),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_742),
.B(n_699),
.Y(n_778)
);

INVxp67_ASAP7_75t_R g779 ( 
.A(n_766),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_735),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_740),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_732),
.B(n_699),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_740),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_741),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_761),
.B(n_772),
.Y(n_785)
);

INVx3_ASAP7_75t_SL g786 ( 
.A(n_739),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_748),
.B(n_746),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_745),
.B(n_752),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_745),
.B(n_752),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_759),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_745),
.B(n_764),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_750),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_736),
.B(n_764),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_736),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_734),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_736),
.B(n_764),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_746),
.B(n_737),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_737),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_759),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_788),
.B(n_768),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_797),
.A2(n_760),
.B(n_770),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_785),
.A2(n_760),
.B1(n_763),
.B2(n_771),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_R g803 ( 
.A(n_786),
.B(n_753),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_792),
.B(n_757),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_798),
.B(n_769),
.C(n_770),
.Y(n_805)
);

NAND3xp33_ASAP7_75t_L g806 ( 
.A(n_798),
.B(n_769),
.C(n_770),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_788),
.B(n_768),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_789),
.B(n_766),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_792),
.B(n_757),
.Y(n_809)
);

OA21x2_ASAP7_75t_L g810 ( 
.A1(n_797),
.A2(n_734),
.B(n_787),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_789),
.B(n_765),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_SL g812 ( 
.A1(n_797),
.A2(n_747),
.B(n_762),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_787),
.B(n_748),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_791),
.B(n_762),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_791),
.B(n_737),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_779),
.B(n_765),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_780),
.B(n_737),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_778),
.B(n_771),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_780),
.B(n_747),
.Y(n_819)
);

NAND4xp25_ASAP7_75t_L g820 ( 
.A(n_782),
.B(n_771),
.C(n_754),
.D(n_755),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_790),
.B(n_749),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_779),
.B(n_765),
.Y(n_822)
);

OAI221xp5_ASAP7_75t_L g823 ( 
.A1(n_773),
.A2(n_749),
.B1(n_756),
.B2(n_758),
.C(n_733),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_790),
.B(n_755),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_782),
.B(n_756),
.C(n_758),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_L g826 ( 
.A(n_778),
.B(n_733),
.C(n_754),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_799),
.B(n_755),
.Y(n_827)
);

NAND4xp25_ASAP7_75t_L g828 ( 
.A(n_777),
.B(n_784),
.C(n_776),
.D(n_795),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_813),
.B(n_799),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_803),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_800),
.B(n_777),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_819),
.B(n_815),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_807),
.B(n_778),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_808),
.B(n_775),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_821),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_811),
.B(n_775),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_804),
.Y(n_837)
);

AND2x4_ASAP7_75t_SL g838 ( 
.A(n_816),
.B(n_776),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_809),
.B(n_784),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_811),
.B(n_796),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_824),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_812),
.B(n_796),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_816),
.B(n_796),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_828),
.B(n_739),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_810),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_829),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_838),
.B(n_822),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_839),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_837),
.Y(n_849)
);

OAI33xp33_ASAP7_75t_L g850 ( 
.A1(n_832),
.A2(n_817),
.A3(n_802),
.B1(n_825),
.B2(n_827),
.B3(n_814),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_836),
.B(n_818),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_836),
.B(n_818),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_841),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_845),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_841),
.Y(n_855)
);

INVxp33_ASAP7_75t_L g856 ( 
.A(n_847),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_847),
.B(n_838),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_847),
.B(n_834),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_848),
.B(n_832),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_849),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_851),
.B(n_834),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_853),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_852),
.B(n_833),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_850),
.Y(n_864)
);

CKINVDCx16_ASAP7_75t_R g865 ( 
.A(n_857),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_862),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_860),
.Y(n_867)
);

BUFx12f_ASAP7_75t_L g868 ( 
.A(n_857),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_859),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_866),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_869),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_867),
.A2(n_864),
.B1(n_856),
.B2(n_845),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_865),
.A2(n_856),
.B1(n_857),
.B2(n_830),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_870),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_871),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_873),
.B(n_868),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_872),
.B(n_867),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_873),
.B(n_850),
.Y(n_878)
);

NOR3xp33_ASAP7_75t_SL g879 ( 
.A(n_877),
.B(n_844),
.C(n_820),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_878),
.A2(n_845),
.B(n_854),
.C(n_842),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_876),
.B(n_854),
.C(n_858),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_875),
.B(n_858),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_874),
.A2(n_861),
.B(n_863),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_876),
.B(n_861),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_874),
.Y(n_885)
);

NOR3xp33_ASAP7_75t_L g886 ( 
.A(n_880),
.B(n_823),
.C(n_855),
.Y(n_886)
);

AOI211xp5_ASAP7_75t_L g887 ( 
.A1(n_881),
.A2(n_884),
.B(n_882),
.C(n_885),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_883),
.B(n_863),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_SL g889 ( 
.A(n_879),
.B(n_822),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_880),
.B(n_846),
.C(n_801),
.Y(n_890)
);

AND3x2_ASAP7_75t_L g891 ( 
.A(n_885),
.B(n_773),
.C(n_831),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_L g892 ( 
.A(n_887),
.B(n_805),
.C(n_806),
.Y(n_892)
);

AOI211xp5_ASAP7_75t_L g893 ( 
.A1(n_889),
.A2(n_803),
.B(n_826),
.C(n_786),
.Y(n_893)
);

NOR4xp25_ASAP7_75t_L g894 ( 
.A(n_888),
.B(n_835),
.C(n_843),
.D(n_831),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_891),
.B(n_833),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_886),
.B(n_835),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_890),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_896),
.Y(n_898)
);

INVxp67_ASAP7_75t_L g899 ( 
.A(n_897),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_895),
.A2(n_892),
.B1(n_893),
.B2(n_894),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_L g901 ( 
.A(n_897),
.B(n_810),
.C(n_795),
.Y(n_901)
);

NOR2x1_ASAP7_75t_L g902 ( 
.A(n_897),
.B(n_843),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_902),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_898),
.B(n_810),
.Y(n_904)
);

CKINVDCx16_ASAP7_75t_R g905 ( 
.A(n_900),
.Y(n_905)
);

NAND4xp75_ASAP7_75t_L g906 ( 
.A(n_899),
.B(n_840),
.C(n_739),
.D(n_793),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_903),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_905),
.B(n_901),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_907),
.Y(n_909)
);

XNOR2xp5_ASAP7_75t_L g910 ( 
.A(n_908),
.B(n_906),
.Y(n_910)
);

OAI221xp5_ASAP7_75t_L g911 ( 
.A1(n_909),
.A2(n_904),
.B1(n_786),
.B2(n_840),
.C(n_795),
.Y(n_911)
);

NOR4xp25_ASAP7_75t_L g912 ( 
.A(n_910),
.B(n_795),
.C(n_783),
.D(n_781),
.Y(n_912)
);

OA21x2_ASAP7_75t_L g913 ( 
.A1(n_911),
.A2(n_734),
.B(n_767),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_912),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_914),
.A2(n_739),
.B1(n_767),
.B2(n_743),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_913),
.A2(n_743),
.B(n_744),
.Y(n_916)
);

CKINVDCx16_ASAP7_75t_R g917 ( 
.A(n_916),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_917),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_918),
.A2(n_913),
.B1(n_915),
.B2(n_739),
.Y(n_919)
);

OAI221xp5_ASAP7_75t_R g920 ( 
.A1(n_919),
.A2(n_774),
.B1(n_754),
.B2(n_755),
.C(n_765),
.Y(n_920)
);

AOI211xp5_ASAP7_75t_L g921 ( 
.A1(n_920),
.A2(n_738),
.B(n_794),
.C(n_793),
.Y(n_921)
);


endmodule