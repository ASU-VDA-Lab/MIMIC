module fake_netlist_1_6449_n_9 (n_3, n_1, n_2, n_0, n_9);
input n_3;
input n_1;
input n_2;
input n_0;
output n_9;
wire n_6;
wire n_4;
wire n_5;
wire n_7;
wire n_8;
NAND3xp33_ASAP7_75t_SL g4 ( .A(n_2), .B(n_3), .C(n_1), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
AOI222xp33_ASAP7_75t_L g7 ( .A1(n_6), .A2(n_4), .B1(n_5), .B2(n_2), .C1(n_3), .C2(n_0), .Y(n_7) );
AOI211xp5_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_0), .B(n_1), .C(n_2), .Y(n_8) );
AOI21xp33_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_1), .B(n_3), .Y(n_9) );
endmodule