module real_aes_15954_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_34;
wire n_12;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_35;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
wire n_33;
wire n_36;
INVx2_ASAP7_75t_L g29 ( .A(n_0), .Y(n_29) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_2), .B(n_7), .Y(n_16) );
AND2x2_ASAP7_75t_L g14 ( .A(n_3), .B(n_15), .Y(n_14) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_3), .Y(n_25) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_4), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_5), .B(n_27), .Y(n_26) );
INVx1_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_9), .A2(n_17), .B(n_22), .Y(n_8) );
NOR2xp33_ASAP7_75t_L g9 ( .A(n_10), .B(n_12), .Y(n_9) );
INVx1_ASAP7_75t_L g33 ( .A(n_10), .Y(n_33) );
INVx1_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
INVxp67_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_14), .B(n_16), .Y(n_13) );
HB1xp67_ASAP7_75t_L g32 ( .A(n_15), .Y(n_32) );
INVx1_ASAP7_75t_L g24 ( .A(n_16), .Y(n_24) );
A2O1A1Ixp33_ASAP7_75t_L g22 ( .A1(n_17), .A2(n_23), .B(n_33), .C(n_34), .Y(n_22) );
INVx1_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
AOI221xp5_ASAP7_75t_SL g23 ( .A1(n_24), .A2(n_25), .B1(n_26), .B2(n_30), .C(n_31), .Y(n_23) );
INVx1_ASAP7_75t_L g30 ( .A(n_25), .Y(n_30) );
NOR2xp33_ASAP7_75t_L g35 ( .A(n_25), .B(n_31), .Y(n_35) );
INVxp67_ASAP7_75t_SL g36 ( .A(n_26), .Y(n_36) );
INVx2_ASAP7_75t_SL g27 ( .A(n_28), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
INVx1_ASAP7_75t_L g31 ( .A(n_32), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_35), .B(n_36), .Y(n_34) );
endmodule