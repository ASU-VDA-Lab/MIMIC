module fake_jpeg_2252_n_154 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_SL g48 ( 
.A(n_9),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_51),
.Y(n_52)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_48),
.B1(n_55),
.B2(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_54),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_38),
.B1(n_37),
.B2(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_52),
.A2(n_38),
.B1(n_41),
.B2(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_20),
.Y(n_98)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_84),
.Y(n_88)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_39),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_42),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_62),
.B1(n_1),
.B2(n_2),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_44),
.B1(n_41),
.B2(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_70),
.B1(n_62),
.B2(n_2),
.Y(n_86)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_44),
.Y(n_85)
);

XNOR2x1_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_19),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_3),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_8),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_22),
.C(n_33),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_116),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_5),
.B(n_8),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_9),
.B(n_10),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_108),
.B(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_24),
.B1(n_32),
.B2(n_30),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_120),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_117),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_118),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_17),
.C(n_27),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_116),
.B(n_126),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_25),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_133),
.Y(n_138)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_103),
.C(n_112),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_137),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_120),
.C(n_111),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_114),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_139),
.A2(n_140),
.B1(n_124),
.B2(n_122),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_104),
.B1(n_113),
.B2(n_10),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_122),
.B1(n_133),
.B2(n_131),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_130),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_143),
.B1(n_129),
.B2(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_145),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_144),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_144),
.B(n_127),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_134),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_13),
.B(n_14),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_152),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_15),
.Y(n_154)
);


endmodule