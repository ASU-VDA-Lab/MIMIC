module fake_jpeg_19660_n_87 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_87);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_87;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_0),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_32),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_51),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_37),
.B1(n_33),
.B2(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_1),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_18),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_59),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx2_ASAP7_75t_SL g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_1),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_2),
.B(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_20),
.B1(n_4),
.B2(n_8),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_71),
.B1(n_11),
.B2(n_14),
.Y(n_75)
);

AO21x2_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_60),
.B(n_13),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_68),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_72),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_79),
.B1(n_15),
.B2(n_16),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_74),
.B1(n_66),
.B2(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_22),
.B(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_24),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_25),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_26),
.Y(n_87)
);


endmodule