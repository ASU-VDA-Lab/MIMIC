module fake_jpeg_11389_n_183 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_183);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_183;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_24),
.C(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_18),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx2_ASAP7_75t_SL g56 ( 
.A(n_40),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_18),
.B1(n_32),
.B2(n_22),
.Y(n_63)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_57),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_42),
.B1(n_38),
.B2(n_36),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_63),
.B1(n_43),
.B2(n_40),
.Y(n_70)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_25),
.B1(n_22),
.B2(n_16),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_39),
.B1(n_34),
.B2(n_20),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_25),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_74),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_37),
.B(n_40),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_79),
.B(n_21),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_42),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_75),
.Y(n_90)
);

FAx1_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_43),
.CI(n_32),
.CON(n_74),
.SN(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_30),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_84),
.Y(n_99)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_19),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_20),
.B(n_19),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_34),
.B1(n_52),
.B2(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_104),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_56),
.B(n_8),
.C(n_10),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_106),
.B1(n_107),
.B2(n_74),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_46),
.B1(n_21),
.B2(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_105),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_46),
.B(n_21),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_21),
.B1(n_2),
.B2(n_5),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_72),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_88),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_80),
.C(n_75),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

BUFx4f_ASAP7_75t_SL g138 ( 
.A(n_115),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_79),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_77),
.C(n_68),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_119),
.Y(n_131)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_124),
.B1(n_107),
.B2(n_95),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_104),
.B1(n_105),
.B2(n_94),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_125),
.B(n_126),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_127),
.A2(n_78),
.B(n_71),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_101),
.B(n_97),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_121),
.B(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_135),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_133),
.B1(n_114),
.B2(n_117),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_98),
.B1(n_74),
.B2(n_96),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_120),
.A2(n_106),
.B1(n_87),
.B2(n_66),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_66),
.B1(n_68),
.B2(n_76),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_140),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_115),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_134),
.A2(n_112),
.B(n_119),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_150),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_127),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_149),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_110),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_113),
.C(n_83),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_118),
.C(n_1),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_135),
.B1(n_128),
.B2(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g160 ( 
.A(n_146),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_149),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_150),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_167),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_166),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_162),
.B(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_145),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_158),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_156),
.B1(n_159),
.B2(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_138),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_139),
.C(n_158),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_173),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_175),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_152),
.A3(n_141),
.B1(n_125),
.B2(n_138),
.C1(n_93),
.C2(n_14),
.Y(n_175)
);

AOI31xp67_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_141),
.A3(n_138),
.B(n_13),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_171),
.B1(n_93),
.B2(n_7),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_179),
.B1(n_176),
.B2(n_172),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_181),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_6),
.Y(n_183)
);


endmodule