module fake_jpeg_18770_n_176 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_35),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_27),
.B(n_5),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_65),
.B1(n_68),
.B2(n_71),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_93),
.B(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_86),
.A2(n_68),
.B1(n_65),
.B2(n_76),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_74),
.B1(n_77),
.B2(n_60),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_79),
.B1(n_74),
.B2(n_60),
.Y(n_103)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_77),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_114),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_104),
.B1(n_98),
.B2(n_90),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_109),
.Y(n_116)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_112),
.Y(n_118)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_73),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_76),
.B1(n_69),
.B2(n_75),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_61),
.B(n_53),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_0),
.B(n_1),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_122),
.B1(n_78),
.B2(n_67),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_54),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_2),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_103),
.A2(n_98),
.B1(n_52),
.B2(n_90),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_73),
.B(n_54),
.C(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_125),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_59),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_3),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_107),
.B1(n_114),
.B2(n_63),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_129),
.A2(n_63),
.B1(n_58),
.B2(n_4),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_139),
.B1(n_129),
.B2(n_119),
.Y(n_143)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_141),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_8),
.B(n_9),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_78),
.C(n_67),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_128),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_133),
.B1(n_12),
.B2(n_13),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_11),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_140),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_6),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_143),
.B(n_146),
.Y(n_158)
);

XOR2x2_ASAP7_75t_SL g144 ( 
.A(n_134),
.B(n_126),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_147),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_32),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_11),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_135),
.C(n_132),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_12),
.B1(n_14),
.B2(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_159),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_155),
.A2(n_156),
.B1(n_153),
.B2(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_144),
.B(n_146),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_157),
.B1(n_156),
.B2(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_163),
.A2(n_164),
.B1(n_157),
.B2(n_162),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_147),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_50),
.B1(n_16),
.B2(n_17),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_15),
.C(n_24),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_25),
.C(n_31),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_171),
.A2(n_36),
.B(n_37),
.Y(n_172)
);

AOI21x1_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_38),
.B(n_40),
.Y(n_173)
);

OAI21x1_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_41),
.B(n_45),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_46),
.C(n_47),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_48),
.B(n_49),
.Y(n_176)
);


endmodule