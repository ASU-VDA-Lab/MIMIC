module fake_netlist_6_682_n_155 (n_16, n_1, n_34, n_9, n_8, n_18, n_10, n_21, n_24, n_37, n_6, n_15, n_33, n_27, n_3, n_14, n_38, n_0, n_39, n_32, n_4, n_36, n_22, n_26, n_13, n_35, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_40, n_155);

input n_16;
input n_1;
input n_34;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_37;
input n_6;
input n_15;
input n_33;
input n_27;
input n_3;
input n_14;
input n_38;
input n_0;
input n_39;
input n_32;
input n_4;
input n_36;
input n_22;
input n_26;
input n_13;
input n_35;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;
input n_40;

output n_155;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_77;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_82;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_108;
wire n_97;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g65 ( 
.A(n_12),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_0),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_1),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVxp67_ASAP7_75t_SL g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_2),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_5),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_53),
.B(n_65),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_46),
.B1(n_52),
.B2(n_45),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_63),
.B(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_61),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_82),
.C(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_86),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_60),
.B(n_56),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_54),
.B(n_52),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_46),
.B(n_27),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_73),
.B(n_6),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_7),
.B(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_86),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_68),
.B(n_82),
.C(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_87),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_76),
.B(n_69),
.C(n_85),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_72),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_71),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_91),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OA211x2_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_85),
.B(n_109),
.C(n_108),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_115),
.A2(n_85),
.B1(n_108),
.B2(n_106),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_107),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_109),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_105),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_120),
.B(n_118),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_97),
.Y(n_131)
);

NAND4xp25_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_76),
.C(n_96),
.D(n_105),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_106),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_119),
.Y(n_134)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_129),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

OAI33xp33_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_7),
.A3(n_114),
.B1(n_106),
.B2(n_88),
.B3(n_20),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_130),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_138),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_137),
.Y(n_146)
);

AND3x1_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_140),
.C(n_125),
.Y(n_147)
);

NOR3x1_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_124),
.C(n_140),
.Y(n_148)
);

AND4x1_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_125),
.C(n_139),
.D(n_131),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_147),
.Y(n_151)
);

OAI322xp33_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_148),
.A3(n_126),
.B1(n_149),
.B2(n_137),
.C1(n_114),
.C2(n_32),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_126),
.B(n_114),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_16),
.B(n_18),
.Y(n_154)
);

AOI221xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_19),
.B1(n_29),
.B2(n_31),
.C(n_33),
.Y(n_155)
);


endmodule