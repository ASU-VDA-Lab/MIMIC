module fake_jpeg_16535_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_2),
.B(n_1),
.Y(n_7)
);

BUFx2_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_SL g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_22),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g16 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_16),
.A2(n_19),
.B1(n_9),
.B2(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_7),
.B(n_0),
.Y(n_18)
);

OAI21xp33_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_20),
.B(n_21),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_7),
.B(n_3),
.Y(n_21)
);

OR2x2_ASAP7_75t_SL g22 ( 
.A(n_10),
.B(n_9),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_25),
.B1(n_9),
.B2(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_19),
.B1(n_12),
.B2(n_15),
.Y(n_25)
);

AOI22x1_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_20),
.B(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_10),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_14),
.C(n_11),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_33),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_34),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_12),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_5),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_8),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_27),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_37),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.C(n_41),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_31),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_26),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_40),
.B(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_44),
.Y(n_46)
);


endmodule