module real_jpeg_7276_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_167;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_1),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_1),
.A2(n_57),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_1),
.A2(n_57),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_1),
.B(n_44),
.C(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_1),
.A2(n_57),
.B1(n_146),
.B2(n_149),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_1),
.A2(n_181),
.B(n_184),
.C(n_187),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_1),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_1),
.B(n_114),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_1),
.B(n_215),
.C(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_1),
.B(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_2),
.A2(n_23),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_23),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_2),
.A2(n_23),
.B1(n_149),
.B2(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_5),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_5),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_6),
.Y(n_154)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_6),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_6),
.Y(n_186)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_8),
.Y(n_149)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_8),
.Y(n_153)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_8),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_8),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_9),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_9),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_189),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_188),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_141),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_14),
.B(n_141),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_95),
.C(n_126),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_15),
.A2(n_16),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_61),
.B1(n_62),
.B2(n_94),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_17),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_28),
.B1(n_42),
.B2(n_53),
.Y(n_17)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_18),
.A2(n_28),
.B1(n_42),
.B2(n_53),
.Y(n_165)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_20),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_27),
.Y(n_131)
);

NAND2x1_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_42),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_39),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_42),
.Y(n_226)
);

AOI22x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_46),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_54),
.A2(n_57),
.B(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_70),
.B2(n_93),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_63),
.B(n_93),
.C(n_94),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_65),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_70),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_80),
.B1(n_86),
.B2(n_88),
.Y(n_70)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_71),
.A2(n_80),
.B1(n_88),
.B2(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_79),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_82),
.Y(n_218)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_85),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_93),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_93),
.B(n_204),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_95),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_224)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_95),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_95),
.B(n_175),
.C(n_225),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_95),
.A2(n_126),
.B1(n_227),
.B2(n_240),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_103),
.B1(n_119),
.B2(n_120),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_97),
.B(n_114),
.Y(n_208)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_103),
.B(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_104),
.B(n_121),
.Y(n_207)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_114),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B1(n_111),
.B2(n_113),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_111),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_134),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_127),
.A2(n_128),
.B1(n_134),
.B2(n_135),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_169),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_162),
.B2(n_163),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_150),
.B1(n_158),
.B2(n_161),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_168),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_164),
.A2(n_165),
.B1(n_205),
.B2(n_206),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_164),
.B(n_205),
.C(n_234),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_179),
.B2(n_180),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_175),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_201),
.Y(n_202)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_237),
.B(n_243),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_231),
.B(n_236),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_221),
.B(n_230),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_203),
.B(n_220),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_200),
.B(n_202),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_219),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_219),
.Y(n_229)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_229),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_229),
.Y(n_230)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_233),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_242),
.Y(n_243)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);


endmodule