module fake_jpeg_8989_n_299 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_20),
.B1(n_22),
.B2(n_28),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_65),
.B1(n_21),
.B2(n_31),
.Y(n_93)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_70),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_64),
.Y(n_79)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_22),
.B1(n_20),
.B2(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_67),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_69),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_44),
.B1(n_28),
.B2(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_77),
.B1(n_82),
.B2(n_58),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_44),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_85),
.C(n_31),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_43),
.B1(n_44),
.B2(n_37),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_20),
.B1(n_22),
.B2(n_27),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_89),
.B1(n_90),
.B2(n_21),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_39),
.C(n_35),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_36),
.B1(n_30),
.B2(n_18),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_24),
.B1(n_30),
.B2(n_18),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_39),
.B(n_35),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_24),
.B(n_25),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_45),
.A2(n_17),
.B(n_26),
.C(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_25),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_32),
.B1(n_31),
.B2(n_17),
.Y(n_117)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_99),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_96),
.A2(n_103),
.B1(n_74),
.B2(n_73),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_51),
.B1(n_46),
.B2(n_54),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_63),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_59),
.B1(n_49),
.B2(n_58),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_72),
.B(n_92),
.C(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_70),
.C(n_69),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_72),
.C(n_77),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_111),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_112),
.B1(n_113),
.B2(n_84),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_25),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_30),
.B1(n_61),
.B2(n_64),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_78),
.A2(n_66),
.B1(n_32),
.B2(n_21),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_90),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_118),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_23),
.B1(n_26),
.B2(n_74),
.Y(n_144)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_91),
.B(n_75),
.C(n_93),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_135),
.B1(n_94),
.B2(n_82),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_96),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_106),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_71),
.Y(n_132)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_143),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_86),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_109),
.B(n_100),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_111),
.B1(n_97),
.B2(n_105),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_26),
.C(n_23),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_87),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_145),
.B1(n_83),
.B2(n_48),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_81),
.B1(n_48),
.B2(n_73),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_153),
.B1(n_160),
.B2(n_166),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_123),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_162),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_34),
.B(n_33),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_120),
.B(n_103),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_154),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_55),
.B(n_67),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_145),
.B(n_119),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_34),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_159),
.C(n_168),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_86),
.Y(n_158)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_140),
.B1(n_124),
.B2(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_120),
.B(n_13),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_132),
.B(n_13),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_83),
.B1(n_60),
.B2(n_50),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_34),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_88),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_143),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_114),
.C(n_110),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_121),
.C(n_141),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_154),
.B(n_159),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_131),
.B1(n_123),
.B2(n_133),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_184),
.B1(n_186),
.B2(n_189),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_185),
.C(n_188),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_123),
.B1(n_129),
.B2(n_125),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_139),
.B1(n_144),
.B2(n_88),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_155),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_136),
.C(n_110),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_136),
.B1(n_57),
.B2(n_33),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_136),
.C(n_34),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_197),
.C(n_166),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_171),
.B1(n_149),
.B2(n_164),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_163),
.B1(n_148),
.B2(n_156),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_156),
.B(n_164),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_165),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_34),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_181),
.B1(n_180),
.B2(n_189),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_213),
.B1(n_219),
.B2(n_221),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_211),
.B1(n_217),
.B2(n_218),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_209),
.C(n_176),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_208),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_177),
.A2(n_155),
.B(n_148),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_214),
.B(n_193),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_160),
.B1(n_173),
.B2(n_146),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_167),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_170),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_8),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_190),
.B1(n_196),
.B2(n_198),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_185),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_226),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_228),
.C(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_183),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_234),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_176),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_203),
.A2(n_188),
.B1(n_191),
.B2(n_5),
.Y(n_236)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_2),
.C(n_3),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_212),
.B(n_10),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_219),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_202),
.B(n_213),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_249),
.B(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_247),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_211),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_239),
.A2(n_199),
.B(n_204),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_230),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_254),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_225),
.A2(n_216),
.B1(n_209),
.B2(n_221),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_253),
.A2(n_236),
.B1(n_240),
.B2(n_227),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_237),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_226),
.C(n_223),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_258),
.C(n_261),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_263),
.B1(n_242),
.B2(n_252),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_222),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_265),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_228),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_233),
.B1(n_229),
.B2(n_205),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_264),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_215),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_244),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_SL g285 ( 
.A1(n_268),
.A2(n_273),
.B(n_11),
.C(n_12),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_250),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_241),
.B(n_247),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_243),
.B1(n_214),
.B2(n_244),
.Y(n_274)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_274),
.A2(n_258),
.A3(n_10),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_234),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_277),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_208),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_263),
.B(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_208),
.Y(n_279)
);

NOR4xp25_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_283),
.C(n_284),
.D(n_11),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_285),
.B1(n_12),
.B2(n_14),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_10),
.B(n_15),
.C(n_6),
.D(n_7),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_9),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_280),
.A2(n_272),
.B(n_11),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_290),
.C(n_16),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_289),
.B(n_291),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_282),
.B(n_272),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_14),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_293),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_16),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_294),
.A2(n_16),
.B(n_3),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_294),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_297),
.A2(n_292),
.B(n_295),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_298),
.B(n_5),
.Y(n_299)
);


endmodule