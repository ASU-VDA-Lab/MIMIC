module fake_jpeg_1167_n_469 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_469);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_469;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_21),
.B(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_51),
.B(n_94),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_56),
.Y(n_163)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_30),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_60),
.A2(n_32),
.B(n_33),
.Y(n_164)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_61),
.Y(n_109)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_64),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_14),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_65),
.B(n_82),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx12f_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_74),
.B(n_75),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_14),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_16),
.B(n_14),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_17),
.B(n_12),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_11),
.Y(n_92)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_24),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_105),
.B(n_138),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_23),
.B1(n_48),
.B2(n_18),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_113),
.A2(n_117),
.B1(n_122),
.B2(n_140),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_82),
.A2(n_50),
.B1(n_47),
.B2(n_28),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_64),
.A2(n_28),
.B1(n_38),
.B2(n_24),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_67),
.A2(n_25),
.B1(n_43),
.B2(n_47),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_128),
.A2(n_32),
.B1(n_23),
.B2(n_34),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_130),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_72),
.B(n_37),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_50),
.B1(n_47),
.B2(n_28),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_93),
.A2(n_50),
.B1(n_38),
.B2(n_49),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_149),
.A2(n_150),
.B1(n_33),
.B2(n_78),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_101),
.A2(n_38),
.B1(n_25),
.B2(n_43),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_77),
.B(n_44),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_158),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_80),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_96),
.B(n_48),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_100),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_39),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_165),
.B(n_175),
.Y(n_228)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_107),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_169),
.Y(n_232)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx3_ASAP7_75t_SL g225 ( 
.A(n_170),
.Y(n_225)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

AO22x1_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_68),
.B1(n_69),
.B2(n_85),
.Y(n_172)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_36),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_37),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_178),
.B(n_194),
.Y(n_237)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

BUFx4f_ASAP7_75t_SL g180 ( 
.A(n_157),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_180),
.Y(n_235)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_184),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx4_ASAP7_75t_SL g231 ( 
.A(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_188),
.A2(n_201),
.B1(n_204),
.B2(n_207),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_189),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_241)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_36),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_192),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_99),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_135),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_34),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_206),
.Y(n_246)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_128),
.A2(n_18),
.B1(n_52),
.B2(n_59),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_117),
.A2(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_202),
.A2(n_115),
.B1(n_110),
.B2(n_119),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_122),
.A2(n_19),
.B1(n_39),
.B2(n_46),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_121),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_121),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_118),
.B(n_19),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_146),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_212),
.B1(n_127),
.B2(n_124),
.Y(n_245)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_220),
.B1(n_223),
.B2(n_110),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_200),
.A2(n_150),
.B1(n_149),
.B2(n_140),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_218),
.A2(n_226),
.B1(n_243),
.B2(n_249),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_155),
.B1(n_148),
.B2(n_123),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_155),
.B1(n_151),
.B2(n_148),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_192),
.A2(n_151),
.B1(n_70),
.B2(n_71),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_175),
.A2(n_147),
.B1(n_127),
.B2(n_124),
.Y(n_243)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

AOI32xp33_ASAP7_75t_L g247 ( 
.A1(n_166),
.A2(n_160),
.A3(n_119),
.B1(n_156),
.B2(n_134),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_203),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_192),
.A2(n_147),
.B1(n_126),
.B2(n_139),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_191),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_251),
.B(n_258),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_199),
.C(n_165),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_274),
.C(n_263),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_215),
.A2(n_202),
.B1(n_207),
.B2(n_172),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_254),
.A2(n_262),
.B1(n_271),
.B2(n_276),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_255),
.A2(n_229),
.B(n_219),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_215),
.A2(n_172),
.B1(n_184),
.B2(n_190),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_256),
.A2(n_261),
.B1(n_265),
.B2(n_214),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_173),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_260),
.A2(n_236),
.B1(n_233),
.B2(n_221),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_174),
.B1(n_179),
.B2(n_181),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_244),
.A2(n_185),
.B1(n_208),
.B2(n_209),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_211),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_266),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_246),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_268),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_238),
.A2(n_183),
.B1(n_196),
.B2(n_197),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_180),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_246),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_180),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_270),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_171),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_217),
.A2(n_220),
.B1(n_241),
.B2(n_218),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_227),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_170),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_213),
.B(n_109),
.C(n_193),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_212),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_275),
.B(n_277),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_247),
.A2(n_210),
.B1(n_129),
.B2(n_109),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_242),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_278),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_213),
.B(n_186),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_225),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_255),
.A2(n_235),
.B(n_230),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_280),
.A2(n_293),
.B(n_137),
.Y(n_327)
);

NAND3xp33_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_289),
.C(n_274),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g286 ( 
.A(n_253),
.B(n_226),
.CI(n_242),
.CON(n_286),
.SN(n_286)
);

MAJIxp5_ASAP7_75t_SL g324 ( 
.A(n_286),
.B(n_163),
.C(n_239),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_230),
.B1(n_219),
.B2(n_234),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_287),
.A2(n_294),
.B1(n_296),
.B2(n_306),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_156),
.B(n_231),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_231),
.B1(n_222),
.B2(n_240),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_291),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_231),
.B1(n_222),
.B2(n_240),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_225),
.B(n_214),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_297),
.A2(n_304),
.B(n_275),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_278),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_163),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_300),
.A2(n_256),
.B1(n_257),
.B2(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_250),
.A2(n_240),
.B1(n_236),
.B2(n_233),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_260),
.B1(n_257),
.B2(n_262),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_221),
.B(n_198),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_250),
.A2(n_216),
.B1(n_176),
.B2(n_137),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_329),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_308),
.A2(n_311),
.B1(n_315),
.B2(n_320),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

OAI21xp33_ASAP7_75t_SL g348 ( 
.A1(n_310),
.A2(n_327),
.B(n_330),
.Y(n_348)
);

XOR2x2_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_258),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_295),
.C(n_284),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_280),
.A2(n_267),
.B(n_273),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_313),
.A2(n_319),
.B(n_293),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_282),
.A2(n_266),
.B1(n_251),
.B2(n_265),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_292),
.B(n_270),
.Y(n_316)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_316),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_285),
.A2(n_279),
.B1(n_272),
.B2(n_269),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_282),
.A2(n_303),
.B1(n_289),
.B2(n_302),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_287),
.A2(n_259),
.B1(n_277),
.B2(n_252),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_321),
.A2(n_300),
.B1(n_296),
.B2(n_294),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_323),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_332),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_252),
.B1(n_216),
.B2(n_33),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_325),
.A2(n_331),
.B1(n_292),
.B2(n_298),
.Y(n_336)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_328),
.Y(n_358)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_305),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_299),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_333),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_334),
.A2(n_335),
.B1(n_340),
.B2(n_341),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_318),
.A2(n_320),
.B1(n_315),
.B2(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_318),
.A2(n_306),
.B1(n_286),
.B2(n_290),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_330),
.A2(n_286),
.B1(n_298),
.B2(n_297),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_283),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_344),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_283),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_312),
.B(n_291),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_345),
.B(n_328),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_286),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_349),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_311),
.A2(n_284),
.B1(n_112),
.B2(n_46),
.Y(n_351)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_310),
.A2(n_313),
.B(n_327),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_354),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_324),
.B(n_239),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_355),
.B(n_357),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_94),
.Y(n_357)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_337),
.Y(n_361)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_352),
.Y(n_362)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_364),
.Y(n_400)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_356),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_365),
.B(n_366),
.Y(n_386)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_358),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_347),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_367),
.B(n_371),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_354),
.A2(n_319),
.B1(n_321),
.B2(n_326),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_369),
.A2(n_372),
.B1(n_350),
.B2(n_355),
.Y(n_389)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_342),
.A2(n_326),
.B1(n_329),
.B2(n_323),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_377),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_345),
.B(n_325),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_353),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_378),
.B(n_379),
.Y(n_385)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_308),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_380),
.B(n_340),
.Y(n_383)
);

XNOR2x1_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_349),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_338),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_394),
.Y(n_404)
);

OAI22x1_ASAP7_75t_L g387 ( 
.A1(n_381),
.A2(n_348),
.B1(n_333),
.B2(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_389),
.A2(n_374),
.B1(n_370),
.B2(n_377),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_360),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_390),
.B(n_10),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_380),
.C(n_375),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_391),
.B(n_393),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_344),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_373),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_338),
.C(n_341),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_376),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_41),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_381),
.B(n_335),
.C(n_357),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_399),
.B(n_401),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_334),
.C(n_112),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_398),
.A2(n_359),
.B(n_374),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_403),
.Y(n_427)
);

AOI211xp5_ASAP7_75t_L g405 ( 
.A1(n_385),
.A2(n_359),
.B(n_369),
.C(n_372),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_405),
.A2(n_406),
.B1(n_412),
.B2(n_413),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_416),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_370),
.Y(n_408)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_409),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_112),
.C(n_41),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_410),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_395),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_SL g414 ( 
.A(n_399),
.B(n_41),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_417),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_10),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_388),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_421),
.B(n_422),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_400),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_392),
.C(n_393),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_426),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_403),
.B(n_383),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_397),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_404),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_401),
.C(n_394),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_8),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_402),
.B(n_384),
.Y(n_430)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_430),
.Y(n_435)
);

O2A1O1Ixp33_ASAP7_75t_SL g432 ( 
.A1(n_427),
.A2(n_402),
.B(n_387),
.C(n_405),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_418),
.B(n_425),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_418),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_410),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_434),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_427),
.A2(n_414),
.B(n_384),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_436),
.A2(n_438),
.B(n_443),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_420),
.A2(n_416),
.B(n_417),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_424),
.A2(n_41),
.B1(n_8),
.B2(n_35),
.Y(n_439)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_439),
.Y(n_451)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_431),
.Y(n_440)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_440),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_442),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_429),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_428),
.C(n_419),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_444),
.A2(n_450),
.B(n_435),
.Y(n_455)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g458 ( 
.A1(n_446),
.A2(n_8),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_447),
.B(n_448),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_41),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_433),
.B(n_41),
.C(n_1),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_445),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_444),
.A2(n_437),
.B(n_436),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_456),
.A2(n_457),
.B(n_458),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_449),
.A2(n_432),
.B(n_439),
.Y(n_457)
);

AOI321xp33_ASAP7_75t_SL g459 ( 
.A1(n_445),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_459),
.B(n_452),
.Y(n_461)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_460),
.Y(n_465)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_461),
.A2(n_463),
.B(n_451),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_453),
.Y(n_463)
);

OAI211xp5_ASAP7_75t_L g466 ( 
.A1(n_464),
.A2(n_462),
.B(n_450),
.C(n_3),
.Y(n_466)
);

OAI321xp33_ASAP7_75t_L g467 ( 
.A1(n_466),
.A2(n_1),
.A3(n_2),
.B1(n_6),
.B2(n_465),
.C(n_458),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_467),
.A2(n_2),
.B(n_6),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_468),
.Y(n_469)
);


endmodule