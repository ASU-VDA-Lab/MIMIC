module fake_jpeg_29471_n_537 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_537);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_537;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_20),
.B(n_9),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_55),
.B(n_58),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_57),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_8),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_59),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_81),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_10),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_63),
.B(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_23),
.B(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_30),
.B(n_7),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_82),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_92),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_88),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_90),
.Y(n_148)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_102),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_30),
.B(n_7),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_41),
.B(n_27),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_105),
.Y(n_156)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_7),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_77),
.A2(n_27),
.B1(n_31),
.B2(n_36),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_110),
.A2(n_133),
.B1(n_144),
.B2(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_18),
.C(n_46),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_114),
.B(n_158),
.C(n_40),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_105),
.A2(n_41),
.B1(n_36),
.B2(n_52),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_121),
.B(n_143),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_17),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_129),
.B(n_155),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_56),
.A2(n_61),
.B1(n_69),
.B2(n_68),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_59),
.A2(n_43),
.B(n_25),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_90),
.A2(n_36),
.B1(n_46),
.B2(n_51),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_51),
.B1(n_22),
.B2(n_43),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_57),
.A2(n_25),
.B1(n_43),
.B2(n_22),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_153),
.A2(n_162),
.B1(n_49),
.B2(n_76),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_65),
.A2(n_37),
.B1(n_52),
.B2(n_17),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_98),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_67),
.B(n_34),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_24),
.C(n_49),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_59),
.B(n_37),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_161),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_60),
.B(n_38),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_70),
.A2(n_34),
.B1(n_38),
.B2(n_32),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_60),
.B(n_32),
.Y(n_165)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_127),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_168),
.B(n_176),
.Y(n_227)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_45),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_171),
.B(n_175),
.Y(n_251)
);

INVx4_ASAP7_75t_SL g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_172),
.Y(n_246)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_174),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_113),
.B(n_45),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_116),
.Y(n_176)
);

BUFx2_ASAP7_75t_SL g177 ( 
.A(n_142),
.Y(n_177)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_177),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_119),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_178),
.Y(n_238)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_180),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_181),
.B(n_182),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_111),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_142),
.A2(n_54),
.B1(n_71),
.B2(n_73),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_183),
.A2(n_193),
.B1(n_218),
.B2(n_53),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_116),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_184),
.B(n_185),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_136),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_186),
.B(n_95),
.Y(n_230)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_187),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_188),
.Y(n_242)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_121),
.B(n_104),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_189),
.B(n_94),
.CI(n_95),
.CON(n_228),
.SN(n_228)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_40),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_192),
.B(n_198),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_25),
.B1(n_24),
.B2(n_48),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_196),
.A2(n_108),
.B1(n_141),
.B2(n_128),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_125),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_197),
.B(n_200),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_114),
.B(n_48),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_112),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_126),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_204),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_110),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_210),
.Y(n_239)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_107),
.Y(n_207)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_207),
.Y(n_253)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_149),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_214),
.Y(n_241)
);

BUFx8_ASAP7_75t_L g212 ( 
.A(n_107),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_212),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_122),
.B(n_48),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_215),
.Y(n_257)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_216),
.A2(n_219),
.B1(n_152),
.B2(n_107),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_217),
.A2(n_85),
.B1(n_80),
.B2(n_79),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_109),
.A2(n_49),
.B1(n_22),
.B2(n_21),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_159),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_148),
.C(n_145),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_221),
.B(n_230),
.C(n_196),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_SL g223 ( 
.A(n_208),
.B(n_144),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_223),
.B(n_215),
.C(n_181),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_108),
.B1(n_141),
.B2(n_135),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_224),
.A2(n_250),
.B1(n_178),
.B2(n_159),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_228),
.B(n_249),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_152),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_235),
.B(n_152),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_170),
.A2(n_190),
.B1(n_148),
.B2(n_188),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_247),
.A2(n_219),
.B1(n_214),
.B2(n_209),
.Y(n_291)
);

AO22x1_ASAP7_75t_L g249 ( 
.A1(n_189),
.A2(n_159),
.B1(n_94),
.B2(n_72),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_150),
.B1(n_146),
.B2(n_123),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_171),
.B(n_132),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_175),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_262),
.B(n_266),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_254),
.B(n_192),
.CI(n_186),
.CON(n_263),
.SN(n_263)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_263),
.B(n_268),
.Y(n_329)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_267),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_254),
.B(n_208),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_218),
.B(n_193),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_270),
.A2(n_283),
.B(n_292),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_233),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_271),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_280),
.Y(n_316)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_274),
.A2(n_277),
.B1(n_282),
.B2(n_284),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_249),
.Y(n_275)
);

NAND2x1_ASAP7_75t_SL g306 ( 
.A(n_275),
.B(n_238),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_276),
.A2(n_279),
.B1(n_287),
.B2(n_291),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_223),
.A2(n_150),
.B1(n_146),
.B2(n_139),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_199),
.C(n_213),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_281),
.C(n_242),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_235),
.B1(n_249),
.B2(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_180),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_124),
.B1(n_201),
.B2(n_169),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_221),
.A2(n_178),
.B(n_194),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_228),
.A2(n_210),
.B1(n_140),
.B2(n_135),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_191),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_285),
.B(n_289),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_L g286 ( 
.A1(n_228),
.A2(n_164),
.B1(n_138),
.B2(n_140),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_234),
.B1(n_238),
.B2(n_130),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_128),
.B1(n_130),
.B2(n_167),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_179),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_236),
.Y(n_290)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_242),
.A2(n_205),
.B1(n_147),
.B2(n_172),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_236),
.Y(n_293)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g294 ( 
.A1(n_225),
.A2(n_219),
.B(n_205),
.C(n_174),
.Y(n_294)
);

AOI21xp33_ASAP7_75t_L g328 ( 
.A1(n_294),
.A2(n_256),
.B(n_212),
.Y(n_328)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_231),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_296),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_255),
.B(n_202),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_297),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_227),
.B(n_239),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_300),
.A2(n_317),
.B(n_320),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_281),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_301),
.A2(n_311),
.B(n_313),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_263),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_234),
.B1(n_238),
.B2(n_220),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_304),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_306),
.A2(n_283),
.B(n_288),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_297),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_308),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_309),
.A2(n_291),
.B1(n_276),
.B2(n_292),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_275),
.B(n_234),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_277),
.A2(n_229),
.B1(n_226),
.B2(n_260),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_312),
.A2(n_314),
.B1(n_287),
.B2(n_267),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_269),
.A2(n_222),
.B1(n_220),
.B2(n_243),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_284),
.A2(n_229),
.B1(n_226),
.B2(n_248),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_298),
.A2(n_245),
.B(n_261),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_298),
.A2(n_245),
.B1(n_253),
.B2(n_237),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_261),
.B(n_195),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_322),
.A2(n_212),
.B(n_207),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_279),
.A2(n_78),
.B1(n_89),
.B2(n_87),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_324),
.A2(n_282),
.B1(n_274),
.B2(n_289),
.Y(n_345)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_268),
.A2(n_260),
.A3(n_248),
.B1(n_243),
.B2(n_237),
.Y(n_327)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_328),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_280),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_262),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_334),
.B(n_367),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_328),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_335),
.B(n_355),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_336),
.A2(n_340),
.B1(n_358),
.B2(n_299),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_338),
.A2(n_362),
.B(n_363),
.Y(n_369)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_305),
.Y(n_339)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_339),
.Y(n_372)
);

INVx8_ASAP7_75t_L g342 ( 
.A(n_310),
.Y(n_342)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_263),
.C(n_272),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_344),
.B(n_348),
.C(n_350),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_345),
.A2(n_360),
.B1(n_346),
.B2(n_343),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_318),
.A2(n_270),
.B1(n_285),
.B2(n_281),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_346),
.A2(n_354),
.B1(n_359),
.B2(n_360),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_347),
.B(n_311),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_278),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_302),
.B(n_266),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_308),
.B(n_265),
.Y(n_351)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_325),
.B(n_271),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_353),
.B(n_365),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_318),
.A2(n_324),
.B1(n_330),
.B2(n_333),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g355 ( 
.A(n_302),
.B(n_294),
.CI(n_293),
.CON(n_355),
.SN(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_294),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_361),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_303),
.A2(n_264),
.B1(n_273),
.B2(n_296),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_333),
.A2(n_264),
.B1(n_290),
.B2(n_253),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_303),
.A2(n_244),
.B1(n_256),
.B2(n_84),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_187),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_317),
.A2(n_173),
.B(n_244),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_323),
.A2(n_53),
.B1(n_1),
.B2(n_2),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_364),
.A2(n_366),
.B1(n_341),
.B2(n_339),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_310),
.B(n_12),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_323),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_3),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_349),
.A2(n_320),
.B(n_322),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_371),
.A2(n_6),
.B(n_11),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_300),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_375),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_374),
.A2(n_378),
.B1(n_398),
.B2(n_357),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_301),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_351),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_376),
.B(n_389),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_337),
.A2(n_315),
.B1(n_306),
.B2(n_319),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_301),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_387),
.Y(n_412)
);

NOR2x1_ASAP7_75t_L g382 ( 
.A(n_356),
.B(n_314),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_382),
.B(n_385),
.Y(n_407)
);

OAI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_337),
.A2(n_309),
.B1(n_327),
.B2(n_306),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_383),
.A2(n_386),
.B1(n_400),
.B2(n_307),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_354),
.A2(n_312),
.B1(n_313),
.B2(n_315),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_342),
.Y(n_388)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_388),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_341),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_359),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_390),
.Y(n_401)
);

AOI22x1_ASAP7_75t_L g392 ( 
.A1(n_349),
.A2(n_311),
.B1(n_299),
.B2(n_305),
.Y(n_392)
);

OA22x2_ASAP7_75t_L g413 ( 
.A1(n_392),
.A2(n_331),
.B1(n_326),
.B2(n_307),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_311),
.Y(n_393)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_393),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_366),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_394),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_361),
.B(n_311),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_21),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_352),
.A2(n_304),
.B(n_321),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_396),
.A2(n_362),
.B(n_355),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_358),
.A2(n_343),
.B1(n_340),
.B2(n_338),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_321),
.Y(n_399)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_399),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_352),
.B(n_357),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_402),
.A2(n_411),
.B(n_416),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_403),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g446 ( 
.A(n_404),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_386),
.A2(n_355),
.B1(n_345),
.B2(n_332),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_408),
.A2(n_415),
.B1(n_378),
.B2(n_371),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_350),
.C(n_332),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_397),
.C(n_373),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_369),
.A2(n_331),
.B(n_364),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_413),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_396),
.A2(n_326),
.B(n_13),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_385),
.B(n_3),
.Y(n_417)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_417),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_422),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_379),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_420),
.B(n_421),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_399),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_392),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_398),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_423),
.A2(n_382),
.B1(n_400),
.B2(n_368),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_381),
.Y(n_424)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_424),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_3),
.Y(n_426)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_426),
.Y(n_431)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_427),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_429),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_441),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_410),
.B(n_380),
.C(n_375),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_440),
.C(n_451),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_387),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_436),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_370),
.C(n_392),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_370),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_391),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_452),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_443),
.A2(n_407),
.B1(n_422),
.B2(n_417),
.Y(n_457)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_409),
.Y(n_444)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_415),
.A2(n_374),
.B1(n_368),
.B2(n_393),
.Y(n_448)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_403),
.A2(n_384),
.B1(n_395),
.B2(n_391),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_449),
.A2(n_453),
.B1(n_429),
.B2(n_425),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_406),
.B(n_21),
.C(n_12),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_11),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_408),
.C(n_407),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_461),
.C(n_465),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_457),
.A2(n_459),
.B1(n_467),
.B2(n_416),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_413),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_460),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_418),
.C(n_404),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_444),
.A2(n_402),
.B(n_440),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_463),
.A2(n_430),
.B(n_453),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_425),
.C(n_401),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_446),
.C(n_436),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_466),
.B(n_469),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_443),
.A2(n_401),
.B1(n_419),
.B2(n_411),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_438),
.Y(n_469)
);

BUFx4f_ASAP7_75t_SL g470 ( 
.A(n_439),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_470),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_450),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_471),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_447),
.B(n_413),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_472),
.B(n_448),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_468),
.A2(n_445),
.B1(n_447),
.B2(n_450),
.Y(n_474)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_474),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_476),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_472),
.A2(n_419),
.B(n_413),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_477),
.Y(n_496)
);

XOR2x1_ASAP7_75t_SL g478 ( 
.A(n_467),
.B(n_460),
.Y(n_478)
);

MAJx2_ASAP7_75t_L g505 ( 
.A(n_478),
.B(n_460),
.C(n_431),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_435),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_483),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_482),
.B(n_488),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_430),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_466),
.A2(n_465),
.B1(n_455),
.B2(n_434),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_490),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_428),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_456),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_454),
.A2(n_437),
.B(n_405),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_458),
.A2(n_437),
.B(n_405),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_489),
.B(n_427),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_462),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_485),
.C(n_456),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_483),
.C(n_479),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_494),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_484),
.B(n_454),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_503),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_505),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_470),
.Y(n_501)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_501),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_473),
.Y(n_502)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_502),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_470),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_431),
.Y(n_504)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_504),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_497),
.A2(n_478),
.B1(n_459),
.B2(n_475),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_514),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_498),
.B(n_481),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_507),
.A2(n_515),
.B(n_493),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_499),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_496),
.A2(n_481),
.B1(n_476),
.B2(n_477),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_492),
.B(n_426),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_491),
.A2(n_487),
.B(n_451),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_516),
.A2(n_510),
.B(n_511),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_SL g527 ( 
.A(n_518),
.B(n_516),
.C(n_515),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g528 ( 
.A(n_520),
.B(n_521),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_SL g522 ( 
.A(n_509),
.B(n_505),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_522),
.A2(n_507),
.B(n_514),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_492),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_523),
.A2(n_524),
.B1(n_517),
.B2(n_500),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_511),
.B(n_500),
.Y(n_524)
);

A2O1A1Ixp33_ASAP7_75t_SL g531 ( 
.A1(n_525),
.A2(n_527),
.B(n_513),
.C(n_423),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_526),
.B(n_519),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_529),
.A2(n_530),
.B(n_531),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_512),
.C(n_506),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_11),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_15),
.B(n_16),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_534),
.A2(n_15),
.B(n_16),
.Y(n_535)
);

AOI221xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_15),
.B1(n_16),
.B2(n_21),
.C(n_389),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_536),
.A2(n_15),
.B(n_16),
.Y(n_537)
);


endmodule