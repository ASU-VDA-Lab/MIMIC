module fake_jpeg_11973_n_99 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_12),
.B(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_2),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_49),
.Y(n_50)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_48),
.B1(n_40),
.B2(n_35),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_37),
.B1(n_39),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_48),
.A2(n_37),
.B1(n_39),
.B2(n_35),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_42),
.B1(n_44),
.B2(n_4),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_47),
.A3(n_46),
.B1(n_41),
.B2(n_49),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_19),
.B(n_6),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_24),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_64),
.Y(n_75)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_44),
.C(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_2),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_17),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_67),
.A2(n_53),
.B1(n_57),
.B2(n_5),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_71),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_76),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_79),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_68),
.Y(n_81)
);

NOR4xp25_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_83),
.C(n_84),
.D(n_8),
.Y(n_86)
);

BUFx24_ASAP7_75t_SL g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_7),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_87),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_69),
.B(n_71),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_82),
.B(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_90),
.B(n_91),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_73),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_92),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_9),
.B(n_10),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_89),
.C(n_70),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_9),
.Y(n_97)
);

OAI221xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.C(n_96),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_13),
.Y(n_99)
);


endmodule