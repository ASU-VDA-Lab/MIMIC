module fake_netlist_5_2278_n_1862 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1862);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1862;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_104),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_78),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_70),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_19),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_87),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_39),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_136),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_103),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_7),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_105),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_64),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_130),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_31),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_1),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_134),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_58),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_55),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_175),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_124),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_155),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_56),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_92),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_149),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_170),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_140),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_157),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_67),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_180),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_43),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_151),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_37),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_70),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_186),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_27),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_41),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_177),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_102),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_59),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_115),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_77),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_23),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_53),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_85),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_46),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_12),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_63),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_90),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_106),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_111),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_69),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_15),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_91),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_86),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_93),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_2),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_55),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_114),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_58),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_179),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_101),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_118),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_165),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_40),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_147),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_36),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_42),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_190),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_25),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_32),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_94),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_46),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_95),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_36),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_108),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_145),
.Y(n_276)
);

BUFx5_ASAP7_75t_L g277 ( 
.A(n_52),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_31),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_167),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_89),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_150),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_159),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_69),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_18),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_139),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_122),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_51),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_97),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_172),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_132),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_5),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_110),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_2),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_79),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_163),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_161),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_82),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_20),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_21),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_142),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_63),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_96),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_27),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_120),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_28),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_171),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_57),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_12),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_181),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_47),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_146),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_73),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_127),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_60),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_81),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_184),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_107),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_4),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_43),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_128),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_168),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_98),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_121),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_11),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_125),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_21),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_34),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_9),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_34),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_113),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_15),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_52),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_62),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_185),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_99),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_18),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_45),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_3),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_72),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_76),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_29),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_35),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_29),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_20),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_148),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_83),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_53),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_23),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_60),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_62),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_26),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_8),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_47),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_26),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_68),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_61),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_154),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_24),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_4),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_71),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_75),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_143),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_152),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_153),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_30),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_45),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_1),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_123),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_9),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_7),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_3),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_33),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_6),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_49),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_10),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_13),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_88),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_32),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_80),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_24),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_25),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_277),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_277),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_277),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_232),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_225),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_215),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_237),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_277),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_277),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_286),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_277),
.Y(n_394)
);

INVxp33_ASAP7_75t_SL g395 ( 
.A(n_194),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_204),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_277),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_277),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_300),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_257),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_318),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_216),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_300),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_300),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_220),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_300),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_194),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_369),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_326),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_221),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_204),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_222),
.Y(n_412)
);

BUFx6f_ASAP7_75t_SL g413 ( 
.A(n_204),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_300),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_300),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_203),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_340),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_364),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_300),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_231),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_300),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_223),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_214),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_214),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_366),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_214),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_366),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_206),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_366),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_293),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_231),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_231),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_214),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_214),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_251),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_251),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_242),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_224),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_332),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_251),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_253),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_230),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_233),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_251),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_251),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_234),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_236),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_206),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_284),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_252),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_239),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_284),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_240),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_284),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_284),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_284),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_253),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_241),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_382),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_250),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_196),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_196),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_234),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_245),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_255),
.Y(n_469)
);

INVxp33_ASAP7_75t_SL g470 ( 
.A(n_209),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_260),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_261),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_253),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_262),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_246),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_246),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_207),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_264),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_263),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_264),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_285),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_481),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_425),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_481),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_423),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_423),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_424),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_408),
.A2(n_209),
.B1(n_371),
.B2(n_212),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_389),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

NAND2xp33_ASAP7_75t_L g491 ( 
.A(n_383),
.B(n_212),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_481),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_386),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_384),
.A2(n_280),
.B(n_198),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_481),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_426),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_481),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_436),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_426),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_436),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_387),
.A2(n_372),
.B1(n_374),
.B2(n_371),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_433),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_434),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_427),
.B(n_199),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_443),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_439),
.A2(n_210),
.B1(n_283),
.B2(n_272),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_402),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_447),
.B(n_400),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_434),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_405),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_443),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_390),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_384),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_410),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_385),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_435),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_407),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_412),
.B(n_228),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_395),
.A2(n_342),
.B1(n_353),
.B2(n_352),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_422),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_385),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_447),
.B(n_199),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_420),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_438),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_440),
.B(n_228),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_463),
.B(n_305),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_442),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_391),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_444),
.B(n_305),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_435),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_391),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_441),
.A2(n_374),
.B1(n_375),
.B2(n_372),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_470),
.A2(n_357),
.B1(n_360),
.B2(n_375),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_445),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_445),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_452),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_388),
.B(n_298),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_446),
.Y(n_541)
);

AND2x2_ASAP7_75t_SL g542 ( 
.A(n_441),
.B(n_198),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_446),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_450),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_450),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_453),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_454),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_453),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_458),
.B(n_294),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_455),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_393),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_471),
.B(n_474),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_416),
.B(n_328),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_455),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_437),
.B(n_328),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_479),
.B(n_280),
.Y(n_557)
);

NOR2x1_ASAP7_75t_L g558 ( 
.A(n_456),
.B(n_363),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_449),
.B(n_348),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_456),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_457),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_396),
.B(n_191),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_482),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_542),
.B(n_458),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_515),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_510),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_483),
.B(n_363),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_L g568 ( 
.A(n_483),
.B(n_394),
.C(n_392),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_542),
.B(n_430),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_517),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_482),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_520),
.B(n_448),
.Y(n_572)
);

INVxp33_ASAP7_75t_L g573 ( 
.A(n_519),
.Y(n_573)
);

AND3x2_ASAP7_75t_L g574 ( 
.A(n_550),
.B(n_269),
.C(n_267),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_517),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_482),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_527),
.B(n_459),
.Y(n_577)
);

BUFx6f_ASAP7_75t_SL g578 ( 
.A(n_527),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_514),
.Y(n_579)
);

INVx5_ASAP7_75t_L g580 ( 
.A(n_515),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_510),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_559),
.B(n_432),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_531),
.B(n_462),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_493),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_493),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_524),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_506),
.B(n_429),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_493),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_523),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_523),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_523),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_550),
.B(n_464),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_SL g594 ( 
.A1(n_506),
.A2(n_348),
.B(n_392),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_530),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_530),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_530),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_482),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_533),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_494),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_533),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_494),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_494),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_533),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_515),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_515),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_485),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_553),
.A2(n_472),
.B1(n_469),
.B2(n_227),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_499),
.Y(n_611)
);

INVx1_ASAP7_75t_SL g612 ( 
.A(n_552),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_482),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_554),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_485),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_495),
.A2(n_397),
.B(n_394),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_549),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_486),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_486),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_487),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_554),
.B(n_429),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_546),
.A2(n_229),
.B1(n_235),
.B2(n_219),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_495),
.Y(n_624)
);

BUFx6f_ASAP7_75t_SL g625 ( 
.A(n_527),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_528),
.B(n_459),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_487),
.Y(n_627)
);

INVx8_ASAP7_75t_L g628 ( 
.A(n_528),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_490),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_499),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_492),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_513),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_490),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_528),
.B(n_460),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_557),
.B(n_396),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_524),
.Y(n_636)
);

BUFx4f_ASAP7_75t_L g637 ( 
.A(n_549),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_549),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_559),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_528),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_562),
.B(n_411),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_549),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_497),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_513),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_513),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_507),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_507),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_556),
.B(n_465),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_556),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_507),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_497),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_535),
.A2(n_379),
.B1(n_381),
.B2(n_377),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_507),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_500),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_500),
.B(n_503),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_525),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_503),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_540),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_539),
.B(n_211),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_504),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_489),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_492),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_509),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_504),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_505),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_505),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_492),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_511),
.B(n_480),
.Y(n_668)
);

INVxp33_ASAP7_75t_L g669 ( 
.A(n_502),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_512),
.B(n_411),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_511),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_518),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_501),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_491),
.A2(n_267),
.B1(n_270),
.B2(n_269),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_484),
.B(n_460),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_488),
.A2(n_270),
.B1(n_339),
.B2(n_274),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_516),
.B(n_473),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_484),
.B(n_461),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_532),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_522),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_532),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_540),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_536),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_536),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_484),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_484),
.B(n_461),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_537),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_537),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_498),
.B(n_397),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_SL g690 ( 
.A1(n_534),
.A2(n_413),
.B1(n_473),
.B2(n_401),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_492),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_501),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_558),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_526),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_541),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_541),
.Y(n_696)
);

BUFx4f_ASAP7_75t_L g697 ( 
.A(n_549),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_543),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_543),
.B(n_480),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_492),
.Y(n_700)
);

INVxp33_ASAP7_75t_L g701 ( 
.A(n_508),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_544),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_498),
.B(n_398),
.Y(n_703)
);

OAI22x1_ASAP7_75t_L g704 ( 
.A1(n_535),
.A2(n_521),
.B1(n_508),
.B2(n_379),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_498),
.B(n_544),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_558),
.A2(n_339),
.B1(n_304),
.B2(n_306),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_545),
.B(n_217),
.Y(n_707)
);

BUFx10_ASAP7_75t_L g708 ( 
.A(n_529),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_501),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_501),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_640),
.B(n_538),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_640),
.A2(n_548),
.B1(n_409),
.B2(n_418),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_693),
.B(n_545),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_693),
.B(n_547),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_587),
.B(n_285),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_628),
.B(n_547),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_614),
.B(n_521),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_647),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_582),
.B(n_451),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_594),
.A2(n_309),
.B(n_311),
.C(n_256),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_647),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_565),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_628),
.B(n_551),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_668),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_628),
.B(n_207),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_653),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_628),
.B(n_551),
.Y(n_727)
);

BUFx12f_ASAP7_75t_L g728 ( 
.A(n_708),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_628),
.B(n_555),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_653),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_669),
.A2(n_344),
.B1(n_345),
.B2(n_338),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_588),
.B(n_555),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_587),
.B(n_285),
.Y(n_733)
);

NAND3xp33_ASAP7_75t_L g734 ( 
.A(n_594),
.B(n_243),
.C(n_238),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_588),
.B(n_561),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_635),
.B(n_636),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_668),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_636),
.B(n_285),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_649),
.B(n_561),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_649),
.B(n_498),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_585),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_656),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_648),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_577),
.B(n_560),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_654),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_639),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_657),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_657),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_699),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_626),
.B(n_634),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_639),
.B(n_192),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_585),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_699),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_655),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_609),
.B(n_615),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_578),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_566),
.B(n_192),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_566),
.B(n_582),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_564),
.B(n_193),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_655),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_615),
.B(n_560),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_648),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_618),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_586),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_618),
.B(n_560),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_619),
.B(n_560),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_619),
.Y(n_767)
);

INVxp33_ASAP7_75t_L g768 ( 
.A(n_622),
.Y(n_768)
);

OAI221xp5_ASAP7_75t_L g769 ( 
.A1(n_674),
.A2(n_351),
.B1(n_367),
.B2(n_373),
.C(n_376),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_586),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_578),
.A2(n_417),
.B1(n_291),
.B2(n_301),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_567),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_581),
.B(n_193),
.Y(n_773)
);

INVx8_ASAP7_75t_L g774 ( 
.A(n_578),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_568),
.B(n_285),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_568),
.B(n_322),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_625),
.A2(n_271),
.B1(n_268),
.B2(n_275),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_567),
.A2(n_377),
.B1(n_381),
.B2(n_299),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_567),
.A2(n_319),
.B1(n_292),
.B2(n_287),
.Y(n_779)
);

BUFx5_ASAP7_75t_L g780 ( 
.A(n_624),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_574),
.Y(n_781)
);

BUFx8_ASAP7_75t_L g782 ( 
.A(n_656),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_620),
.B(n_627),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_660),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_589),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_565),
.B(n_322),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_567),
.B(n_465),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_627),
.Y(n_788)
);

OAI221xp5_ASAP7_75t_L g789 ( 
.A1(n_676),
.A2(n_258),
.B1(n_289),
.B2(n_288),
.C(n_279),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_664),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_629),
.B(n_560),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_629),
.B(n_633),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_633),
.B(n_501),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_643),
.B(n_501),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_643),
.B(n_218),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_589),
.Y(n_796)
);

O2A1O1Ixp5_ASAP7_75t_L g797 ( 
.A1(n_616),
.A2(n_317),
.B(n_248),
.C(n_249),
.Y(n_797)
);

INVx8_ASAP7_75t_L g798 ( 
.A(n_625),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_651),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_565),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_658),
.B(n_247),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_682),
.B(n_623),
.Y(n_802)
);

XOR2xp5_ASAP7_75t_L g803 ( 
.A(n_579),
.B(n_276),
.Y(n_803)
);

CKINVDCx16_ASAP7_75t_R g804 ( 
.A(n_708),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_708),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_651),
.B(n_226),
.Y(n_806)
);

AO22x2_ASAP7_75t_L g807 ( 
.A1(n_593),
.A2(n_254),
.B1(n_244),
.B2(n_265),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_665),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_665),
.B(n_273),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_573),
.B(n_466),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_606),
.B(n_207),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_572),
.B(n_195),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_606),
.B(n_322),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_SL g814 ( 
.A(n_625),
.B(n_413),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_600),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_584),
.A2(n_331),
.B1(n_290),
.B2(n_282),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_608),
.B(n_322),
.Y(n_817)
);

OAI22xp33_ASAP7_75t_L g818 ( 
.A1(n_701),
.A2(n_334),
.B1(n_278),
.B2(n_266),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_664),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_612),
.B(n_259),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_641),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_666),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_679),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_624),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_624),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_608),
.B(n_322),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_708),
.Y(n_827)
);

INVx8_ASAP7_75t_L g828 ( 
.A(n_659),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_569),
.A2(n_336),
.B1(n_281),
.B2(n_296),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_666),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_679),
.B(n_207),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_681),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_671),
.B(n_295),
.Y(n_833)
);

INVx8_ASAP7_75t_L g834 ( 
.A(n_659),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_704),
.A2(n_419),
.B1(n_403),
.B2(n_404),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_SL g836 ( 
.A(n_661),
.B(n_413),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_672),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_672),
.B(n_307),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_704),
.A2(n_421),
.B1(n_403),
.B2(n_404),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_707),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_600),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_683),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_659),
.A2(n_314),
.B1(n_358),
.B2(n_346),
.Y(n_843)
);

NAND2x1p5_ASAP7_75t_L g844 ( 
.A(n_683),
.B(n_310),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_681),
.B(n_207),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_602),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_607),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_688),
.B(n_313),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_688),
.B(n_316),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_695),
.B(n_341),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_684),
.B(n_207),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_602),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_659),
.A2(n_361),
.B1(n_197),
.B2(n_200),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_610),
.B(n_333),
.C(n_329),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_696),
.B(n_399),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_670),
.B(n_195),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_659),
.A2(n_347),
.B1(n_297),
.B2(n_303),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_702),
.B(n_399),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_702),
.B(n_406),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_685),
.B(n_406),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_684),
.B(n_207),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_677),
.B(n_197),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_687),
.B(n_207),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_687),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_698),
.B(n_414),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_698),
.B(n_312),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_R g867 ( 
.A(n_804),
.B(n_663),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_825),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_728),
.Y(n_869)
);

BUFx4f_ASAP7_75t_SL g870 ( 
.A(n_805),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_736),
.B(n_570),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_R g872 ( 
.A(n_814),
.B(n_680),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_742),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_812),
.B(n_570),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_743),
.B(n_707),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_768),
.B(n_694),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_746),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_745),
.Y(n_878)
);

INVx5_ASAP7_75t_L g879 ( 
.A(n_825),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_L g880 ( 
.A(n_712),
.B(n_652),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_756),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_768),
.B(n_690),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_747),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_747),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_722),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_748),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_810),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_805),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_762),
.B(n_707),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_784),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_784),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_746),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_756),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_722),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_790),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_790),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_756),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_759),
.A2(n_707),
.B1(n_705),
.B2(n_575),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_819),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_754),
.B(n_707),
.Y(n_900)
);

O2A1O1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_731),
.A2(n_689),
.B(n_703),
.C(n_595),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_827),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_763),
.B(n_575),
.Y(n_903)
);

INVx3_ASAP7_75t_SL g904 ( 
.A(n_774),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_SL g905 ( 
.A(n_854),
.B(n_652),
.C(n_308),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_767),
.B(n_583),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_780),
.B(n_580),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_819),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_788),
.B(n_799),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_758),
.B(n_590),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_825),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_825),
.B(n_617),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_827),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_760),
.A2(n_706),
.B1(n_596),
.B2(n_597),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_823),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_780),
.B(n_580),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_808),
.B(n_822),
.Y(n_917)
);

OAI22xp5_ASAP7_75t_SL g918 ( 
.A1(n_803),
.A2(n_350),
.B1(n_302),
.B2(n_315),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_823),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_780),
.B(n_580),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_832),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_830),
.B(n_590),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_782),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_797),
.A2(n_616),
.B(n_592),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_750),
.A2(n_592),
.B(n_591),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_724),
.B(n_673),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_832),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_758),
.B(n_591),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_847),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_737),
.B(n_673),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_824),
.B(n_617),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_864),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_716),
.A2(n_697),
.B(n_637),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_837),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_741),
.Y(n_935)
);

INVx4_ASAP7_75t_SL g936 ( 
.A(n_847),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_807),
.A2(n_601),
.B1(n_605),
.B2(n_599),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_847),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_717),
.B(n_595),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_719),
.B(n_320),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_772),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_780),
.B(n_580),
.Y(n_942)
);

AOI22x1_ASAP7_75t_L g943 ( 
.A1(n_800),
.A2(n_710),
.B1(n_709),
.B2(n_673),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_802),
.B(n_599),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_782),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_774),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_847),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_774),
.Y(n_948)
);

AND2x6_ASAP7_75t_L g949 ( 
.A(n_824),
.B(n_692),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_798),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_798),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_752),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_798),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_842),
.B(n_605),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_807),
.A2(n_603),
.B1(n_414),
.B2(n_415),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_749),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_764),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_755),
.B(n_603),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_753),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_783),
.B(n_563),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_792),
.B(n_713),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_787),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_714),
.B(n_563),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_711),
.B(n_692),
.Y(n_964)
);

INVx5_ASAP7_75t_L g965 ( 
.A(n_787),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_781),
.B(n_692),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_772),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_779),
.B(n_709),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_828),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_740),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_770),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_779),
.B(n_709),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_732),
.B(n_735),
.Y(n_973)
);

NAND3xp33_ASAP7_75t_SL g974 ( 
.A(n_843),
.B(n_327),
.C(n_325),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_773),
.B(n_821),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_785),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_718),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_793),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_796),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_815),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_739),
.B(n_563),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_771),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_828),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_794),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_840),
.B(n_734),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_757),
.B(n_751),
.Y(n_986)
);

NOR2xp67_ASAP7_75t_L g987 ( 
.A(n_773),
.B(n_675),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_820),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_721),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_757),
.B(n_563),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_816),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_828),
.Y(n_992)
);

OR2x6_ASAP7_75t_L g993 ( 
.A(n_834),
.B(n_840),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_751),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_731),
.A2(n_678),
.B(n_686),
.C(n_630),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_834),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_726),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_841),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_834),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_730),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_846),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_835),
.B(n_571),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_835),
.B(n_571),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_844),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_852),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_801),
.Y(n_1006)
);

INVx8_ASAP7_75t_L g1007 ( 
.A(n_836),
.Y(n_1007)
);

NOR2x1p5_ASAP7_75t_L g1008 ( 
.A(n_795),
.B(n_337),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_807),
.A2(n_415),
.B1(n_421),
.B2(n_419),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_839),
.B(n_571),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_778),
.B(n_343),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_778),
.B(n_349),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_839),
.B(n_571),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_761),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_844),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_765),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_R g1017 ( 
.A(n_856),
.B(n_200),
.Y(n_1017)
);

NAND3xp33_ASAP7_75t_SL g1018 ( 
.A(n_857),
.B(n_356),
.C(n_354),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_856),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_860),
.B(n_576),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_806),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_L g1022 ( 
.A(n_723),
.B(n_607),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_866),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_766),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_791),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_865),
.Y(n_1026)
);

OR2x6_ASAP7_75t_L g1027 ( 
.A(n_720),
.B(n_468),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_855),
.B(n_637),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_858),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_866),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_862),
.B(n_468),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_775),
.A2(n_776),
.B1(n_789),
.B2(n_769),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_727),
.A2(n_697),
.B(n_617),
.Y(n_1033)
);

CKINVDCx6p67_ASAP7_75t_R g1034 ( 
.A(n_809),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_744),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_729),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_831),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_818),
.B(n_355),
.Y(n_1038)
);

NOR2x1_ASAP7_75t_L g1039 ( 
.A(n_946),
.B(n_833),
.Y(n_1039)
);

CKINVDCx11_ASAP7_75t_R g1040 ( 
.A(n_923),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_877),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_L g1042 ( 
.A(n_905),
.B(n_862),
.C(n_818),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_873),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_884),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_934),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_986),
.A2(n_853),
.B(n_738),
.C(n_715),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_892),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_868),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_884),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1022),
.A2(n_725),
.B(n_697),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_975),
.B(n_777),
.Y(n_1051)
);

CKINVDCx20_ASAP7_75t_R g1052 ( 
.A(n_867),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1019),
.A2(n_849),
.B1(n_848),
.B2(n_838),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_887),
.B(n_829),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_973),
.A2(n_642),
.B(n_617),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_878),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_975),
.A2(n_850),
.B(n_738),
.C(n_733),
.Y(n_1057)
);

NOR2xp67_ASAP7_75t_SL g1058 ( 
.A(n_879),
.B(n_965),
.Y(n_1058)
);

OAI221xp5_ASAP7_75t_L g1059 ( 
.A1(n_1038),
.A2(n_359),
.B1(n_370),
.B2(n_368),
.C(n_859),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_994),
.B(n_715),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_940),
.B(n_733),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_939),
.B(n_786),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_867),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_883),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_891),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_939),
.B(n_786),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_961),
.A2(n_638),
.B(n_642),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1032),
.A2(n_863),
.B1(n_861),
.B2(n_851),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1032),
.A2(n_863),
.B1(n_861),
.B2(n_851),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_911),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_991),
.A2(n_845),
.B1(n_831),
.B2(n_826),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1033),
.A2(n_638),
.B(n_642),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_993),
.B(n_845),
.Y(n_1073)
);

AOI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_882),
.A2(n_811),
.B1(n_365),
.B2(n_362),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_994),
.A2(n_826),
.B(n_817),
.C(n_813),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1029),
.B(n_576),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_1006),
.B(n_813),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1038),
.A2(n_817),
.B(n_646),
.C(n_650),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_944),
.A2(n_201),
.B1(n_202),
.B2(n_205),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_933),
.A2(n_638),
.B(n_642),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_910),
.B(n_576),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_876),
.B(n_202),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_892),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_910),
.B(n_598),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_1011),
.A2(n_646),
.B(n_650),
.C(n_645),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_928),
.B(n_598),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_962),
.B(n_965),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_895),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_962),
.B(n_205),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_948),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_931),
.A2(n_607),
.B(n_613),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1011),
.A2(n_646),
.B(n_650),
.C(n_645),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_928),
.B(n_598),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_879),
.A2(n_607),
.B(n_613),
.Y(n_1094)
);

OAI22x1_ASAP7_75t_L g1095 ( 
.A1(n_1012),
.A2(n_208),
.B1(n_213),
.B2(n_380),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_876),
.B(n_208),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_944),
.A2(n_213),
.B1(n_378),
.B2(n_380),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_R g1098 ( 
.A(n_950),
.B(n_378),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1009),
.A2(n_475),
.B1(n_478),
.B2(n_476),
.Y(n_1099)
);

AOI21xp33_ASAP7_75t_L g1100 ( 
.A1(n_1012),
.A2(n_321),
.B(n_323),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_993),
.B(n_475),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_882),
.A2(n_630),
.B(n_604),
.C(n_644),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1021),
.B(n_598),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1020),
.A2(n_613),
.B(n_621),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_911),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_SL g1106 ( 
.A(n_904),
.B(n_298),
.Y(n_1106)
);

AOI222xp33_ASAP7_75t_L g1107 ( 
.A1(n_880),
.A2(n_298),
.B1(n_476),
.B2(n_478),
.C1(n_324),
.C2(n_335),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_SL g1108 ( 
.A1(n_982),
.A2(n_918),
.B1(n_988),
.B2(n_888),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_872),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_941),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_985),
.A2(n_700),
.B1(n_691),
.B2(n_667),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_967),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1028),
.A2(n_621),
.B(n_496),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_868),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1009),
.A2(n_700),
.B1(n_691),
.B2(n_667),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_970),
.B(n_631),
.Y(n_1116)
);

BUFx8_ASAP7_75t_L g1117 ( 
.A(n_945),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_SL g1118 ( 
.A(n_904),
.B(n_611),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_872),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_902),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_962),
.B(n_631),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_913),
.Y(n_1122)
);

AO32x1_ASAP7_75t_L g1123 ( 
.A1(n_1031),
.A2(n_644),
.A3(n_632),
.B1(n_477),
.B2(n_8),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_974),
.A2(n_662),
.B(n_477),
.C(n_6),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_886),
.Y(n_1125)
);

AND3x1_ASAP7_75t_SL g1126 ( 
.A(n_1008),
.B(n_0),
.C(n_5),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_1007),
.B(n_496),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_965),
.A2(n_0),
.B1(n_10),
.B2(n_11),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1035),
.B(n_496),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1018),
.A2(n_13),
.B(n_14),
.C(n_16),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1026),
.B(n_74),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_967),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_968),
.A2(n_14),
.B(n_17),
.C(n_19),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_968),
.A2(n_972),
.B(n_909),
.C(n_917),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1034),
.B(n_17),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_972),
.A2(n_22),
.B(n_28),
.C(n_30),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_955),
.A2(n_22),
.B1(n_33),
.B2(n_35),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_SL g1138 ( 
.A1(n_1017),
.A2(n_1007),
.B1(n_870),
.B2(n_1023),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_955),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_1139)
);

INVx3_ASAP7_75t_SL g1140 ( 
.A(n_869),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1026),
.B(n_129),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_935),
.Y(n_1142)
);

O2A1O1Ixp5_ASAP7_75t_L g1143 ( 
.A1(n_964),
.A2(n_131),
.B(n_189),
.C(n_188),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_L g1144 ( 
.A1(n_964),
.A2(n_100),
.B(n_187),
.C(n_183),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_870),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_907),
.A2(n_920),
.B(n_916),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_956),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1030),
.B(n_38),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_871),
.B(n_40),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_987),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_990),
.A2(n_133),
.B(n_178),
.Y(n_1151)
);

NOR2xp67_ASAP7_75t_L g1152 ( 
.A(n_959),
.B(n_116),
.Y(n_1152)
);

NOR2x2_ASAP7_75t_L g1153 ( 
.A(n_1027),
.B(n_952),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_966),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_965),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_881),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_881),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_916),
.A2(n_135),
.B(n_173),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_920),
.A2(n_137),
.B(n_169),
.Y(n_1159)
);

AO21x1_ASAP7_75t_L g1160 ( 
.A1(n_874),
.A2(n_48),
.B(n_50),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_942),
.A2(n_84),
.B(n_166),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_900),
.B(n_50),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_957),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_SL g1164 ( 
.A(n_932),
.B(n_51),
.C(n_54),
.Y(n_1164)
);

NOR2xp67_ASAP7_75t_L g1165 ( 
.A(n_1015),
.B(n_138),
.Y(n_1165)
);

OAI22x1_ASAP7_75t_L g1166 ( 
.A1(n_900),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_890),
.Y(n_1167)
);

INVx5_ASAP7_75t_L g1168 ( 
.A(n_929),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1015),
.B(n_59),
.Y(n_1169)
);

BUFx8_ASAP7_75t_SL g1170 ( 
.A(n_893),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_893),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_966),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_875),
.B(n_61),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1045),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1080),
.A2(n_943),
.B(n_924),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1082),
.B(n_1014),
.Y(n_1176)
);

AO21x2_ASAP7_75t_L g1177 ( 
.A1(n_1050),
.A2(n_925),
.B(n_898),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1096),
.B(n_1016),
.Y(n_1178)
);

NAND2x1_ASAP7_75t_L g1179 ( 
.A(n_1058),
.B(n_929),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1057),
.A2(n_1003),
.A3(n_1002),
.B(n_1010),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1051),
.B(n_1025),
.Y(n_1181)
);

NOR4xp25_ASAP7_75t_L g1182 ( 
.A(n_1130),
.B(n_937),
.C(n_901),
.D(n_995),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1043),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1134),
.A2(n_912),
.B(n_958),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1042),
.A2(n_1107),
.B1(n_1059),
.B2(n_1148),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_1168),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_SL g1187 ( 
.A1(n_1160),
.A2(n_937),
.B(n_1013),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1048),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1060),
.B(n_1061),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1137),
.A2(n_914),
.B1(n_1004),
.B2(n_889),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_R g1191 ( 
.A(n_1063),
.B(n_897),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1044),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1040),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1137),
.A2(n_914),
.B1(n_1004),
.B2(n_889),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_1047),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1154),
.B(n_1027),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1147),
.B(n_1054),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1172),
.B(n_1027),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1171),
.B(n_951),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1083),
.Y(n_1200)
);

AO21x1_ASAP7_75t_L g1201 ( 
.A1(n_1046),
.A2(n_984),
.B(n_978),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1149),
.B(n_1024),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1113),
.A2(n_1104),
.B(n_1091),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1055),
.A2(n_960),
.B(n_963),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1138),
.B(n_1036),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1120),
.B(n_930),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1139),
.A2(n_969),
.B1(n_983),
.B2(n_999),
.Y(n_1207)
);

AO32x2_ASAP7_75t_L g1208 ( 
.A1(n_1139),
.A2(n_903),
.A3(n_954),
.B1(n_906),
.B2(n_922),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1067),
.A2(n_981),
.B(n_1036),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1068),
.A2(n_919),
.A3(n_899),
.B(n_908),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1062),
.A2(n_1036),
.B(n_929),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1066),
.A2(n_1036),
.B(n_929),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1049),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_1068),
.A2(n_896),
.A3(n_915),
.B(n_1037),
.Y(n_1214)
);

AOI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1081),
.A2(n_989),
.B(n_1000),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1125),
.A2(n_996),
.B1(n_969),
.B2(n_999),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1081),
.A2(n_997),
.B(n_1005),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1084),
.A2(n_1093),
.B(n_1086),
.Y(n_1218)
);

OAI22x1_ASAP7_75t_L g1219 ( 
.A1(n_1162),
.A2(n_930),
.B1(n_926),
.B2(n_1001),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1069),
.A2(n_927),
.A3(n_921),
.B(n_980),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1155),
.B(n_1168),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1053),
.B(n_926),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1069),
.A2(n_971),
.A3(n_998),
.B(n_979),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1124),
.A2(n_976),
.B(n_885),
.C(n_894),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1100),
.A2(n_977),
.B(n_996),
.C(n_992),
.Y(n_1225)
);

AOI221xp5_ASAP7_75t_SL g1226 ( 
.A1(n_1133),
.A2(n_1136),
.B1(n_1128),
.B2(n_1150),
.C(n_1095),
.Y(n_1226)
);

NOR2x1_ASAP7_75t_R g1227 ( 
.A(n_1090),
.B(n_953),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1103),
.B(n_977),
.Y(n_1228)
);

NOR4xp25_ASAP7_75t_L g1229 ( 
.A(n_1100),
.B(n_947),
.C(n_938),
.D(n_66),
.Y(n_1229)
);

NOR3xp33_ASAP7_75t_L g1230 ( 
.A(n_1135),
.B(n_999),
.C(n_996),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1109),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1094),
.A2(n_949),
.B(n_936),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1077),
.A2(n_992),
.B1(n_983),
.B2(n_969),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1101),
.B(n_949),
.Y(n_1234)
);

AOI21xp33_ASAP7_75t_L g1235 ( 
.A1(n_1079),
.A2(n_1097),
.B(n_1071),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1102),
.A2(n_1141),
.B(n_1131),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1074),
.B(n_949),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1167),
.B(n_64),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1110),
.B(n_1112),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1141),
.A2(n_144),
.B(n_158),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1085),
.A2(n_160),
.B(n_141),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1143),
.A2(n_65),
.B(n_66),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1144),
.A2(n_1129),
.B(n_1116),
.Y(n_1243)
);

BUFx10_ASAP7_75t_L g1244 ( 
.A(n_1101),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1142),
.B(n_1163),
.Y(n_1245)
);

AO21x1_ASAP7_75t_L g1246 ( 
.A1(n_1071),
.A2(n_1075),
.B(n_1078),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1116),
.A2(n_1076),
.B(n_1151),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1076),
.B(n_1088),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1152),
.A2(n_1073),
.B(n_1165),
.C(n_1092),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1156),
.Y(n_1250)
);

AOI21xp33_ASAP7_75t_L g1251 ( 
.A1(n_1079),
.A2(n_1097),
.B(n_1089),
.Y(n_1251)
);

NOR2xp67_ASAP7_75t_SL g1252 ( 
.A(n_1157),
.B(n_1168),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1108),
.A2(n_1166),
.B1(n_1132),
.B2(n_1122),
.Y(n_1253)
);

AND2x6_ASAP7_75t_L g1254 ( 
.A(n_1073),
.B(n_1070),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1173),
.B(n_1065),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_SL g1256 ( 
.A1(n_1158),
.A2(n_1159),
.B(n_1161),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1056),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1115),
.A2(n_1099),
.A3(n_1123),
.B(n_1064),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1118),
.A2(n_1087),
.B(n_1039),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1169),
.B(n_1119),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1170),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1111),
.A2(n_1121),
.B(n_1070),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1099),
.A2(n_1164),
.B(n_1123),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_1048),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1106),
.B(n_1145),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1105),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1126),
.A2(n_1153),
.A3(n_1127),
.B(n_1114),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1127),
.B(n_1048),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1140),
.B(n_1127),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1117),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1098),
.A2(n_1057),
.A3(n_1160),
.B(n_1069),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1117),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1057),
.A2(n_1160),
.A3(n_1068),
.B(n_1069),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1082),
.B(n_975),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1082),
.B(n_975),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1043),
.B(n_612),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1050),
.A2(n_628),
.B(n_1134),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1042),
.A2(n_812),
.B(n_986),
.C(n_975),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_SL g1279 ( 
.A(n_1058),
.B(n_1019),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1154),
.B(n_993),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1154),
.B(n_717),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1080),
.A2(n_1072),
.B(n_1146),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1050),
.A2(n_628),
.B(n_1134),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1040),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1041),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1045),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1082),
.B(n_975),
.Y(n_1287)
);

OR2x6_ASAP7_75t_L g1288 ( 
.A(n_1157),
.B(n_993),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1058),
.B(n_1155),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1050),
.A2(n_1080),
.B(n_1072),
.Y(n_1290)
);

AOI211x1_ASAP7_75t_L g1291 ( 
.A1(n_1137),
.A2(n_1139),
.B(n_1160),
.C(n_1128),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1042),
.A2(n_812),
.B(n_986),
.C(n_975),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1080),
.A2(n_1072),
.B(n_1146),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1082),
.B(n_1019),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1050),
.A2(n_628),
.B(n_1134),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_1052),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1080),
.A2(n_1072),
.B(n_1146),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1080),
.A2(n_1072),
.B(n_1146),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1082),
.B(n_975),
.Y(n_1299)
);

AOI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1042),
.A2(n_1038),
.B1(n_731),
.B2(n_818),
.C(n_1012),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1050),
.A2(n_628),
.B(n_1134),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1174),
.Y(n_1302)
);

OA21x2_ASAP7_75t_L g1303 ( 
.A1(n_1175),
.A2(n_1236),
.B(n_1218),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1189),
.B(n_1197),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1203),
.A2(n_1293),
.B(n_1282),
.Y(n_1305)
);

O2A1O1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1278),
.A2(n_1292),
.B(n_1275),
.C(n_1287),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1246),
.A2(n_1201),
.A3(n_1295),
.B(n_1283),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1183),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1223),
.Y(n_1309)
);

OA21x2_ASAP7_75t_L g1310 ( 
.A1(n_1236),
.A2(n_1298),
.B(n_1297),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1254),
.Y(n_1311)
);

INVx8_ASAP7_75t_L g1312 ( 
.A(n_1268),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1277),
.A2(n_1301),
.B(n_1209),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1281),
.B(n_1206),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1294),
.A2(n_1253),
.B1(n_1299),
.B2(n_1274),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_1193),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1196),
.B(n_1198),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1176),
.B(n_1178),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_L g1319 ( 
.A(n_1231),
.B(n_1276),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1204),
.A2(n_1184),
.B(n_1290),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1225),
.A2(n_1249),
.B(n_1241),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1186),
.B(n_1252),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1290),
.A2(n_1177),
.B(n_1241),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1220),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1177),
.A2(n_1181),
.B(n_1256),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1300),
.B(n_1202),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1211),
.A2(n_1212),
.B(n_1215),
.Y(n_1327)
);

OR2x6_ASAP7_75t_L g1328 ( 
.A(n_1259),
.B(n_1207),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1253),
.A2(n_1194),
.B1(n_1190),
.B2(n_1279),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1223),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1286),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1199),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1199),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1262),
.A2(n_1240),
.B(n_1232),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1244),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1223),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1235),
.A2(n_1187),
.B(n_1182),
.Y(n_1337)
);

INVx4_ASAP7_75t_L g1338 ( 
.A(n_1186),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1224),
.A2(n_1226),
.B(n_1222),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1247),
.A2(n_1243),
.B(n_1216),
.Y(n_1340)
);

CKINVDCx6p67_ASAP7_75t_R g1341 ( 
.A(n_1261),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1185),
.A2(n_1291),
.B1(n_1272),
.B2(n_1296),
.Y(n_1342)
);

NAND2x1p5_ASAP7_75t_L g1343 ( 
.A(n_1205),
.B(n_1179),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_SL g1344 ( 
.A(n_1284),
.B(n_1227),
.Y(n_1344)
);

AOI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1219),
.A2(n_1237),
.B(n_1242),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1255),
.B(n_1183),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1254),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1195),
.B(n_1260),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1226),
.A2(n_1248),
.B(n_1251),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1251),
.A2(n_1228),
.B(n_1238),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1191),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1242),
.A2(n_1233),
.B(n_1245),
.Y(n_1352)
);

O2A1O1Ixp33_ASAP7_75t_SL g1353 ( 
.A1(n_1233),
.A2(n_1245),
.B(n_1265),
.C(n_1257),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1289),
.A2(n_1221),
.B(n_1213),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1273),
.A2(n_1208),
.B(n_1192),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1182),
.A2(n_1279),
.B(n_1230),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1280),
.B(n_1234),
.Y(n_1357)
);

INVx4_ASAP7_75t_SL g1358 ( 
.A(n_1254),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1214),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1266),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1188),
.Y(n_1361)
);

OR2x6_ASAP7_75t_L g1362 ( 
.A(n_1288),
.B(n_1268),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1273),
.A2(n_1208),
.B(n_1210),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1263),
.A2(n_1200),
.B1(n_1254),
.B2(n_1285),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_L g1365 ( 
.A(n_1229),
.B(n_1269),
.C(n_1250),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1220),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1270),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1268),
.A2(n_1288),
.B(n_1210),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1210),
.A2(n_1180),
.B(n_1273),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1244),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1180),
.A2(n_1271),
.B(n_1258),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1258),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_1188),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1227),
.B(n_1188),
.Y(n_1374)
);

AO32x2_ASAP7_75t_L g1375 ( 
.A1(n_1271),
.A2(n_1258),
.A3(n_1180),
.B1(n_1267),
.B2(n_1264),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1278),
.A2(n_812),
.B(n_1292),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1274),
.A2(n_1287),
.B1(n_1299),
.B2(n_1275),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1281),
.B(n_1206),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1193),
.Y(n_1379)
);

OA21x2_ASAP7_75t_L g1380 ( 
.A1(n_1175),
.A2(n_1236),
.B(n_1218),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1278),
.A2(n_812),
.B(n_1292),
.Y(n_1382)
);

AOI21xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1294),
.A2(n_1019),
.B(n_804),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1203),
.A2(n_1293),
.B(n_1282),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1203),
.A2(n_1293),
.B(n_1282),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1175),
.A2(n_1236),
.B(n_1218),
.Y(n_1386)
);

AOI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1215),
.A2(n_1217),
.B(n_1184),
.Y(n_1387)
);

BUFx10_ASAP7_75t_L g1388 ( 
.A(n_1193),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1183),
.Y(n_1390)
);

OAI221xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1300),
.A2(n_1185),
.B1(n_521),
.B2(n_535),
.C(n_508),
.Y(n_1391)
);

BUFx4_ASAP7_75t_SL g1392 ( 
.A(n_1272),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1277),
.A2(n_1295),
.B(n_1283),
.Y(n_1393)
);

INVx2_ASAP7_75t_SL g1394 ( 
.A(n_1239),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1186),
.B(n_1058),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1200),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1300),
.A2(n_1235),
.B(n_1292),
.C(n_1278),
.Y(n_1399)
);

NAND3x1_ASAP7_75t_L g1400 ( 
.A(n_1294),
.B(n_1038),
.C(n_1300),
.Y(n_1400)
);

NAND3xp33_ASAP7_75t_L g1401 ( 
.A(n_1300),
.B(n_1042),
.C(n_1185),
.Y(n_1401)
);

AOI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1215),
.A2(n_1217),
.B(n_1184),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1185),
.B(n_1300),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1188),
.Y(n_1404)
);

INVx5_ASAP7_75t_L g1405 ( 
.A(n_1268),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1203),
.A2(n_1293),
.B(n_1282),
.Y(n_1407)
);

AO31x2_ASAP7_75t_L g1408 ( 
.A1(n_1246),
.A2(n_1201),
.A3(n_1218),
.B(n_1277),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1296),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1294),
.A2(n_1019),
.B1(n_1275),
.B2(n_1274),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1223),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1203),
.A2(n_1293),
.B(n_1282),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1278),
.A2(n_812),
.B(n_1292),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1239),
.B(n_1189),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1281),
.B(n_1206),
.Y(n_1415)
);

CKINVDCx11_ASAP7_75t_R g1416 ( 
.A(n_1296),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1174),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1278),
.A2(n_812),
.B(n_1292),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1294),
.A2(n_1019),
.B1(n_1275),
.B2(n_1274),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1300),
.A2(n_1235),
.B(n_1292),
.C(n_1278),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1203),
.A2(n_1293),
.B(n_1282),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1300),
.A2(n_1294),
.B1(n_1019),
.B2(n_1042),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1317),
.B(n_1314),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1332),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1416),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1400),
.A2(n_1422),
.B1(n_1391),
.B2(n_1329),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1377),
.B(n_1318),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1377),
.B(n_1389),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1389),
.B(n_1396),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1396),
.B(n_1326),
.Y(n_1430)
);

XOR2xp5_ASAP7_75t_L g1431 ( 
.A(n_1409),
.B(n_1316),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1323),
.A2(n_1340),
.B(n_1320),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1304),
.B(n_1381),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1376),
.A2(n_1413),
.B(n_1382),
.Y(n_1434)
);

INVx5_ASAP7_75t_L g1435 ( 
.A(n_1362),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1378),
.B(n_1415),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1302),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1320),
.A2(n_1321),
.B(n_1323),
.Y(n_1438)
);

O2A1O1Ixp5_ASAP7_75t_L g1439 ( 
.A1(n_1403),
.A2(n_1418),
.B(n_1420),
.C(n_1399),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1398),
.B(n_1406),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1397),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1332),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1414),
.B(n_1403),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1394),
.B(n_1357),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1348),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1351),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1346),
.B(n_1401),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1308),
.B(n_1390),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1357),
.B(n_1329),
.Y(n_1449)
);

INVx5_ASAP7_75t_SL g1450 ( 
.A(n_1341),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1409),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1331),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1324),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1306),
.B(n_1410),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_SL g1455 ( 
.A1(n_1391),
.A2(n_1356),
.B(n_1325),
.C(n_1347),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1419),
.B(n_1399),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1369),
.A2(n_1327),
.B(n_1371),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1366),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1365),
.B(n_1420),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1315),
.A2(n_1342),
.B1(n_1362),
.B2(n_1356),
.Y(n_1460)
);

CKINVDCx16_ASAP7_75t_R g1461 ( 
.A(n_1344),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1333),
.Y(n_1462)
);

NOR2xp67_ASAP7_75t_L g1463 ( 
.A(n_1351),
.B(n_1383),
.Y(n_1463)
);

BUFx12f_ASAP7_75t_L g1464 ( 
.A(n_1416),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1310),
.A2(n_1393),
.B(n_1313),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1362),
.A2(n_1395),
.B(n_1322),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1333),
.B(n_1360),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1417),
.B(n_1337),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1319),
.B(n_1349),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1337),
.B(n_1350),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1312),
.A2(n_1405),
.B(n_1364),
.C(n_1374),
.Y(n_1471)
);

A2O1A1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1312),
.A2(n_1405),
.B(n_1364),
.C(n_1374),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1350),
.B(n_1312),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1373),
.B(n_1361),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1361),
.B(n_1404),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1310),
.A2(n_1393),
.B(n_1303),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1353),
.A2(n_1343),
.B(n_1328),
.C(n_1350),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1303),
.A2(n_1386),
.B(n_1380),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1395),
.A2(n_1322),
.B(n_1370),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1343),
.A2(n_1328),
.B(n_1339),
.C(n_1347),
.Y(n_1480)
);

CKINVDCx8_ASAP7_75t_R g1481 ( 
.A(n_1316),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1370),
.A2(n_1338),
.B(n_1328),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1358),
.B(n_1405),
.Y(n_1483)
);

O2A1O1Ixp5_ASAP7_75t_L g1484 ( 
.A1(n_1368),
.A2(n_1345),
.B(n_1402),
.C(n_1387),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1358),
.B(n_1311),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1338),
.A2(n_1358),
.B(n_1339),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1311),
.B(n_1354),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1339),
.A2(n_1359),
.B(n_1411),
.C(n_1309),
.Y(n_1488)
);

OAI31xp33_ASAP7_75t_L g1489 ( 
.A1(n_1309),
.A2(n_1411),
.A3(n_1330),
.B(n_1336),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1367),
.A2(n_1335),
.B1(n_1379),
.B2(n_1404),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1367),
.A2(n_1335),
.B1(n_1379),
.B2(n_1404),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1361),
.B(n_1375),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1408),
.B(n_1355),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1336),
.A2(n_1372),
.B(n_1380),
.C(n_1386),
.Y(n_1494)
);

O2A1O1Ixp5_ASAP7_75t_L g1495 ( 
.A1(n_1372),
.A2(n_1408),
.B(n_1307),
.C(n_1375),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1375),
.B(n_1355),
.Y(n_1496)
);

O2A1O1Ixp33_ASAP7_75t_L g1497 ( 
.A1(n_1355),
.A2(n_1363),
.B(n_1375),
.C(n_1408),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1352),
.B(n_1388),
.Y(n_1498)
);

AOI21x1_ASAP7_75t_SL g1499 ( 
.A1(n_1307),
.A2(n_1408),
.B(n_1334),
.Y(n_1499)
);

AND2x2_ASAP7_75t_SL g1500 ( 
.A(n_1363),
.B(n_1392),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1307),
.B(n_1305),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1388),
.B(n_1363),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1392),
.A2(n_1421),
.B(n_1384),
.C(n_1385),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1407),
.A2(n_1300),
.B(n_1401),
.C(n_1185),
.Y(n_1504)
);

A2O1A1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1412),
.A2(n_1300),
.B(n_1401),
.C(n_1185),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1403),
.A2(n_1292),
.B(n_1278),
.C(n_1275),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1401),
.B(n_1300),
.C(n_1403),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1400),
.A2(n_1019),
.B1(n_1294),
.B2(n_1422),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1403),
.A2(n_1292),
.B(n_1278),
.C(n_1275),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1317),
.B(n_1314),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_SL g1511 ( 
.A1(n_1326),
.A2(n_986),
.B(n_1274),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1324),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1409),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1320),
.A2(n_1321),
.B(n_1323),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1332),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1323),
.A2(n_1340),
.B(n_1320),
.Y(n_1516)
);

NOR2xp67_ASAP7_75t_L g1517 ( 
.A(n_1304),
.B(n_1250),
.Y(n_1517)
);

O2A1O1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1403),
.A2(n_1292),
.B(n_1278),
.C(n_1275),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1400),
.A2(n_1019),
.B1(n_1294),
.B2(n_1422),
.Y(n_1519)
);

NOR2xp67_ASAP7_75t_L g1520 ( 
.A(n_1304),
.B(n_1250),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1302),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1320),
.A2(n_1321),
.B(n_1323),
.Y(n_1522)
);

AOI21x1_ASAP7_75t_SL g1523 ( 
.A1(n_1326),
.A2(n_986),
.B(n_1274),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1397),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1358),
.B(n_1362),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1410),
.B(n_1294),
.Y(n_1526)
);

O2A1O1Ixp5_ASAP7_75t_L g1527 ( 
.A1(n_1403),
.A2(n_1382),
.B(n_1413),
.C(n_1376),
.Y(n_1527)
);

BUFx12f_ASAP7_75t_L g1528 ( 
.A(n_1416),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1492),
.B(n_1496),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1435),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1438),
.A2(n_1522),
.B(n_1514),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1438),
.A2(n_1522),
.B(n_1514),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1470),
.B(n_1468),
.Y(n_1533)
);

OAI33xp33_ASAP7_75t_L g1534 ( 
.A1(n_1426),
.A2(n_1519),
.A3(n_1508),
.B1(n_1507),
.B2(n_1428),
.B3(n_1459),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1427),
.B(n_1430),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1453),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1434),
.B(n_1477),
.Y(n_1537)
);

OR2x6_ASAP7_75t_L g1538 ( 
.A(n_1477),
.B(n_1480),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1457),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1476),
.A2(n_1465),
.B(n_1478),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1469),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1458),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1501),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1512),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1502),
.B(n_1501),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1437),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1525),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1495),
.B(n_1473),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1498),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1487),
.Y(n_1550)
);

BUFx12f_ASAP7_75t_L g1551 ( 
.A(n_1425),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1445),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1456),
.A2(n_1454),
.B1(n_1526),
.B2(n_1460),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1521),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1443),
.B(n_1429),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1495),
.B(n_1432),
.Y(n_1556)
);

AOI222xp33_ASAP7_75t_L g1557 ( 
.A1(n_1440),
.A2(n_1505),
.B1(n_1504),
.B2(n_1433),
.C1(n_1464),
.C2(n_1528),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1516),
.B(n_1500),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1488),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1488),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1489),
.B(n_1452),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1455),
.B(n_1471),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1497),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1497),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1494),
.B(n_1527),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1484),
.A2(n_1527),
.B(n_1439),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1442),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1484),
.B(n_1439),
.Y(n_1568)
);

NAND3x1_ASAP7_75t_L g1569 ( 
.A(n_1449),
.B(n_1444),
.C(n_1467),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1448),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1423),
.B(n_1510),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1503),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1506),
.Y(n_1573)
);

AO21x2_ASAP7_75t_L g1574 ( 
.A1(n_1472),
.A2(n_1486),
.B(n_1518),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1441),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1506),
.Y(n_1576)
);

AO21x2_ASAP7_75t_L g1577 ( 
.A1(n_1509),
.A2(n_1518),
.B(n_1499),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1447),
.B(n_1509),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1525),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1539),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1529),
.B(n_1436),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1541),
.B(n_1520),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1529),
.B(n_1475),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1533),
.B(n_1524),
.Y(n_1584)
);

NAND3xp33_ASAP7_75t_L g1585 ( 
.A(n_1557),
.B(n_1517),
.C(n_1479),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1543),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1541),
.B(n_1474),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1543),
.Y(n_1588)
);

NOR2xp67_ASAP7_75t_L g1589 ( 
.A(n_1533),
.B(n_1490),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1546),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1546),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1546),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1533),
.B(n_1491),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1544),
.Y(n_1594)
);

AOI222xp33_ASAP7_75t_L g1595 ( 
.A1(n_1534),
.A2(n_1463),
.B1(n_1513),
.B2(n_1451),
.C1(n_1450),
.C2(n_1446),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1567),
.Y(n_1596)
);

OAI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1578),
.A2(n_1461),
.B1(n_1515),
.B2(n_1462),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1553),
.A2(n_1483),
.B1(n_1466),
.B2(n_1450),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1548),
.B(n_1499),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1536),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1548),
.B(n_1424),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1548),
.B(n_1483),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1558),
.B(n_1485),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1554),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_SL g1605 ( 
.A1(n_1578),
.A2(n_1450),
.B1(n_1523),
.B2(n_1511),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1567),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_L g1607 ( 
.A(n_1574),
.B(n_1482),
.Y(n_1607)
);

OAI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1585),
.A2(n_1553),
.B1(n_1557),
.B2(n_1562),
.C(n_1537),
.Y(n_1608)
);

NOR4xp25_ASAP7_75t_SL g1609 ( 
.A(n_1594),
.B(n_1575),
.C(n_1572),
.D(n_1549),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1586),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1602),
.B(n_1545),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1582),
.B(n_1535),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1590),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1586),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1600),
.B(n_1549),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1590),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1595),
.A2(n_1534),
.B1(n_1537),
.B2(n_1573),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1590),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1580),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1600),
.B(n_1563),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1602),
.B(n_1550),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1585),
.A2(n_1562),
.B1(n_1576),
.B2(n_1573),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1602),
.B(n_1550),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1591),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1595),
.A2(n_1537),
.B1(n_1576),
.B2(n_1574),
.Y(n_1625)
);

NOR4xp25_ASAP7_75t_SL g1626 ( 
.A(n_1594),
.B(n_1575),
.C(n_1572),
.D(n_1559),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1605),
.A2(n_1562),
.B1(n_1537),
.B2(n_1569),
.Y(n_1627)
);

OAI211xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1582),
.A2(n_1535),
.B(n_1555),
.C(n_1552),
.Y(n_1628)
);

OAI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1605),
.A2(n_1537),
.B1(n_1569),
.B2(n_1538),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1598),
.A2(n_1537),
.B1(n_1569),
.B2(n_1538),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1586),
.B(n_1588),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1583),
.B(n_1550),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1598),
.A2(n_1574),
.B1(n_1532),
.B2(n_1531),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1592),
.Y(n_1634)
);

OAI31xp33_ASAP7_75t_L g1635 ( 
.A1(n_1597),
.A2(n_1568),
.A3(n_1565),
.B(n_1555),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1607),
.A2(n_1538),
.B1(n_1552),
.B2(n_1579),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1596),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1586),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1583),
.B(n_1550),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1592),
.Y(n_1640)
);

OAI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1589),
.A2(n_1538),
.B1(n_1570),
.B2(n_1565),
.C(n_1564),
.Y(n_1641)
);

OAI211xp5_ASAP7_75t_L g1642 ( 
.A1(n_1589),
.A2(n_1565),
.B(n_1568),
.C(n_1566),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1597),
.A2(n_1538),
.B1(n_1579),
.B2(n_1547),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1593),
.A2(n_1531),
.B1(n_1532),
.B2(n_1577),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1601),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1584),
.Y(n_1646)
);

OA222x2_ASAP7_75t_L g1647 ( 
.A1(n_1593),
.A2(n_1538),
.B1(n_1561),
.B2(n_1560),
.C1(n_1559),
.C2(n_1601),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1587),
.B(n_1570),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1592),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1619),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1613),
.Y(n_1651)
);

AND2x6_ASAP7_75t_SL g1652 ( 
.A(n_1612),
.B(n_1551),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1613),
.Y(n_1653)
);

INVx4_ASAP7_75t_SL g1654 ( 
.A(n_1637),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1646),
.B(n_1584),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1619),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1616),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1637),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1616),
.Y(n_1659)
);

AO21x1_ASAP7_75t_L g1660 ( 
.A1(n_1635),
.A2(n_1599),
.B(n_1568),
.Y(n_1660)
);

NOR2x1_ASAP7_75t_L g1661 ( 
.A(n_1642),
.B(n_1596),
.Y(n_1661)
);

CKINVDCx16_ASAP7_75t_R g1662 ( 
.A(n_1627),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1618),
.Y(n_1663)
);

INVxp67_ASAP7_75t_SL g1664 ( 
.A(n_1620),
.Y(n_1664)
);

OR2x6_ASAP7_75t_L g1665 ( 
.A(n_1629),
.B(n_1530),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1624),
.Y(n_1666)
);

INVxp67_ASAP7_75t_SL g1667 ( 
.A(n_1615),
.Y(n_1667)
);

NOR2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1647),
.B(n_1551),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1631),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1624),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1615),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1648),
.B(n_1606),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1644),
.A2(n_1540),
.B(n_1556),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1645),
.Y(n_1674)
);

OR2x6_ASAP7_75t_L g1675 ( 
.A(n_1630),
.B(n_1530),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1631),
.B(n_1645),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1628),
.B(n_1551),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_SL g1678 ( 
.A(n_1635),
.B(n_1606),
.C(n_1593),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1631),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1610),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1621),
.B(n_1599),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1651),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1664),
.B(n_1622),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_SL g1684 ( 
.A(n_1662),
.B(n_1661),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1662),
.A2(n_1608),
.B1(n_1531),
.B2(n_1532),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1654),
.B(n_1647),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1651),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1676),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1680),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1654),
.B(n_1669),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1653),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1654),
.B(n_1621),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1654),
.B(n_1623),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1654),
.B(n_1623),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1653),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1668),
.A2(n_1625),
.B1(n_1633),
.B2(n_1617),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1667),
.B(n_1601),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1657),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1657),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1668),
.A2(n_1643),
.B1(n_1636),
.B2(n_1641),
.Y(n_1700)
);

NAND3xp33_ASAP7_75t_L g1701 ( 
.A(n_1661),
.B(n_1626),
.C(n_1609),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1671),
.B(n_1581),
.Y(n_1702)
);

NAND4xp25_ASAP7_75t_L g1703 ( 
.A(n_1678),
.B(n_1599),
.C(n_1587),
.D(n_1560),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1669),
.B(n_1681),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1677),
.A2(n_1638),
.B1(n_1614),
.B2(n_1610),
.C(n_1604),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1680),
.Y(n_1706)
);

OAI33xp33_ASAP7_75t_L g1707 ( 
.A1(n_1659),
.A2(n_1604),
.A3(n_1649),
.B1(n_1640),
.B2(n_1634),
.B3(n_1542),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1679),
.B(n_1638),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1665),
.A2(n_1566),
.B1(n_1561),
.B2(n_1571),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1650),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1679),
.B(n_1676),
.Y(n_1711)
);

NOR2xp67_ASAP7_75t_L g1712 ( 
.A(n_1679),
.B(n_1634),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1676),
.B(n_1611),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1650),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1655),
.B(n_1665),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1676),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1665),
.B(n_1632),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1663),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1690),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1686),
.B(n_1665),
.Y(n_1720)
);

NOR2x1p5_ASAP7_75t_SL g1721 ( 
.A(n_1689),
.B(n_1656),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1686),
.B(n_1675),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1682),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1697),
.B(n_1672),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1689),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1692),
.B(n_1675),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1692),
.B(n_1675),
.Y(n_1727)
);

NAND2x1p5_ASAP7_75t_L g1728 ( 
.A(n_1690),
.B(n_1658),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1693),
.B(n_1675),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1689),
.Y(n_1730)
);

OR2x6_ASAP7_75t_L g1731 ( 
.A(n_1701),
.B(n_1675),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1706),
.B(n_1663),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1697),
.B(n_1660),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1682),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1706),
.B(n_1666),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1687),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1693),
.B(n_1694),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1687),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1710),
.Y(n_1739)
);

NAND2x1_ASAP7_75t_SL g1740 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1710),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1691),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1691),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1710),
.Y(n_1744)
);

AOI21xp33_ASAP7_75t_L g1745 ( 
.A1(n_1684),
.A2(n_1660),
.B(n_1673),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1695),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1695),
.Y(n_1747)
);

A2O1A1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1684),
.A2(n_1652),
.B(n_1674),
.C(n_1603),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1713),
.B(n_1688),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1683),
.B(n_1670),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1714),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1713),
.B(n_1639),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1688),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1716),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1698),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1730),
.B(n_1683),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1737),
.B(n_1716),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1737),
.B(n_1704),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1719),
.B(n_1685),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1723),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1719),
.B(n_1705),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1755),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1755),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1728),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1754),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1723),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1748),
.A2(n_1696),
.B1(n_1700),
.B2(n_1701),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1734),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1728),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1730),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1725),
.Y(n_1771)
);

OR2x6_ASAP7_75t_L g1772 ( 
.A(n_1728),
.B(n_1688),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1740),
.Y(n_1773)
);

CKINVDCx16_ASAP7_75t_R g1774 ( 
.A(n_1731),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1733),
.B(n_1724),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1740),
.Y(n_1776)
);

INVx2_ASAP7_75t_SL g1777 ( 
.A(n_1753),
.Y(n_1777)
);

INVx4_ASAP7_75t_L g1778 ( 
.A(n_1753),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1731),
.A2(n_1715),
.B1(n_1702),
.B2(n_1709),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1734),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1753),
.Y(n_1781)
);

OAI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1745),
.A2(n_1703),
.B(n_1705),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1770),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1771),
.Y(n_1784)
);

AOI222xp33_ASAP7_75t_L g1785 ( 
.A1(n_1767),
.A2(n_1721),
.B1(n_1720),
.B2(n_1750),
.C1(n_1709),
.C2(n_1722),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1758),
.B(n_1722),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1765),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1774),
.B(n_1725),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1758),
.B(n_1750),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1782),
.A2(n_1745),
.B(n_1720),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1756),
.B(n_1764),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1779),
.A2(n_1731),
.B(n_1733),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1756),
.B(n_1769),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1760),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1777),
.B(n_1749),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1777),
.B(n_1749),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_SL g1797 ( 
.A1(n_1761),
.A2(n_1731),
.B1(n_1729),
.B2(n_1726),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1775),
.B(n_1724),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1778),
.Y(n_1799)
);

AOI221x1_ASAP7_75t_L g1800 ( 
.A1(n_1778),
.A2(n_1781),
.B1(n_1776),
.B2(n_1773),
.C(n_1759),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1757),
.B(n_1703),
.Y(n_1801)
);

OAI322xp33_ASAP7_75t_L g1802 ( 
.A1(n_1775),
.A2(n_1773),
.A3(n_1776),
.B1(n_1760),
.B2(n_1780),
.C1(n_1763),
.C2(n_1762),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1778),
.B(n_1726),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1786),
.B(n_1757),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1803),
.Y(n_1805)
);

INVxp33_ASAP7_75t_L g1806 ( 
.A(n_1788),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1785),
.A2(n_1731),
.B1(n_1772),
.B2(n_1757),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1783),
.B(n_1781),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1787),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1784),
.B(n_1781),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1803),
.B(n_1772),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1797),
.B(n_1727),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1800),
.B(n_1762),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1799),
.B(n_1772),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1795),
.B(n_1727),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1796),
.B(n_1729),
.Y(n_1816)
);

OAI211xp5_ASAP7_75t_L g1817 ( 
.A1(n_1807),
.A2(n_1790),
.B(n_1792),
.C(n_1793),
.Y(n_1817)
);

AOI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1813),
.A2(n_1802),
.B(n_1791),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1807),
.A2(n_1802),
.B(n_1798),
.Y(n_1819)
);

AOI221x1_ASAP7_75t_L g1820 ( 
.A1(n_1808),
.A2(n_1799),
.B1(n_1794),
.B2(n_1780),
.C(n_1766),
.Y(n_1820)
);

OAI211xp5_ASAP7_75t_L g1821 ( 
.A1(n_1805),
.A2(n_1801),
.B(n_1789),
.C(n_1766),
.Y(n_1821)
);

OAI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1812),
.A2(n_1772),
.B1(n_1715),
.B2(n_1732),
.C(n_1735),
.Y(n_1822)
);

NOR4xp25_ASAP7_75t_L g1823 ( 
.A(n_1809),
.B(n_1768),
.C(n_1763),
.D(n_1732),
.Y(n_1823)
);

NOR4xp25_ASAP7_75t_L g1824 ( 
.A(n_1808),
.B(n_1810),
.C(n_1814),
.D(n_1815),
.Y(n_1824)
);

NOR2x1_ASAP7_75t_L g1825 ( 
.A(n_1811),
.B(n_1768),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1810),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1806),
.A2(n_1735),
.B1(n_1742),
.B2(n_1747),
.C(n_1746),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1825),
.Y(n_1828)
);

OAI21xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1818),
.A2(n_1816),
.B(n_1804),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1817),
.A2(n_1814),
.B(n_1811),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1819),
.A2(n_1688),
.B1(n_1751),
.B2(n_1739),
.Y(n_1831)
);

AOI211xp5_ASAP7_75t_L g1832 ( 
.A1(n_1824),
.A2(n_1742),
.B(n_1738),
.C(n_1747),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1826),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1828),
.Y(n_1834)
);

NAND3xp33_ASAP7_75t_L g1835 ( 
.A(n_1830),
.B(n_1831),
.C(n_1829),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1833),
.B(n_1821),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1832),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1828),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1829),
.B(n_1823),
.Y(n_1839)
);

NOR3xp33_ASAP7_75t_L g1840 ( 
.A(n_1830),
.B(n_1822),
.C(n_1827),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_R g1841 ( 
.A(n_1836),
.B(n_1481),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1840),
.B(n_1820),
.Y(n_1842)
);

OAI22xp33_ASAP7_75t_SL g1843 ( 
.A1(n_1839),
.A2(n_1736),
.B1(n_1738),
.B2(n_1746),
.Y(n_1843)
);

AOI321xp33_ASAP7_75t_L g1844 ( 
.A1(n_1837),
.A2(n_1739),
.A3(n_1751),
.B1(n_1744),
.B2(n_1741),
.C(n_1743),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1835),
.A2(n_1736),
.B1(n_1743),
.B2(n_1712),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1842),
.B(n_1834),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1843),
.B(n_1838),
.Y(n_1847)
);

XNOR2xp5_ASAP7_75t_L g1848 ( 
.A(n_1845),
.B(n_1431),
.Y(n_1848)
);

NAND3x1_ASAP7_75t_L g1849 ( 
.A(n_1847),
.B(n_1841),
.C(n_1844),
.Y(n_1849)
);

AOI322xp5_ASAP7_75t_L g1850 ( 
.A1(n_1849),
.A2(n_1848),
.A3(n_1846),
.B1(n_1739),
.B2(n_1751),
.C1(n_1744),
.C2(n_1741),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1850),
.B(n_1721),
.Y(n_1851)
);

AOI222xp33_ASAP7_75t_L g1852 ( 
.A1(n_1850),
.A2(n_1744),
.B1(n_1741),
.B2(n_1707),
.C1(n_1712),
.C2(n_1699),
.Y(n_1852)
);

INVx4_ASAP7_75t_L g1853 ( 
.A(n_1851),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1852),
.B(n_1752),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1854),
.Y(n_1855)
);

OAI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1853),
.A2(n_1714),
.B1(n_1711),
.B2(n_1698),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1855),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1857),
.B(n_1853),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_SL g1859 ( 
.A1(n_1858),
.A2(n_1856),
.B(n_1717),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1859),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1711),
.B1(n_1708),
.B2(n_1717),
.Y(n_1861)
);

AOI211xp5_ASAP7_75t_L g1862 ( 
.A1(n_1861),
.A2(n_1714),
.B(n_1718),
.C(n_1699),
.Y(n_1862)
);


endmodule