module real_jpeg_23529_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_66),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_2),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_72),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_5),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_5),
.A2(n_67),
.B1(n_68),
.B2(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_93),
.Y(n_124)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_8),
.A2(n_45),
.B1(n_54),
.B2(n_55),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_8),
.A2(n_45),
.B1(n_67),
.B2(n_68),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_9),
.A2(n_39),
.B1(n_54),
.B2(n_55),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_9),
.A2(n_39),
.B1(n_67),
.B2(n_68),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_49),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_10),
.A2(n_49),
.B1(n_67),
.B2(n_68),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_10),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_12),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_67),
.C(n_85),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_77),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_12),
.B(n_61),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_12),
.A2(n_69),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_12),
.B(n_98),
.Y(n_220)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_15),
.Y(n_172)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_15),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_112),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_19),
.B(n_112),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_80),
.C(n_100),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_20),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_62),
.B2(n_79),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_46),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_23),
.B(n_46),
.C(n_79),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_37),
.B2(n_43),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_25),
.A2(n_75),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_25),
.A2(n_44),
.B1(n_98),
.B2(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_27),
.A2(n_30),
.B(n_75),
.C(n_78),
.Y(n_74)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_29),
.C(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_29),
.A2(n_30),
.B1(n_53),
.B2(n_56),
.Y(n_57)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g197 ( 
.A(n_30),
.B(n_77),
.CON(n_197),
.SN(n_197)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_30),
.B(n_54),
.C(n_56),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_58),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_51),
.B1(n_61),
.B2(n_96),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_50),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_50),
.A2(n_52),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_51),
.A2(n_61),
.B1(n_197),
.B2(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_52)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_53),
.A2(n_55),
.B(n_197),
.C(n_198),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_54),
.A2(n_55),
.B1(n_85),
.B2(n_87),
.Y(n_84)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_55),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_59),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_61),
.B(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_74),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_63),
.B(n_74),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_65),
.A2(n_130),
.B(n_132),
.Y(n_221)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_70),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_68),
.B1(n_85),
.B2(n_87),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_68),
.B(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_71),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_107),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_69),
.A2(n_129),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_69),
.A2(n_73),
.B1(n_170),
.B2(n_179),
.Y(n_189)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_70),
.Y(n_186)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.CON(n_75),
.SN(n_75)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_77),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_77),
.B(n_88),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_80),
.A2(n_100),
.B1(n_101),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_80),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_95),
.C(n_97),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_81),
.A2(n_82),
.B1(n_95),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_89),
.B(n_91),
.Y(n_82)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_83),
.A2(n_88),
.B1(n_109),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_83),
.A2(n_88),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_83),
.A2(n_88),
.B1(n_155),
.B2(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_83),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_90),
.B(n_94),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_94),
.A2(n_111),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_95),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_96),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_97),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_108),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_108),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_104),
.A2(n_131),
.B(n_168),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_138),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_125),
.B1(n_136),
.B2(n_137),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_133),
.B2(n_134),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_247),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_242),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_232),
.B(n_241),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_210),
.B(n_231),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_193),
.B(n_209),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_165),
.B(n_192),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_156),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_152),
.B1(n_153),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_208)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_176),
.B(n_191),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_174),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_173),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_187),
.B(n_190),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_183),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_188),
.B(n_189),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_208),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_208),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_203),
.C(n_206),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_207),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_211),
.B(n_212),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_223),
.B2(n_224),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_226),
.C(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_219),
.C(n_222),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_229),
.B2(n_230),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_240),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_236),
.C(n_237),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_244),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);


endmodule