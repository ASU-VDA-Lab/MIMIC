module fake_jpeg_1909_n_123 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_123);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_6),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_49),
.Y(n_60)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_35),
.B1(n_41),
.B2(n_43),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_46),
.B1(n_49),
.B2(n_33),
.Y(n_68)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_38),
.B(n_47),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_41),
.B1(n_35),
.B2(n_38),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_50),
.C(n_34),
.Y(n_69)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_0),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_55),
.B1(n_57),
.B2(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_0),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_55),
.B1(n_57),
.B2(n_38),
.Y(n_78)
);

NOR3xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_76),
.C(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_1),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_83),
.B1(n_67),
.B2(n_31),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_57),
.B(n_52),
.Y(n_82)
);

XOR2x1_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_29),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_88),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_90),
.A2(n_76),
.B(n_77),
.C(n_7),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_94),
.Y(n_97)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp67_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_103),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_26),
.C(n_25),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_99),
.C(n_100),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_23),
.C(n_22),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_5),
.B(n_6),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_89),
.B1(n_86),
.B2(n_13),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_20),
.B(n_19),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_104),
.C(n_90),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_9),
.C(n_10),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_10),
.B(n_11),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_109),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_110),
.B(n_112),
.Y(n_116)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_107),
.A2(n_104),
.B(n_96),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_114),
.C(n_110),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_105),
.C(n_12),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_118),
.B1(n_116),
.B2(n_14),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_11),
.C(n_12),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_13),
.C(n_14),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_15),
.C(n_16),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_15),
.B(n_16),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_17),
.Y(n_123)
);


endmodule