module fake_jpeg_19538_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_55),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_15),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_54),
.B(n_75),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_67),
.Y(n_113)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_64),
.Y(n_89)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_18),
.B(n_3),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_71),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_3),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_73),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_19),
.B(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_84),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_19),
.A2(n_4),
.B(n_6),
.Y(n_82)
);

OR2x2_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_6),
.Y(n_124)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_86),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_85),
.A2(n_38),
.B1(n_8),
.B2(n_9),
.Y(n_132)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_14),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_29),
.B1(n_25),
.B2(n_39),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_88),
.A2(n_106),
.B1(n_108),
.B2(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_25),
.B1(n_29),
.B2(n_39),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_91),
.A2(n_109),
.B1(n_112),
.B2(n_117),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_30),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_139),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_45),
.B(n_20),
.C(n_30),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_132),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_29),
.B1(n_37),
.B2(n_36),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_41),
.B1(n_37),
.B2(n_36),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_47),
.A2(n_42),
.B1(n_34),
.B2(n_24),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_52),
.A2(n_33),
.B1(n_41),
.B2(n_22),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_74),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_67),
.A2(n_33),
.B1(n_22),
.B2(n_26),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_62),
.A2(n_30),
.B1(n_34),
.B2(n_42),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_124),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_56),
.A2(n_42),
.B1(n_34),
.B2(n_30),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_78),
.B1(n_64),
.B2(n_69),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_71),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_51),
.B1(n_68),
.B2(n_59),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_SL g136 ( 
.A(n_79),
.B(n_7),
.C(n_9),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_136),
.B(n_10),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_65),
.B1(n_76),
.B2(n_77),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_72),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_10),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_142),
.A2(n_145),
.B1(n_168),
.B2(n_173),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_86),
.B1(n_83),
.B2(n_66),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

NOR2x1_ASAP7_75t_R g149 ( 
.A(n_99),
.B(n_63),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_156),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_100),
.B(n_60),
.Y(n_155)
);

AND2x4_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_45),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_45),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_159),
.Y(n_190)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_132),
.A2(n_75),
.B1(n_57),
.B2(n_50),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_158),
.A2(n_176),
.B1(n_184),
.B2(n_166),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_94),
.B(n_84),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_163),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_58),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_169),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_92),
.B(n_44),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_134),
.Y(n_216)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_164),
.Y(n_221)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_166),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_107),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_60),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_172),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_118),
.B(n_81),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_178),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_113),
.B(n_72),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_103),
.A2(n_53),
.B1(n_72),
.B2(n_13),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_90),
.B(n_11),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_179),
.Y(n_209)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_89),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_103),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_177),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_105),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_128),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_182),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx12_ASAP7_75t_R g183 ( 
.A(n_128),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_133),
.Y(n_213)
);

AND2x2_ASAP7_75t_SL g184 ( 
.A(n_132),
.B(n_93),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_184),
.A2(n_95),
.B(n_133),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_132),
.B1(n_102),
.B2(n_89),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_135),
.B1(n_98),
.B2(n_95),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_110),
.B(n_129),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_96),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_96),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_187),
.B(n_197),
.Y(n_252)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_109),
.B(n_89),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_189),
.A2(n_202),
.B(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_193),
.B(n_215),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_143),
.B(n_104),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_214),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_104),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_147),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_224),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_203),
.B(n_161),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_156),
.B(n_111),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_98),
.C(n_114),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_204),
.A2(n_217),
.B1(n_185),
.B2(n_151),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_157),
.B(n_121),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_114),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_216),
.B(n_162),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_144),
.A2(n_122),
.B1(n_134),
.B2(n_184),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_218),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_147),
.Y(n_224)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_151),
.B(n_122),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_176),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_227),
.B(n_234),
.Y(n_279)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_184),
.B1(n_178),
.B2(n_158),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_230),
.A2(n_255),
.B1(n_189),
.B2(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_231),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_207),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_220),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_151),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_241),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_238),
.A2(n_245),
.B1(n_247),
.B2(n_250),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_239),
.A2(n_258),
.B(n_203),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_171),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_249),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_141),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_211),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_242),
.B(n_246),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_204),
.A2(n_145),
.B1(n_142),
.B2(n_158),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_220),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_158),
.B1(n_159),
.B2(n_140),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_248),
.A2(n_254),
.B(n_257),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_169),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_202),
.A2(n_140),
.B1(n_186),
.B2(n_152),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_202),
.A2(n_173),
.B1(n_150),
.B2(n_176),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_253),
.A2(n_222),
.B1(n_212),
.B2(n_188),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_221),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_205),
.A2(n_181),
.B1(n_176),
.B2(n_160),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_190),
.B(n_176),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_261),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_221),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_199),
.A2(n_163),
.B(n_162),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_259),
.A2(n_216),
.B(n_199),
.Y(n_269)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_201),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_190),
.B(n_175),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_262),
.A2(n_265),
.B1(n_274),
.B2(n_284),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_212),
.C(n_225),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_235),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_189),
.B1(n_188),
.B2(n_222),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_269),
.A2(n_271),
.B(n_280),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_251),
.A2(n_199),
.B(n_215),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_276),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_252),
.B(n_209),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_210),
.C(n_192),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_286),
.C(n_290),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_216),
.B(n_206),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_224),
.C(n_198),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_281),
.B(n_283),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_240),
.B(n_252),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_233),
.A2(n_218),
.B1(n_193),
.B2(n_214),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_241),
.B(n_218),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_256),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_249),
.B(n_218),
.C(n_208),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_233),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_287),
.A2(n_288),
.B1(n_250),
.B2(n_285),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_244),
.A2(n_200),
.B1(n_223),
.B2(n_195),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_232),
.B(n_200),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_292),
.A2(n_306),
.B(n_309),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_235),
.B1(n_238),
.B2(n_253),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_293),
.A2(n_298),
.B1(n_308),
.B2(n_310),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_294),
.B(n_295),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_232),
.B(n_258),
.C(n_259),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_280),
.A2(n_234),
.B1(n_242),
.B2(n_243),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_296),
.A2(n_307),
.B(n_271),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_227),
.Y(n_297)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_297),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_273),
.A2(n_257),
.B1(n_254),
.B2(n_246),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_299),
.A2(n_303),
.B1(n_284),
.B2(n_267),
.Y(n_322)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_287),
.A2(n_231),
.B1(n_229),
.B2(n_228),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_243),
.Y(n_304)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_304),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_286),
.A2(n_236),
.B1(n_183),
.B2(n_165),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_223),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_274),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_195),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_315),
.Y(n_319)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_275),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_313),
.A2(n_317),
.B1(n_273),
.B2(n_170),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_322),
.A2(n_329),
.B1(n_336),
.B2(n_312),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_330),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_282),
.C(n_277),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_327),
.B(n_331),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_310),
.A2(n_267),
.B1(n_290),
.B2(n_278),
.Y(n_329)
);

OAI322xp33_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_283),
.A3(n_276),
.B1(n_282),
.B2(n_272),
.C1(n_269),
.C2(n_278),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_268),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_268),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_333),
.B(n_334),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_201),
.C(n_165),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_291),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_339),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_303),
.A2(n_201),
.B1(n_148),
.B2(n_167),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_148),
.C(n_219),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_337),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_301),
.B(n_154),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_337),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_219),
.C(n_180),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_341),
.A2(n_299),
.B1(n_294),
.B2(n_322),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_297),
.Y(n_342)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_342),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_326),
.A2(n_295),
.B(n_315),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_344),
.A2(n_356),
.B(n_346),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_345),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_347),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_311),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_349),
.B(n_351),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_339),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_352),
.A2(n_329),
.B1(n_318),
.B2(n_308),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_328),
.A2(n_301),
.B(n_296),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_357),
.B(n_335),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_360),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_355),
.B(n_334),
.C(n_327),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_333),
.C(n_331),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_362),
.B(n_370),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_363),
.A2(n_369),
.B1(n_365),
.B2(n_367),
.Y(n_382)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_366),
.Y(n_373)
);

AO221x1_ASAP7_75t_L g368 ( 
.A1(n_349),
.A2(n_332),
.B1(n_325),
.B2(n_306),
.C(n_313),
.Y(n_368)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_368),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_341),
.A2(n_332),
.B1(n_312),
.B2(n_338),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_182),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_371),
.A2(n_356),
.B(n_350),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_375),
.Y(n_387)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_361),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_361),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_376),
.B(n_382),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_350),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_378),
.A2(n_364),
.B(n_342),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_371),
.Y(n_385)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_360),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_381),
.B(n_358),
.Y(n_383)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_383),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_377),
.B(n_370),
.C(n_362),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_390),
.C(n_357),
.Y(n_392)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_385),
.B(n_391),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_372),
.A2(n_351),
.B(n_353),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_386),
.A2(n_348),
.B1(n_344),
.B2(n_366),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_373),
.A2(n_364),
.B1(n_352),
.B2(n_343),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_389),
.A2(n_378),
.B1(n_374),
.B2(n_347),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_379),
.B(n_340),
.C(n_369),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_392),
.B(n_393),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_395),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_388),
.A2(n_348),
.B1(n_167),
.B2(n_146),
.Y(n_395)
);

AOI21xp33_ASAP7_75t_L g398 ( 
.A1(n_396),
.A2(n_387),
.B(n_385),
.Y(n_398)
);

OAI321xp33_ASAP7_75t_L g403 ( 
.A1(n_398),
.A2(n_146),
.A3(n_164),
.B1(n_392),
.B2(n_397),
.C(n_401),
.Y(n_403)
);

A2O1A1O1Ixp25_ASAP7_75t_L g399 ( 
.A1(n_397),
.A2(n_384),
.B(n_390),
.C(n_164),
.D(n_154),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_399),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_403),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_402),
.Y(n_405)
);

AO21x1_ASAP7_75t_L g406 ( 
.A1(n_405),
.A2(n_400),
.B(n_404),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_406),
.Y(n_407)
);


endmodule