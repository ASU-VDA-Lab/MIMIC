module fake_jpeg_24489_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_18),
.Y(n_58)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_32),
.B1(n_27),
.B2(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_62),
.B1(n_31),
.B2(n_20),
.Y(n_77)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_32),
.B1(n_19),
.B2(n_34),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_34),
.B1(n_26),
.B2(n_28),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_21),
.B(n_33),
.C(n_19),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_25),
.B(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_29),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_29),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_65),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_32),
.B1(n_17),
.B2(n_31),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_17),
.Y(n_68)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_78),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_42),
.B1(n_22),
.B2(n_34),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_70),
.A2(n_86),
.B1(n_96),
.B2(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_36),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_24),
.B(n_33),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_82),
.B1(n_94),
.B2(n_100),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_31),
.B1(n_20),
.B2(n_27),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_61),
.B1(n_23),
.B2(n_20),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_24),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_90),
.Y(n_116)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_93),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_92),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_50),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_41),
.B1(n_37),
.B2(n_44),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_26),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_28),
.B1(n_22),
.B2(n_23),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_63),
.B(n_28),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_66),
.A2(n_41),
.B1(n_37),
.B2(n_44),
.Y(n_102)
);

AOI22x1_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_36),
.B1(n_39),
.B2(n_66),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_90),
.B1(n_85),
.B2(n_83),
.Y(n_145)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_113),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_66),
.B1(n_49),
.B2(n_41),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_91),
.B1(n_99),
.B2(n_94),
.Y(n_135)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_89),
.B1(n_84),
.B2(n_44),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_125),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_36),
.Y(n_119)
);

XOR2x1_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_39),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_129),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_88),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_81),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_105),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_71),
.B(n_72),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_148),
.B(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_137),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_87),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_141),
.C(n_144),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_139),
.B1(n_145),
.B2(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_95),
.B1(n_73),
.B2(n_89),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_68),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_111),
.B1(n_124),
.B2(n_104),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_147),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_73),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_117),
.B1(n_126),
.B2(n_127),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_76),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_104),
.A2(n_84),
.B1(n_67),
.B2(n_39),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_150),
.B1(n_124),
.B2(n_109),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_107),
.A2(n_67),
.B1(n_98),
.B2(n_39),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_155),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_98),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_78),
.C(n_69),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_125),
.C(n_103),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_151),
.B(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_164),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_140),
.A2(n_115),
.B(n_111),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_163),
.A2(n_174),
.B(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_172),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_170),
.A2(n_150),
.B1(n_135),
.B2(n_132),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_141),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_107),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_106),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_176),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_106),
.C(n_105),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_16),
.C(n_3),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_179),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_198),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_191),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_183),
.A2(n_194),
.B(n_179),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_139),
.C(n_151),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_196),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_144),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_193),
.C(n_169),
.Y(n_206)
);

OAI322xp33_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_156),
.A3(n_137),
.B1(n_147),
.B2(n_16),
.C1(n_33),
.C2(n_21),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_158),
.C(n_174),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_118),
.B1(n_113),
.B2(n_108),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_157),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_177),
.A2(n_33),
.B(n_3),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_128),
.B1(n_48),
.B2(n_92),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_203),
.B(n_194),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_171),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_206),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_163),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_207),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_160),
.C(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_205),
.C(n_208),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_186),
.C(n_190),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_172),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_168),
.C(n_166),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_159),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_2),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_161),
.C(n_170),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_196),
.C(n_164),
.Y(n_220)
);

OAI31xp33_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_187),
.A3(n_185),
.B(n_183),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_219),
.B(n_221),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_182),
.B1(n_191),
.B2(n_195),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_224),
.B1(n_6),
.B2(n_7),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_8),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_226),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_48),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_2),
.C(n_4),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_10),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_203),
.B(n_2),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_201),
.B1(n_5),
.B2(n_6),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_232),
.C(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_231),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_8),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_10),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_223),
.C(n_214),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_SL g237 ( 
.A(n_234),
.B(n_218),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

OAI221xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_225),
.B1(n_214),
.B2(n_223),
.C(n_14),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_235),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_232),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_246),
.C(n_245),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_229),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_236),
.B1(n_11),
.B2(n_13),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_243),
.B(n_11),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_253),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_250),
.A2(n_10),
.B(n_15),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_15),
.Y(n_255)
);


endmodule