module fake_netlist_6_4762_n_810 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_810);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_810;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

BUFx3_ASAP7_75t_L g183 ( 
.A(n_75),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_67),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_18),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_92),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_16),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_34),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_55),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_60),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_107),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_71),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_56),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_124),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_29),
.Y(n_203)
);

BUFx2_ASAP7_75t_SL g204 ( 
.A(n_43),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_101),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_13),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_141),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_64),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_44),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_58),
.B(n_161),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_84),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_61),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_146),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_40),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_38),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_121),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_140),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_39),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_23),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_12),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_42),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_110),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_85),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_129),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_32),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_37),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_182),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_87),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_27),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_89),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_155),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_6),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_63),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_30),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_2),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_2),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_171),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_68),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_23),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_47),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_8),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_25),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_119),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_41),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_76),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_52),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_112),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_0),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_106),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_131),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_96),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_17),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_18),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_175),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_123),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_148),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_208),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_183),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_225),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_183),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_225),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_206),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_186),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_193),
.B(n_5),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_209),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_193),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_189),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_190),
.A2(n_7),
.B(n_8),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_208),
.B(n_26),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_211),
.B(n_28),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_31),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_248),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_195),
.B(n_9),
.Y(n_299)
);

BUFx12f_ASAP7_75t_L g300 ( 
.A(n_191),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_187),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_264),
.Y(n_303)
);

AND2x6_ASAP7_75t_L g304 ( 
.A(n_236),
.B(n_181),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_246),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_236),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_184),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_185),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_188),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_192),
.B(n_11),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_196),
.B(n_33),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_199),
.B(n_35),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_200),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_203),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_205),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g317 ( 
.A1(n_213),
.A2(n_13),
.B(n_14),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_194),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_214),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_219),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_267),
.B(n_187),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_267),
.B(n_235),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_289),
.Y(n_325)
);

NOR2x1p5_ASAP7_75t_L g326 ( 
.A(n_285),
.B(n_197),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_221),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_270),
.B(n_226),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_283),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_285),
.B(n_235),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g332 ( 
.A(n_265),
.B(n_211),
.C(n_201),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_298),
.B(n_262),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_309),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_298),
.B(n_262),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_307),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_280),
.B(n_237),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_307),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_230),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_287),
.B(n_198),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

NAND3x1_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_250),
.C(n_231),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_300),
.Y(n_348)
);

AND3x2_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_254),
.C(n_232),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_270),
.B(n_233),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_288),
.A2(n_228),
.B1(n_216),
.B2(n_223),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_287),
.B(n_202),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_238),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_297),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_283),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_297),
.Y(n_358)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_296),
.B(n_259),
.C(n_207),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_270),
.B(n_210),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_297),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_312),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_272),
.B(n_312),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_L g365 ( 
.A(n_304),
.B(n_212),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_288),
.A2(n_204),
.B1(n_247),
.B2(n_258),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_271),
.B(n_240),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_282),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_272),
.B(n_271),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_272),
.B(n_244),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_245),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_313),
.Y(n_374)
);

OR2x6_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_276),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_313),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_279),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_288),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_368),
.B(n_300),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_303),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_342),
.B(n_318),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_351),
.B(n_318),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_324),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_303),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_347),
.A2(n_277),
.B1(n_291),
.B2(n_354),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_371),
.B(n_215),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_330),
.B(n_308),
.Y(n_388)
);

A2O1A1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_373),
.A2(n_317),
.B(n_314),
.C(n_320),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_327),
.A2(n_286),
.B1(n_317),
.B2(n_308),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_328),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_L g393 ( 
.A(n_332),
.B(n_304),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_306),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_330),
.B(n_217),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_366),
.B(n_303),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_303),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_324),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_306),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_327),
.A2(n_286),
.B1(n_314),
.B2(n_320),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_327),
.Y(n_402)
);

O2A1O1Ixp5_ASAP7_75t_L g403 ( 
.A1(n_343),
.A2(n_314),
.B(n_316),
.C(n_315),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_336),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_303),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_353),
.B(n_303),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_322),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_357),
.B(n_319),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_359),
.B(n_344),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_326),
.A2(n_269),
.B1(n_220),
.B2(n_222),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_331),
.B(n_218),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_356),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_338),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_333),
.B(n_319),
.Y(n_417)
);

OR2x6_ASAP7_75t_L g418 ( 
.A(n_335),
.B(n_323),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_338),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_341),
.B(n_310),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_324),
.Y(n_421)
);

NAND2x1p5_ASAP7_75t_L g422 ( 
.A(n_340),
.B(n_286),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_L g423 ( 
.A(n_370),
.B(n_257),
.C(n_284),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_334),
.B(n_310),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_337),
.B(n_315),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_365),
.A2(n_316),
.B(n_305),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_341),
.Y(n_427)
);

OR2x6_ASAP7_75t_L g428 ( 
.A(n_329),
.B(n_279),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_345),
.B(n_227),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_345),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_346),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

A2O1A1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_350),
.A2(n_305),
.B(n_273),
.C(n_301),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_352),
.B(n_229),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_355),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_355),
.B(n_358),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_361),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_361),
.B(n_234),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_402),
.A2(n_365),
.B(n_340),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_399),
.Y(n_442)
);

O2A1O1Ixp33_ASAP7_75t_L g443 ( 
.A1(n_378),
.A2(n_372),
.B(n_294),
.C(n_284),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_374),
.B(n_349),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_367),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_408),
.A2(n_340),
.B1(n_251),
.B2(n_253),
.Y(n_446)
);

BUFx4f_ASAP7_75t_L g447 ( 
.A(n_418),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_381),
.A2(n_367),
.B(n_325),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_405),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_367),
.Y(n_451)
);

NAND2x1p5_ASAP7_75t_L g452 ( 
.A(n_377),
.B(n_286),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_385),
.A2(n_325),
.B(n_362),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_422),
.A2(n_362),
.B(n_304),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_325),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_376),
.B(n_325),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_376),
.B(n_325),
.Y(n_458)
);

AO21x1_ASAP7_75t_L g459 ( 
.A1(n_393),
.A2(n_273),
.B(n_281),
.Y(n_459)
);

NOR3xp33_ASAP7_75t_L g460 ( 
.A(n_379),
.B(n_348),
.C(n_294),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_396),
.A2(n_281),
.B(n_292),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_394),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_397),
.A2(n_292),
.B(n_293),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_382),
.B(n_348),
.Y(n_464)
);

O2A1O1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_433),
.A2(n_295),
.B(n_278),
.C(n_266),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_376),
.B(n_304),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_387),
.B(n_241),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_376),
.B(n_304),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_409),
.B(n_295),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_380),
.B(n_304),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_419),
.A2(n_301),
.B(n_293),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_391),
.B(n_290),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_390),
.A2(n_418),
.B1(n_428),
.B2(n_401),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_429),
.A2(n_278),
.B(n_274),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_435),
.A2(n_274),
.B(n_268),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

NOR2x1p5_ASAP7_75t_L g477 ( 
.A(n_406),
.B(n_266),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_418),
.A2(n_268),
.B1(n_290),
.B2(n_108),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_440),
.A2(n_290),
.B(n_105),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_386),
.A2(n_290),
.B1(n_104),
.B2(n_109),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_392),
.B(n_404),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_415),
.B(n_290),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_413),
.B(n_14),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_428),
.B(n_426),
.Y(n_484)
);

CKINVDCx6p67_ASAP7_75t_R g485 ( 
.A(n_375),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_386),
.A2(n_290),
.B1(n_111),
.B2(n_113),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_437),
.A2(n_407),
.B(n_420),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_436),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_403),
.A2(n_99),
.B(n_176),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_411),
.A2(n_97),
.B(n_174),
.Y(n_490)
);

INVx8_ASAP7_75t_L g491 ( 
.A(n_375),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_375),
.B(n_15),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_427),
.A2(n_95),
.B(n_173),
.Y(n_493)
);

AO22x1_ASAP7_75t_L g494 ( 
.A1(n_423),
.A2(n_412),
.B1(n_425),
.B2(n_424),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_416),
.A2(n_94),
.B(n_172),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_430),
.Y(n_496)
);

O2A1O1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_389),
.A2(n_15),
.B(n_17),
.C(n_19),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_410),
.B(n_19),
.Y(n_498)
);

OAI321xp33_ASAP7_75t_L g499 ( 
.A1(n_383),
.A2(n_20),
.A3(n_21),
.B1(n_22),
.B2(n_24),
.C(n_25),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_439),
.A2(n_114),
.B(n_168),
.Y(n_500)
);

AO21x1_ASAP7_75t_L g501 ( 
.A1(n_431),
.A2(n_20),
.B(n_21),
.Y(n_501)
);

NAND3xp33_ASAP7_75t_L g502 ( 
.A(n_434),
.B(n_115),
.C(n_167),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_438),
.A2(n_100),
.B(n_166),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_395),
.B(n_22),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_384),
.A2(n_117),
.B1(n_36),
.B2(n_45),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_384),
.Y(n_506)
);

A2O1A1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_398),
.A2(n_421),
.B(n_414),
.C(n_24),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_421),
.A2(n_46),
.B(n_48),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_398),
.B(n_49),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_492),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_445),
.A2(n_421),
.B(n_414),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_450),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_448),
.A2(n_54),
.B(n_57),
.Y(n_513)
);

AO31x2_ASAP7_75t_L g514 ( 
.A1(n_459),
.A2(n_59),
.A3(n_62),
.B(n_65),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_469),
.B(n_66),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_473),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_484),
.A2(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_455),
.B(n_78),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_441),
.A2(n_79),
.B(n_80),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_461),
.A2(n_180),
.B(n_82),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_487),
.A2(n_165),
.B(n_83),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_476),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_481),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_462),
.B(n_81),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_451),
.A2(n_86),
.B(n_88),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_464),
.B(n_90),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_449),
.B(n_91),
.Y(n_527)
);

AO32x2_ASAP7_75t_L g528 ( 
.A1(n_478),
.A2(n_480),
.A3(n_446),
.B1(n_499),
.B2(n_497),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_496),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_457),
.A2(n_93),
.B(n_118),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_458),
.A2(n_120),
.B(n_122),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_454),
.A2(n_125),
.B(n_126),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_443),
.A2(n_127),
.B(n_128),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_483),
.A2(n_130),
.B(n_132),
.C(n_133),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_456),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_466),
.A2(n_134),
.B(n_135),
.Y(n_536)
);

CKINVDCx6p67_ASAP7_75t_R g537 ( 
.A(n_485),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_452),
.A2(n_136),
.B(n_137),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_491),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_468),
.A2(n_138),
.B(n_139),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_476),
.Y(n_541)
);

AO31x2_ASAP7_75t_L g542 ( 
.A1(n_501),
.A2(n_143),
.A3(n_144),
.B(n_145),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_467),
.B(n_147),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_494),
.B(n_149),
.Y(n_544)
);

AOI211x1_ASAP7_75t_L g545 ( 
.A1(n_498),
.A2(n_150),
.B(n_154),
.C(n_157),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_442),
.B(n_158),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_447),
.B(n_159),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_488),
.B(n_160),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_491),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_488),
.Y(n_550)
);

OAI21xp33_ASAP7_75t_L g551 ( 
.A1(n_460),
.A2(n_162),
.B(n_163),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_506),
.Y(n_552)
);

NOR2xp67_ASAP7_75t_L g553 ( 
.A(n_444),
.B(n_486),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_453),
.A2(n_470),
.B(n_472),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_452),
.A2(n_482),
.B(n_463),
.Y(n_555)
);

AO21x1_ASAP7_75t_L g556 ( 
.A1(n_503),
.A2(n_509),
.B(n_504),
.Y(n_556)
);

NAND3xp33_ASAP7_75t_SL g557 ( 
.A(n_505),
.B(n_507),
.C(n_489),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_506),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_471),
.A2(n_465),
.B(n_479),
.Y(n_559)
);

OA22x2_ASAP7_75t_L g560 ( 
.A1(n_447),
.A2(n_491),
.B1(n_477),
.B2(n_502),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_490),
.A2(n_493),
.B(n_495),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_500),
.A2(n_474),
.B(n_475),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_456),
.A2(n_502),
.B(n_508),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_456),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_473),
.A2(n_368),
.B1(n_378),
.B2(n_351),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_469),
.B(n_368),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_541),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_523),
.B(n_566),
.Y(n_568)
);

CKINVDCx8_ASAP7_75t_R g569 ( 
.A(n_549),
.Y(n_569)
);

NOR2xp67_ASAP7_75t_SL g570 ( 
.A(n_533),
.B(n_543),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_527),
.B(n_553),
.Y(n_571)
);

OA21x2_ASAP7_75t_L g572 ( 
.A1(n_511),
.A2(n_521),
.B(n_538),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_565),
.B(n_529),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_539),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_529),
.B(n_515),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_554),
.A2(n_561),
.B(n_520),
.Y(n_576)
);

AOI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_510),
.A2(n_560),
.B(n_524),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_527),
.B(n_546),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_541),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_564),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_512),
.B(n_528),
.Y(n_581)
);

INVx6_ASAP7_75t_L g582 ( 
.A(n_535),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_512),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_544),
.A2(n_510),
.B1(n_522),
.B2(n_550),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_558),
.B(n_552),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_537),
.B(n_558),
.Y(n_586)
);

INVx8_ASAP7_75t_L g587 ( 
.A(n_535),
.Y(n_587)
);

AO31x2_ASAP7_75t_L g588 ( 
.A1(n_556),
.A2(n_516),
.A3(n_563),
.B(n_534),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_545),
.A2(n_518),
.B1(n_535),
.B2(n_517),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_559),
.A2(n_532),
.B(n_555),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_548),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_526),
.B(n_551),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_513),
.B(n_519),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_562),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_528),
.B(n_547),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_557),
.A2(n_525),
.B(n_540),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_536),
.A2(n_530),
.B(n_531),
.Y(n_597)
);

AOI22x1_ASAP7_75t_L g598 ( 
.A1(n_528),
.A2(n_563),
.B1(n_533),
.B2(n_477),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_542),
.B(n_514),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_514),
.A2(n_554),
.B(n_461),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_542),
.B(n_514),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_542),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_529),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_566),
.A2(n_368),
.B1(n_565),
.B2(n_351),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_541),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_564),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_554),
.A2(n_461),
.B(n_561),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_523),
.B(n_566),
.Y(n_608)
);

OAI21x1_ASAP7_75t_L g609 ( 
.A1(n_554),
.A2(n_461),
.B(n_561),
.Y(n_609)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_554),
.A2(n_461),
.B(n_561),
.Y(n_610)
);

BUFx2_ASAP7_75t_SL g611 ( 
.A(n_539),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_608),
.B(n_568),
.Y(n_612)
);

OA21x2_ASAP7_75t_L g613 ( 
.A1(n_600),
.A2(n_602),
.B(n_599),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_567),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_587),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_571),
.B(n_578),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_583),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_583),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_567),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_604),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_580),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_595),
.B(n_578),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_595),
.B(n_573),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_571),
.B(n_579),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_571),
.B(n_605),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_603),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_581),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_581),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_587),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_580),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_575),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_587),
.Y(n_632)
);

OAI22xp33_ASAP7_75t_L g633 ( 
.A1(n_592),
.A2(n_577),
.B1(n_569),
.B2(n_606),
.Y(n_633)
);

NAND2x1p5_ASAP7_75t_L g634 ( 
.A(n_593),
.B(n_570),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_584),
.B(n_588),
.Y(n_635)
);

OAI222xp33_ASAP7_75t_L g636 ( 
.A1(n_598),
.A2(n_570),
.B1(n_589),
.B2(n_569),
.C1(n_574),
.C2(n_591),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_587),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_582),
.Y(n_638)
);

NOR2x1_ASAP7_75t_SL g639 ( 
.A(n_602),
.B(n_594),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_582),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_585),
.B(n_588),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_585),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_585),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_601),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_596),
.A2(n_611),
.B1(n_601),
.B2(n_582),
.Y(n_645)
);

AO21x2_ASAP7_75t_L g646 ( 
.A1(n_576),
.A2(n_590),
.B(n_600),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_588),
.B(n_586),
.Y(n_647)
);

NOR2x1_ASAP7_75t_L g648 ( 
.A(n_636),
.B(n_601),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_622),
.B(n_588),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_624),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_615),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_623),
.B(n_588),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_622),
.B(n_572),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_624),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_623),
.B(n_572),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_631),
.B(n_572),
.Y(n_656)
);

CKINVDCx8_ASAP7_75t_R g657 ( 
.A(n_629),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_625),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_631),
.B(n_593),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_615),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_612),
.B(n_620),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_647),
.B(n_590),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_617),
.B(n_593),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_613),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_613),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_627),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_615),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_625),
.B(n_582),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_635),
.B(n_607),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_616),
.B(n_609),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_613),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_617),
.B(n_597),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_621),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_628),
.B(n_610),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_644),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_618),
.B(n_614),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_634),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_626),
.A2(n_645),
.B1(n_633),
.B2(n_635),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_616),
.B(n_642),
.Y(n_679)
);

NOR2x1_ASAP7_75t_SL g680 ( 
.A(n_644),
.B(n_646),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_618),
.B(n_619),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_664),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_677),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_649),
.B(n_641),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_661),
.B(n_626),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_650),
.B(n_616),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_649),
.B(n_641),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_655),
.B(n_641),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_655),
.B(n_641),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_652),
.B(n_646),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_654),
.B(n_658),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_664),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_653),
.B(n_642),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_653),
.B(n_643),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_679),
.B(n_643),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_665),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_652),
.B(n_634),
.Y(n_697)
);

OR2x6_ASAP7_75t_L g698 ( 
.A(n_677),
.B(n_634),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_656),
.B(n_639),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_656),
.B(n_639),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_668),
.B(n_630),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_651),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_675),
.B(n_646),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_676),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_651),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_662),
.B(n_638),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_670),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_672),
.A2(n_632),
.B(n_638),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_675),
.B(n_640),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_679),
.B(n_638),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_662),
.B(n_669),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_666),
.B(n_640),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_651),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_701),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_711),
.B(n_690),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_682),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_684),
.B(n_674),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_684),
.B(n_674),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_691),
.B(n_685),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_682),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_687),
.B(n_669),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_692),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_692),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_687),
.B(n_680),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_697),
.B(n_680),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_693),
.B(n_659),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_693),
.B(n_659),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_697),
.B(n_671),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_704),
.B(n_678),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_707),
.B(n_677),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_688),
.B(n_689),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_688),
.B(n_671),
.Y(n_732)
);

AND2x4_ASAP7_75t_L g733 ( 
.A(n_707),
.B(n_677),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_711),
.B(n_690),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_708),
.B(n_648),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_698),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_715),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_715),
.B(n_706),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_734),
.Y(n_739)
);

OAI21xp33_ASAP7_75t_L g740 ( 
.A1(n_735),
.A2(n_648),
.B(n_709),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_720),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_731),
.B(n_700),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_730),
.B(n_699),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_730),
.B(n_699),
.Y(n_744)
);

NOR2x1p5_ASAP7_75t_L g745 ( 
.A(n_729),
.B(n_710),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_734),
.B(n_703),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_720),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_719),
.B(n_703),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_714),
.B(n_700),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_722),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_731),
.B(n_694),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_722),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_723),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_728),
.B(n_696),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_716),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_749),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_741),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_739),
.B(n_732),
.Y(n_758)
);

OAI32xp33_ASAP7_75t_L g759 ( 
.A1(n_740),
.A2(n_724),
.A3(n_736),
.B1(n_726),
.B2(n_727),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_747),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_748),
.B(n_721),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_750),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_742),
.B(n_739),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_748),
.A2(n_686),
.B1(n_736),
.B2(n_698),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_752),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_753),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_738),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_756),
.B(n_737),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_761),
.A2(n_745),
.B1(n_746),
.B2(n_743),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_767),
.B(n_751),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_759),
.A2(n_698),
.B(n_746),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_758),
.A2(n_743),
.B1(n_744),
.B2(n_725),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_SL g773 ( 
.A(n_771),
.B(n_758),
.C(n_763),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_769),
.A2(n_764),
.B1(n_744),
.B2(n_733),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_768),
.B(n_766),
.C(n_765),
.Y(n_775)
);

AOI221xp5_ASAP7_75t_L g776 ( 
.A1(n_772),
.A2(n_762),
.B1(n_760),
.B2(n_673),
.C(n_757),
.Y(n_776)
);

OAI21xp5_ASAP7_75t_L g777 ( 
.A1(n_770),
.A2(n_757),
.B(n_755),
.Y(n_777)
);

NAND4xp75_ASAP7_75t_L g778 ( 
.A(n_774),
.B(n_776),
.C(n_777),
.D(n_773),
.Y(n_778)
);

NOR3xp33_ASAP7_75t_L g779 ( 
.A(n_775),
.B(n_667),
.C(n_712),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_775),
.Y(n_780)
);

NAND4xp75_ASAP7_75t_L g781 ( 
.A(n_780),
.B(n_712),
.C(n_667),
.D(n_702),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_779),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_782),
.B(n_778),
.Y(n_783)
);

NOR2x1_ASAP7_75t_L g784 ( 
.A(n_781),
.B(n_660),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_783),
.B(n_754),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_784),
.B(n_660),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_784),
.Y(n_787)
);

INVx4_ASAP7_75t_L g788 ( 
.A(n_787),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_785),
.A2(n_695),
.B1(n_713),
.B2(n_705),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_786),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_789),
.A2(n_657),
.B1(n_733),
.B2(n_730),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_788),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_790),
.B(n_638),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_792),
.B(n_790),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_793),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_791),
.B(n_718),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_792),
.A2(n_629),
.B(n_637),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_794),
.A2(n_629),
.B(n_637),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_795),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_796),
.A2(n_695),
.B1(n_683),
.B2(n_637),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_797),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_794),
.A2(n_637),
.B(n_681),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_794),
.B(n_637),
.Y(n_803)
);

NAND2x1_ASAP7_75t_L g804 ( 
.A(n_799),
.B(n_640),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_803),
.A2(n_640),
.B(n_663),
.Y(n_805)
);

OR4x2_ASAP7_75t_L g806 ( 
.A(n_801),
.B(n_717),
.C(n_695),
.D(n_721),
.Y(n_806)
);

AO21x2_ASAP7_75t_L g807 ( 
.A1(n_805),
.A2(n_798),
.B(n_802),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_804),
.B(n_800),
.Y(n_808)
);

XOR2xp5_ASAP7_75t_L g809 ( 
.A(n_808),
.B(n_806),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_809),
.A2(n_807),
.B1(n_670),
.B2(n_694),
.Y(n_810)
);


endmodule