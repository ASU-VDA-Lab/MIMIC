module fake_jpeg_3249_n_214 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_214);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_214;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_1),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_78),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_63),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_86),
.B(n_90),
.C(n_82),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_63),
.B1(n_60),
.B2(n_67),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_78),
.B1(n_76),
.B2(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_56),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_79),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_58),
.B1(n_67),
.B2(n_59),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_91),
.B1(n_72),
.B2(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_62),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_95),
.Y(n_124)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_72),
.B1(n_88),
.B2(n_70),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_71),
.B(n_70),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_52),
.B(n_65),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_109),
.Y(n_126)
);

OA22x2_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_72),
.B1(n_53),
.B2(n_58),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_106),
.Y(n_112)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_71),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_81),
.B1(n_86),
.B2(n_51),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_121),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_68),
.B1(n_52),
.B2(n_51),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_8),
.B(n_9),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_2),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_53),
.B1(n_64),
.B2(n_55),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_53),
.B1(n_64),
.B2(n_4),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_23),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_127),
.C(n_128),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_50),
.B1(n_49),
.B2(n_48),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_47),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_46),
.Y(n_139)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_136),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_94),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_147),
.C(n_152),
.Y(n_158)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_141),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_98),
.B(n_5),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_12),
.B(n_13),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_142),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_6),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_SL g145 ( 
.A(n_110),
.B(n_7),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_118),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_39),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_128),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_151),
.B(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_10),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_150),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_12),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_35),
.B1(n_33),
.B2(n_32),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_152),
.B(n_14),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_158),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_170),
.Y(n_176)
);

AOI22x1_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_131),
.B1(n_125),
.B2(n_30),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_SL g185 ( 
.A1(n_160),
.A2(n_163),
.B(n_16),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_161),
.B(n_171),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_28),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_167),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_27),
.B(n_26),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_145),
.B1(n_151),
.B2(n_18),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_25),
.C(n_24),
.Y(n_170)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_153),
.A2(n_159),
.B(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_180),
.Y(n_194)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_146),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_182),
.Y(n_195)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_185),
.C(n_163),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_162),
.C(n_170),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_190),
.C(n_181),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_189),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_177),
.B(n_166),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_194),
.B(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_200),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_199),
.C(n_191),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_192),
.A2(n_173),
.B(n_157),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_173),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_17),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_185),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_191),
.B1(n_193),
.B2(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_203),
.B(n_205),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

OAI321xp33_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_206),
.A3(n_196),
.B1(n_200),
.B2(n_20),
.C(n_17),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_207),
.B1(n_19),
.B2(n_20),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_22),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_18),
.C(n_21),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_21),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_22),
.Y(n_214)
);


endmodule