module fake_jpeg_26104_n_342 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_54),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_43),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_51),
.Y(n_73)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_26),
.B1(n_32),
.B2(n_22),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_47),
.B1(n_32),
.B2(n_22),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_72),
.A2(n_87),
.B1(n_91),
.B2(n_99),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_74),
.B(n_83),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_47),
.B1(n_32),
.B2(n_38),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_26),
.B1(n_32),
.B2(n_24),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_26),
.B1(n_20),
.B2(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_90),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g81 ( 
.A(n_56),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_26),
.B1(n_20),
.B2(n_21),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_95),
.B1(n_100),
.B2(n_25),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_41),
.B1(n_39),
.B2(n_48),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_49),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_28),
.B(n_35),
.Y(n_109)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_20),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_94),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_61),
.A2(n_23),
.B1(n_21),
.B2(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_23),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_17),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_40),
.B1(n_17),
.B2(n_35),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_21),
.B1(n_35),
.B2(n_17),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_18),
.C(n_25),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_101),
.B(n_72),
.CI(n_94),
.CON(n_147),
.SN(n_147)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_126),
.Y(n_145)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_112),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_98),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_64),
.B1(n_28),
.B2(n_30),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_143)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_62),
.C(n_68),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_25),
.B1(n_30),
.B2(n_28),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_30),
.B1(n_68),
.B2(n_36),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_80),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_73),
.B1(n_85),
.B2(n_82),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_93),
.Y(n_129)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_133),
.Y(n_168)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_97),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_149),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_90),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_141),
.Y(n_165)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_140),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_148),
.B(n_125),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_77),
.Y(n_141)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_73),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_122),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_74),
.B(n_99),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_25),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_154),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_75),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_73),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_156),
.A2(n_85),
.B(n_126),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_25),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_159),
.B(n_173),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_135),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_125),
.B(n_113),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_142),
.B1(n_153),
.B2(n_155),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_131),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_182),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_151),
.B1(n_148),
.B2(n_152),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_84),
.B1(n_25),
.B2(n_34),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_103),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_113),
.B1(n_118),
.B2(n_123),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_176),
.B1(n_185),
.B2(n_139),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_175),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_130),
.A2(n_123),
.B1(n_85),
.B2(n_116),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_SL g193 ( 
.A1(n_177),
.A2(n_180),
.B(n_147),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_70),
.C(n_114),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_186),
.C(n_27),
.Y(n_221)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_138),
.B(n_70),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_188),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_82),
.Y(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_145),
.A2(n_116),
.B1(n_82),
.B2(n_84),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_70),
.C(n_62),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_27),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_70),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_25),
.Y(n_202)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_139),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_196),
.Y(n_228)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_194),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_195),
.A2(n_200),
.B1(n_163),
.B2(n_1),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_166),
.B(n_176),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_133),
.Y(n_199)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_221),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_153),
.B1(n_137),
.B2(n_84),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_209),
.B1(n_172),
.B2(n_181),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_206),
.A2(n_163),
.B1(n_181),
.B2(n_18),
.Y(n_239)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_215),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_174),
.B1(n_170),
.B2(n_179),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_160),
.B(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_62),
.Y(n_213)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g216 ( 
.A1(n_164),
.A2(n_27),
.A3(n_18),
.B1(n_10),
.B2(n_11),
.Y(n_216)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_159),
.B(n_18),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_178),
.Y(n_230)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_220),
.Y(n_231)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_161),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_167),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_0),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_226),
.A2(n_240),
.B(n_245),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_222),
.B1(n_219),
.B2(n_197),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_234),
.Y(n_263)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_183),
.C(n_161),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_246),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_177),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_186),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_236),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_190),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_239),
.A2(n_205),
.B1(n_247),
.B2(n_208),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_8),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_243),
.C(n_194),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_9),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_9),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_9),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_223),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_249),
.B(n_251),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_250),
.A2(n_211),
.B1(n_232),
.B2(n_224),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_222),
.B(n_203),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_237),
.Y(n_252)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_230),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_256),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_202),
.C(n_194),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_262),
.C(n_234),
.Y(n_277)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_229),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_195),
.C(n_206),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_207),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_270),
.B1(n_7),
.B2(n_14),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_241),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_269),
.B(n_208),
.Y(n_285)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_266),
.B1(n_250),
.B2(n_251),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_272),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_284),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_288),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_235),
.C(n_236),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_280),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_238),
.C(n_241),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_216),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_285),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_211),
.C(n_11),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_286),
.B(n_287),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_7),
.C(n_14),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_260),
.B1(n_256),
.B2(n_267),
.Y(n_289)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_272),
.B(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_264),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_300),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_298),
.A2(n_286),
.B1(n_271),
.B2(n_284),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_270),
.B(n_259),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_299),
.A2(n_281),
.B(n_275),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_262),
.B1(n_253),
.B2(n_11),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_5),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_303),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_277),
.B(n_5),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_302),
.B(n_12),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_5),
.Y(n_303)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_290),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_305),
.B(n_309),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_280),
.C(n_287),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_311),
.C(n_312),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_282),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_0),
.B(n_1),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_291),
.A2(n_12),
.B1(n_13),
.B2(n_16),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_12),
.C(n_13),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_16),
.B1(n_1),
.B2(n_2),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_13),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_16),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_315),
.A2(n_302),
.B(n_301),
.Y(n_318)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_318),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_294),
.C(n_303),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_294),
.C(n_298),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_323),
.B(n_310),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_324),
.C(n_314),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_325),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_331),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_304),
.C(n_312),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_324),
.A2(n_308),
.B(n_2),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_332),
.B(n_308),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_326),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_336),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_333),
.B(n_335),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_328),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_0),
.C(n_2),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_340),
.B(n_0),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_4),
.Y(n_342)
);


endmodule