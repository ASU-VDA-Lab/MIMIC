module real_jpeg_9281_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_1),
.A2(n_21),
.B1(n_22),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_2),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_8),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_9),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_9),
.A2(n_21),
.B1(n_22),
.B2(n_45),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_10),
.A2(n_21),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_10),
.B(n_21),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_56),
.B1(n_93),
.B2(n_94),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_72),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_71),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_63),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_49),
.B2(n_62),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_20),
.A2(n_25),
.B1(n_28),
.B2(n_67),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_26),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_21),
.A2(n_22),
.B1(n_40),
.B2(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_21),
.B(n_40),
.Y(n_51)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_22),
.A2(n_36),
.B1(n_42),
.B2(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_25),
.A2(n_28),
.B1(n_67),
.B2(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_28),
.B(n_38),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_29),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_29),
.B(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_29),
.B(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_30),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_38),
.CON(n_36),
.SN(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_40),
.Y(n_42)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_38),
.B(n_94),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_56),
.B(n_59),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_58),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_69),
.B(n_70),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_77),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_58),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_58),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_63),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.CI(n_68),
.CON(n_63),
.SN(n_63)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_101),
.B(n_104),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_89),
.B(n_100),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_88),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_88),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_83),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_95),
.B(n_99),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);


endmodule