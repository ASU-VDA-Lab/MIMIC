module fake_jpeg_6353_n_11 (n_3, n_2, n_1, n_0, n_4, n_11);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_11;

wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

NOR2xp33_ASAP7_75t_SL g5 ( 
.A(n_0),
.B(n_1),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_0),
.Y(n_6)
);

A2O1A1O1Ixp25_ASAP7_75t_L g7 ( 
.A1(n_6),
.A2(n_0),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_7)
);

MAJIxp5_ASAP7_75t_L g8 ( 
.A(n_7),
.B(n_5),
.C(n_2),
.Y(n_8)
);

MAJIxp5_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_5),
.C(n_4),
.Y(n_9)
);

OAI21xp5_ASAP7_75t_SL g10 ( 
.A1(n_9),
.A2(n_4),
.B(n_1),
.Y(n_10)
);

NOR3xp33_ASAP7_75t_SL g11 ( 
.A(n_10),
.B(n_3),
.C(n_7),
.Y(n_11)
);


endmodule