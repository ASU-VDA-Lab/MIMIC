module fake_jpeg_14695_n_47 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_47);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_47;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_32;

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_6),
.B(n_9),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_17),
.B1(n_19),
.B2(n_3),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_19),
.B1(n_22),
.B2(n_20),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_18),
.B1(n_20),
.B2(n_4),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_22),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_33),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_17),
.C(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_27),
.B1(n_2),
.B2(n_4),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_32),
.A2(n_18),
.B1(n_5),
.B2(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_38),
.B(n_7),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_8),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_29),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B(n_10),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_40),
.A3(n_41),
.B1(n_24),
.B2(n_13),
.Y(n_47)
);


endmodule