module fake_aes_11785_n_671 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_671);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_671;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_17), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_66), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_1), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_20), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_60), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_16), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_34), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_22), .Y(n_83) );
INVxp33_ASAP7_75t_SL g84 ( .A(n_53), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_14), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_50), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_56), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_36), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_3), .Y(n_89) );
CKINVDCx14_ASAP7_75t_R g90 ( .A(n_63), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_59), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_55), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_38), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_47), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_52), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_61), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_12), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_45), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_28), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_8), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_26), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
BUFx3_ASAP7_75t_L g103 ( .A(n_24), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_35), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_7), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_7), .Y(n_106) );
INVxp33_ASAP7_75t_SL g107 ( .A(n_6), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_51), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_62), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_18), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_32), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_10), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_48), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_21), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_49), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_43), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_64), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_12), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_13), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_54), .Y(n_122) );
AND3x2_ASAP7_75t_L g123 ( .A(n_89), .B(n_0), .C(n_1), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_99), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_89), .B(n_121), .Y(n_126) );
AND2x6_ASAP7_75t_L g127 ( .A(n_103), .B(n_29), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
CKINVDCx6p67_ASAP7_75t_R g129 ( .A(n_87), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_107), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_108), .B(n_2), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_77), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
CKINVDCx16_ASAP7_75t_R g139 ( .A(n_90), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_121), .B(n_4), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_76), .B(n_5), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_103), .Y(n_143) );
NOR3xp33_ASAP7_75t_L g144 ( .A(n_81), .B(n_5), .C(n_6), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_83), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
BUFx2_ASAP7_75t_L g148 ( .A(n_76), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_86), .B(n_8), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_88), .Y(n_150) );
OR2x6_ASAP7_75t_L g151 ( .A(n_78), .B(n_9), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_88), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
CKINVDCx6p67_ASAP7_75t_R g154 ( .A(n_91), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_92), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_97), .B(n_100), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_85), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_116), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_116), .B(n_9), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_119), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_119), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_122), .B(n_10), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_148), .B(n_120), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
AND2x2_ASAP7_75t_L g166 ( .A(n_148), .B(n_120), .Y(n_166) );
AO22x2_ASAP7_75t_L g167 ( .A1(n_149), .A2(n_106), .B1(n_112), .B2(n_115), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_126), .B(n_102), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_124), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_127), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_124), .Y(n_172) );
NOR2xp33_ASAP7_75t_SL g173 ( .A(n_129), .B(n_104), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_137), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_139), .B(n_84), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_139), .B(n_84), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_129), .B(n_118), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_129), .B(n_117), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_124), .Y(n_181) );
INVx4_ASAP7_75t_L g182 ( .A(n_127), .Y(n_182) );
BUFx10_ASAP7_75t_L g183 ( .A(n_126), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_156), .B(n_114), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_132), .B(n_107), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_124), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_158), .B(n_113), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_132), .B(n_98), .Y(n_188) );
NAND3xp33_ASAP7_75t_L g189 ( .A(n_134), .B(n_111), .C(n_93), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_124), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_124), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_126), .B(n_109), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_126), .B(n_94), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_127), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_146), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_134), .B(n_101), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_146), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_143), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_136), .B(n_96), .Y(n_200) );
INVx1_ASAP7_75t_SL g201 ( .A(n_133), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_141), .B(n_95), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_125), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_125), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_149), .B(n_40), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_152), .Y(n_207) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_163), .A2(n_41), .B(n_75), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_125), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_136), .B(n_110), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_149), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_127), .Y(n_212) );
INVx3_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_160), .B(n_11), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_138), .B(n_105), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_152), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_160), .B(n_11), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_160), .B(n_13), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_135), .B(n_14), .Y(n_219) );
AO22x2_ASAP7_75t_L g220 ( .A1(n_144), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_151), .A2(n_15), .B1(n_18), .B2(n_19), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_135), .B(n_19), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_164), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_183), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
AND3x2_ASAP7_75t_SL g226 ( .A(n_173), .B(n_154), .C(n_151), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_167), .A2(n_151), .B1(n_133), .B2(n_141), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_185), .B(n_157), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_167), .A2(n_151), .B1(n_140), .B2(n_130), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_183), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_183), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_219), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_164), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_219), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_196), .B(n_140), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_219), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_167), .A2(n_130), .B1(n_161), .B2(n_147), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_179), .B(n_157), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_171), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_199), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_179), .B(n_123), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_222), .Y(n_243) );
INVx5_ASAP7_75t_L g244 ( .A(n_222), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_167), .A2(n_145), .B1(n_161), .B2(n_150), .Y(n_245) );
BUFx4f_ASAP7_75t_L g246 ( .A(n_196), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_171), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_182), .B(n_145), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_166), .B(n_154), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_166), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_192), .B(n_150), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_214), .A2(n_217), .B1(n_218), .B2(n_201), .Y(n_252) );
INVx8_ASAP7_75t_L g253 ( .A(n_214), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_168), .B(n_135), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_222), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_176), .A2(n_135), .B(n_153), .C(n_138), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_165), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_168), .B(n_153), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_214), .Y(n_260) );
AND2x6_ASAP7_75t_L g261 ( .A(n_214), .B(n_153), .Y(n_261) );
INVxp67_ASAP7_75t_SL g262 ( .A(n_217), .Y(n_262) );
INVx4_ASAP7_75t_L g263 ( .A(n_217), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_165), .Y(n_264) );
INVx4_ASAP7_75t_L g265 ( .A(n_217), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_218), .Y(n_266) );
AND3x2_ASAP7_75t_SL g267 ( .A(n_221), .B(n_162), .C(n_159), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_202), .B(n_147), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_180), .Y(n_269) );
INVx8_ASAP7_75t_L g270 ( .A(n_218), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_168), .B(n_193), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_199), .Y(n_272) );
INVx4_ASAP7_75t_L g273 ( .A(n_218), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_169), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_180), .A2(n_142), .B1(n_153), .B2(n_155), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_202), .B(n_142), .Y(n_276) );
AND2x4_ASAP7_75t_SL g277 ( .A(n_221), .B(n_162), .Y(n_277) );
BUFx8_ASAP7_75t_L g278 ( .A(n_168), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_169), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_193), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_174), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_178), .B(n_159), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_210), .B(n_215), .Y(n_283) );
BUFx4f_ASAP7_75t_SL g284 ( .A(n_193), .Y(n_284) );
NAND2xp33_ASAP7_75t_SL g285 ( .A(n_177), .B(n_162), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_268), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_253), .Y(n_287) );
NOR2x1_ASAP7_75t_SL g288 ( .A(n_263), .B(n_182), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_253), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_228), .A2(n_176), .B(n_213), .C(n_211), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_278), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_278), .Y(n_292) );
INVx4_ASAP7_75t_L g293 ( .A(n_253), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_238), .B(n_188), .Y(n_294) );
CKINVDCx11_ASAP7_75t_R g295 ( .A(n_242), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_238), .Y(n_296) );
NAND2xp33_ASAP7_75t_L g297 ( .A(n_261), .B(n_171), .Y(n_297) );
CKINVDCx11_ASAP7_75t_R g298 ( .A(n_242), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_254), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_254), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_259), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_270), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_270), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_262), .B(n_193), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_258), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_223), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_264), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_274), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_262), .B(n_176), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
INVx2_ASAP7_75t_SL g312 ( .A(n_270), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_277), .A2(n_176), .B1(n_213), .B2(n_211), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_281), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_227), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_284), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_284), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_263), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_240), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_261), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g322 ( .A1(n_228), .A2(n_184), .B1(n_187), .B2(n_220), .C1(n_197), .C2(n_200), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_265), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_252), .A2(n_220), .B1(n_213), .B2(n_211), .Y(n_324) );
NOR2xp67_ASAP7_75t_SL g325 ( .A(n_265), .B(n_182), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_248), .A2(n_212), .B(n_182), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_276), .B(n_211), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_261), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_260), .A2(n_212), .B(n_213), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_261), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_229), .A2(n_220), .B1(n_189), .B2(n_206), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_276), .B(n_198), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_233), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_286), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_322), .A2(n_282), .B1(n_237), .B2(n_232), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_331), .B(n_285), .C(n_275), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_296), .B(n_250), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_332), .Y(n_338) );
OR2x6_ASAP7_75t_L g339 ( .A(n_293), .B(n_273), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_294), .B(n_269), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_294), .B(n_246), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_332), .B(n_246), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_316), .A2(n_243), .B1(n_255), .B2(n_236), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_293), .B(n_273), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_320), .Y(n_345) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_307), .Y(n_346) );
AOI211xp5_ASAP7_75t_L g347 ( .A1(n_333), .A2(n_249), .B(n_283), .C(n_235), .Y(n_347) );
AOI222xp33_ASAP7_75t_L g348 ( .A1(n_315), .A2(n_220), .B1(n_271), .B2(n_251), .C1(n_260), .C2(n_267), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_302), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_293), .B(n_244), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_304), .A2(n_266), .B1(n_256), .B2(n_234), .Y(n_351) );
OAI21x1_ASAP7_75t_L g352 ( .A1(n_308), .A2(n_206), .B(n_234), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_304), .B(n_245), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_306), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_324), .A2(n_239), .B1(n_256), .B2(n_244), .Y(n_355) );
NAND2x1_ASAP7_75t_L g356 ( .A(n_302), .B(n_266), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_309), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_308), .A2(n_251), .B1(n_280), .B2(n_189), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_315), .A2(n_244), .B1(n_206), .B2(n_267), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
OAI22xp33_ASAP7_75t_SL g361 ( .A1(n_291), .A2(n_226), .B1(n_244), .B2(n_159), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_307), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_314), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_348), .A2(n_313), .B1(n_299), .B2(n_305), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_335), .A2(n_311), .B1(n_327), .B2(n_300), .Y(n_365) );
BUFx8_ASAP7_75t_L g366 ( .A(n_350), .Y(n_366) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_352), .A2(n_297), .B(n_290), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_345), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_338), .B(n_301), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_335), .B(n_310), .Y(n_370) );
BUFx12f_ASAP7_75t_L g371 ( .A(n_339), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_342), .B(n_311), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_328), .B1(n_310), .B2(n_155), .Y(n_373) );
INVx2_ASAP7_75t_SL g374 ( .A(n_344), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_354), .B(n_287), .Y(n_375) );
CKINVDCx9p33_ASAP7_75t_R g376 ( .A(n_341), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_346), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_357), .B(n_287), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_363), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_352), .A2(n_297), .B(n_320), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_351), .B(n_302), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_345), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_359), .A2(n_318), .B1(n_317), .B2(n_323), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_340), .B(n_302), .Y(n_385) );
AOI222xp33_ASAP7_75t_L g386 ( .A1(n_334), .A2(n_298), .B1(n_295), .B2(n_291), .C1(n_292), .C2(n_317), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_336), .B(n_125), .C(n_131), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_345), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_362), .A2(n_318), .B1(n_319), .B2(n_323), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_343), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_379), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_366), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_379), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_385), .Y(n_394) );
OA21x2_ASAP7_75t_L g395 ( .A1(n_367), .A2(n_152), .B(n_155), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_364), .A2(n_347), .B1(n_292), .B2(n_337), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_365), .A2(n_361), .B1(n_355), .B2(n_351), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_369), .B(n_343), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_372), .B(n_349), .Y(n_399) );
AOI33xp33_ASAP7_75t_L g400 ( .A1(n_375), .A2(n_128), .A3(n_131), .B1(n_358), .B2(n_226), .B3(n_207), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_369), .B(n_360), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_373), .A2(n_358), .B1(n_339), .B2(n_328), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_365), .A2(n_339), .B1(n_289), .B2(n_312), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_366), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_368), .Y(n_405) );
INVxp67_ASAP7_75t_L g406 ( .A(n_386), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_390), .B(n_360), .Y(n_407) );
OAI33xp33_ASAP7_75t_L g408 ( .A1(n_390), .A2(n_131), .A3(n_128), .B1(n_174), .B2(n_175), .B3(n_195), .Y(n_408) );
OAI222xp33_ASAP7_75t_L g409 ( .A1(n_374), .A2(n_344), .B1(n_350), .B2(n_360), .C1(n_321), .C2(n_330), .Y(n_409) );
OAI211xp5_ASAP7_75t_L g410 ( .A1(n_386), .A2(n_128), .B(n_356), .C(n_257), .Y(n_410) );
AOI322xp5_ASAP7_75t_L g411 ( .A1(n_377), .A2(n_195), .A3(n_216), .B1(n_207), .B2(n_198), .C1(n_175), .C2(n_143), .Y(n_411) );
AO22x1_ASAP7_75t_L g412 ( .A1(n_366), .A2(n_350), .B1(n_330), .B2(n_321), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_375), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
AO21x2_ASAP7_75t_L g416 ( .A1(n_367), .A2(n_170), .B(n_186), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_375), .B(n_216), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_373), .A2(n_329), .B(n_272), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_371), .A2(n_289), .B1(n_303), .B2(n_312), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_372), .B(n_303), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_370), .A2(n_319), .B1(n_323), .B2(n_208), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_370), .A2(n_371), .B1(n_381), .B2(n_385), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_381), .Y(n_423) );
AND2x4_ASAP7_75t_SL g424 ( .A(n_374), .B(n_319), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_368), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_391), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_416), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_415), .B(n_368), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_415), .B(n_382), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_392), .B(n_371), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_423), .B(n_374), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_423), .B(n_382), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_416), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_391), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_406), .A2(n_378), .B1(n_383), .B2(n_389), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_397), .A2(n_378), .B1(n_387), .B2(n_376), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_393), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_393), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_407), .B(n_388), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_396), .B(n_378), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_407), .B(n_388), .Y(n_441) );
AOI222xp33_ASAP7_75t_SL g442 ( .A1(n_414), .A2(n_127), .B1(n_186), .B2(n_170), .C1(n_204), .C2(n_191), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_416), .Y(n_443) );
OAI21x1_ASAP7_75t_L g444 ( .A1(n_395), .A2(n_380), .B(n_384), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_394), .B(n_388), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_410), .A2(n_387), .B(n_380), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_417), .B(n_384), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_405), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_425), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_404), .B(n_208), .Y(n_450) );
OAI33xp33_ASAP7_75t_L g451 ( .A1(n_398), .A2(n_170), .A3(n_186), .B1(n_205), .B2(n_204), .B3(n_181), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_425), .B(n_384), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_401), .B(n_382), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_417), .B(n_208), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_401), .B(n_125), .Y(n_455) );
AOI221xp5_ASAP7_75t_SL g456 ( .A1(n_402), .A2(n_125), .B1(n_191), .B2(n_209), .C(n_205), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_422), .B(n_405), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_395), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_399), .B(n_172), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_392), .A2(n_413), .B1(n_404), .B2(n_403), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_395), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_399), .B(n_181), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_400), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_392), .A2(n_127), .B1(n_241), .B2(n_199), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_413), .B(n_23), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_420), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_413), .B(n_209), .Y(n_467) );
AOI33xp33_ASAP7_75t_L g468 ( .A1(n_419), .A2(n_190), .A3(n_172), .B1(n_225), .B2(n_224), .B3(n_231), .Y(n_468) );
OAI22xp5_ASAP7_75t_SL g469 ( .A1(n_420), .A2(n_25), .B1(n_27), .B2(n_30), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_418), .Y(n_470) );
NOR2x1_ASAP7_75t_SL g471 ( .A(n_412), .B(n_320), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_421), .B(n_190), .Y(n_472) );
INVx5_ASAP7_75t_L g473 ( .A(n_412), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_424), .A2(n_127), .B1(n_288), .B2(n_203), .Y(n_474) );
AND4x1_ASAP7_75t_L g475 ( .A(n_465), .B(n_408), .C(n_325), .D(n_411), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_439), .B(n_424), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_439), .B(n_31), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_441), .B(n_33), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_440), .A2(n_127), .B1(n_203), .B2(n_320), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_441), .B(n_37), .Y(n_480) );
AND2x4_ASAP7_75t_SL g481 ( .A(n_466), .B(n_409), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_473), .B(n_320), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_466), .B(n_39), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_453), .B(n_42), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_453), .B(n_44), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_426), .Y(n_486) );
OR2x4_ASAP7_75t_L g487 ( .A(n_450), .B(n_46), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_463), .A2(n_203), .B1(n_171), .B2(n_194), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_428), .B(n_57), .Y(n_489) );
AOI332xp33_ASAP7_75t_L g490 ( .A1(n_426), .A2(n_65), .A3(n_67), .B1(n_68), .B2(n_69), .B3(n_70), .C1(n_71), .C2(n_72), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_434), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_448), .Y(n_492) );
NAND4xp25_ASAP7_75t_SL g493 ( .A(n_468), .B(n_73), .C(n_230), .D(n_288), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_434), .B(n_171), .Y(n_495) );
NAND3xp33_ASAP7_75t_SL g496 ( .A(n_430), .B(n_212), .C(n_326), .Y(n_496) );
OAI211xp5_ASAP7_75t_SL g497 ( .A1(n_435), .A2(n_325), .B(n_212), .C(n_194), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_451), .A2(n_171), .B(n_194), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_437), .Y(n_500) );
OAI31xp33_ASAP7_75t_L g501 ( .A1(n_460), .A2(n_194), .A3(n_240), .B(n_247), .Y(n_501) );
OAI31xp33_ASAP7_75t_SL g502 ( .A1(n_436), .A2(n_194), .A3(n_247), .B(n_240), .Y(n_502) );
NAND4xp25_ASAP7_75t_SL g503 ( .A(n_435), .B(n_194), .C(n_247), .D(n_456), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_428), .B(n_429), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_429), .B(n_457), .Y(n_505) );
NAND4xp25_ASAP7_75t_SL g506 ( .A(n_456), .B(n_442), .C(n_474), .D(n_463), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_448), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_438), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_473), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_438), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_457), .B(n_432), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_448), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_432), .B(n_449), .Y(n_513) );
NAND2x1_ASAP7_75t_L g514 ( .A(n_449), .B(n_458), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_473), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_469), .A2(n_466), .B1(n_470), .B2(n_431), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_432), .B(n_452), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_452), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_447), .B(n_445), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_431), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_462), .B(n_455), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_458), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_432), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_462), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_455), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_459), .Y(n_526) );
NAND3xp33_ASAP7_75t_SL g527 ( .A(n_467), .B(n_446), .C(n_454), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_470), .B(n_467), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_461), .B(n_427), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_461), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_427), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_482), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_494), .B(n_427), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_486), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_526), .B(n_473), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_486), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_505), .B(n_433), .Y(n_537) );
OAI31xp33_ASAP7_75t_L g538 ( .A1(n_493), .A2(n_469), .A3(n_472), .B(n_433), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_507), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_507), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_517), .B(n_433), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_524), .B(n_473), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g543 ( .A(n_506), .B(n_472), .C(n_443), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_509), .B(n_473), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_491), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_491), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_505), .B(n_443), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_517), .B(n_443), .Y(n_548) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_527), .B(n_444), .C(n_471), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_529), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_504), .B(n_444), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_504), .B(n_471), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_511), .B(n_464), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_509), .B(n_515), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_511), .B(n_513), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_514), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_519), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_514), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_518), .B(n_520), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_476), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_498), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_513), .B(n_518), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_498), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_508), .B(n_510), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_521), .B(n_481), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_515), .B(n_523), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_500), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_529), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_528), .B(n_492), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_500), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_522), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_523), .B(n_522), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_510), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_481), .B(n_475), .Y(n_574) );
XOR2x2_ASAP7_75t_L g575 ( .A(n_476), .B(n_516), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_525), .B(n_530), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_530), .B(n_512), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_512), .B(n_531), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_531), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_489), .B(n_477), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_489), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_562), .B(n_487), .Y(n_582) );
NAND2xp33_ASAP7_75t_SL g583 ( .A(n_557), .B(n_515), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_557), .B(n_487), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_562), .B(n_487), .Y(n_585) );
XOR2x2_ASAP7_75t_L g586 ( .A(n_575), .B(n_485), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_571), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_569), .B(n_485), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_569), .B(n_484), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_534), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_540), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_559), .B(n_484), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_534), .Y(n_593) );
XOR2xp5_ASAP7_75t_L g594 ( .A(n_575), .B(n_477), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_555), .B(n_478), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_536), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_555), .B(n_478), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_536), .Y(n_598) );
XOR2xp5_ASAP7_75t_L g599 ( .A(n_581), .B(n_480), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_551), .B(n_480), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_551), .B(n_495), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_571), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_541), .B(n_495), .Y(n_603) );
AOI32xp33_ASAP7_75t_L g604 ( .A1(n_574), .A2(n_497), .A3(n_490), .B1(n_479), .B2(n_502), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_545), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_545), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_546), .Y(n_607) );
NAND2xp33_ASAP7_75t_SL g608 ( .A(n_554), .B(n_483), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_541), .B(n_501), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_560), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_552), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_565), .B(n_503), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_546), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_537), .B(n_488), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_547), .B(n_496), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_550), .B(n_499), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_561), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_561), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_567), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_538), .A2(n_558), .B(n_556), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g621 ( .A1(n_554), .A2(n_544), .B(n_543), .C(n_549), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_535), .B(n_576), .C(n_579), .Y(n_622) );
NAND2x1_ASAP7_75t_L g623 ( .A(n_554), .B(n_544), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_548), .B(n_568), .Y(n_624) );
NAND2x1_ASAP7_75t_L g625 ( .A(n_544), .B(n_566), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_553), .A2(n_542), .B1(n_580), .B2(n_548), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_567), .A2(n_573), .B1(n_570), .B2(n_563), .C(n_564), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_550), .B(n_568), .Y(n_628) );
XNOR2x1_ASAP7_75t_L g629 ( .A(n_553), .B(n_566), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_570), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_573), .Y(n_631) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_566), .B(n_533), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_572), .B(n_577), .Y(n_633) );
AOI21xp33_ASAP7_75t_L g634 ( .A1(n_532), .A2(n_533), .B(n_579), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_532), .B(n_539), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_532), .B(n_539), .Y(n_636) );
XNOR2x1_ASAP7_75t_L g637 ( .A(n_572), .B(n_577), .Y(n_637) );
XNOR2x1_ASAP7_75t_L g638 ( .A(n_578), .B(n_532), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_591), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_594), .A2(n_621), .B1(n_638), .B2(n_623), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_628), .B(n_637), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g642 ( .A1(n_612), .A2(n_615), .B(n_584), .Y(n_642) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_620), .A2(n_612), .B(n_584), .C(n_610), .Y(n_643) );
NAND3xp33_ASAP7_75t_SL g644 ( .A(n_583), .B(n_625), .C(n_604), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_634), .A2(n_627), .B1(n_622), .B2(n_583), .C(n_626), .Y(n_645) );
XOR2xp5_ASAP7_75t_L g646 ( .A(n_586), .B(n_599), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_607), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_629), .B(n_633), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_586), .A2(n_609), .B1(n_608), .B2(n_632), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_634), .A2(n_608), .B(n_582), .C(n_585), .Y(n_650) );
OA22x2_ASAP7_75t_L g651 ( .A1(n_611), .A2(n_597), .B1(n_595), .B2(n_588), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_644), .A2(n_643), .B(n_640), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g653 ( .A(n_649), .B(n_609), .C(n_614), .D(n_627), .Y(n_653) );
OAI22x1_ASAP7_75t_L g654 ( .A1(n_646), .A2(n_636), .B1(n_635), .B2(n_589), .Y(n_654) );
NOR2x1p5_ASAP7_75t_L g655 ( .A(n_641), .B(n_628), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g656 ( .A1(n_649), .A2(n_600), .B(n_592), .C(n_616), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_645), .A2(n_601), .B(n_603), .C(n_624), .Y(n_657) );
NAND3xp33_ASAP7_75t_SL g658 ( .A(n_650), .B(n_601), .C(n_603), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_L g659 ( .A1(n_652), .A2(n_642), .B(n_639), .C(n_648), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_654), .Y(n_660) );
AOI211xp5_ASAP7_75t_L g661 ( .A1(n_658), .A2(n_647), .B(n_651), .C(n_532), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_653), .A2(n_605), .B1(n_630), .B2(n_590), .Y(n_662) );
OAI22xp5_ASAP7_75t_SL g663 ( .A1(n_660), .A2(n_657), .B1(n_656), .B2(n_655), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_661), .A2(n_606), .B1(n_619), .B2(n_593), .Y(n_664) );
XOR2xp5_ASAP7_75t_L g665 ( .A(n_662), .B(n_618), .Y(n_665) );
OAI22xp5_ASAP7_75t_SL g666 ( .A1(n_663), .A2(n_659), .B1(n_631), .B2(n_596), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_665), .A2(n_664), .B1(n_598), .B2(n_613), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_667), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_668), .Y(n_669) );
OR4x1_ASAP7_75t_L g670 ( .A(n_669), .B(n_666), .C(n_617), .D(n_602), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_578), .B1(n_587), .B2(n_602), .C(n_666), .Y(n_671) );
endmodule