module fake_jpeg_12842_n_417 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_417);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_417;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_71),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_14),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_70),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_60),
.Y(n_99)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_65),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g78 ( 
.A(n_64),
.Y(n_78)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_34),
.B(n_37),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_69),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_15),
.B(n_13),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_73),
.Y(n_111)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_15),
.B1(n_37),
.B2(n_19),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_75),
.A2(n_84),
.B1(n_106),
.B2(n_18),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_81),
.A2(n_94),
.B(n_101),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_16),
.B1(n_33),
.B2(n_27),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_39),
.A2(n_16),
.B1(n_33),
.B2(n_27),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_110),
.B1(n_113),
.B2(n_17),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_16),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_88),
.B(n_103),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_25),
.C(n_36),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_25),
.B1(n_36),
.B2(n_18),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_50),
.B(n_37),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_49),
.A2(n_19),
.B1(n_33),
.B2(n_27),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_19),
.B1(n_32),
.B2(n_31),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_109),
.A2(n_67),
.B(n_66),
.C(n_72),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_41),
.A2(n_36),
.B1(n_32),
.B2(n_31),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_42),
.A2(n_32),
.B1(n_31),
.B2(n_25),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_64),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_56),
.Y(n_144)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_118),
.A2(n_143),
.B1(n_48),
.B2(n_102),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_71),
.B1(n_64),
.B2(n_59),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_120),
.Y(n_189)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_24),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_140),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_123),
.Y(n_195)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_71),
.B1(n_59),
.B2(n_53),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_144),
.B1(n_152),
.B2(n_155),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_12),
.C(n_13),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_127),
.B(n_136),
.Y(n_181)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_132),
.A2(n_99),
.B1(n_76),
.B2(n_95),
.Y(n_191)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_65),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_142),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_17),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_73),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_111),
.B(n_38),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_108),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_147),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_77),
.B(n_69),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_149),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_154),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_100),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_107),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_153),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_77),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_107),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_99),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_130),
.C(n_137),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_166),
.C(n_186),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_101),
.Y(n_166)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_109),
.B(n_92),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_188),
.B(n_22),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_113),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_185),
.Y(n_200)
);

NOR2xp67_ASAP7_75t_R g180 ( 
.A(n_143),
.B(n_52),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_SL g233 ( 
.A(n_180),
.B(n_2),
.C(n_3),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_114),
.B1(n_105),
.B2(n_76),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_SL g229 ( 
.A1(n_184),
.A2(n_187),
.B(n_0),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_105),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_89),
.C(n_68),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_17),
.B(n_18),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_117),
.B1(n_146),
.B2(n_149),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_116),
.B(n_124),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_24),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_157),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_190),
.C(n_183),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_199),
.A2(n_202),
.B1(n_224),
.B2(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_201),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_149),
.B1(n_146),
.B2(n_128),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_158),
.A2(n_134),
.B(n_133),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_203),
.A2(n_214),
.B(n_215),
.Y(n_236)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_205),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_158),
.A2(n_132),
.B1(n_152),
.B2(n_131),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_206),
.A2(n_207),
.B1(n_213),
.B2(n_227),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_178),
.A2(n_120),
.B1(n_90),
.B2(n_125),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_159),
.B(n_135),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_209),
.B(n_210),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_172),
.B(n_155),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_167),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_220),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_177),
.A2(n_90),
.B1(n_83),
.B2(n_89),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_182),
.A2(n_121),
.B(n_52),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_171),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_216),
.B(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_221),
.Y(n_270)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_163),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_166),
.B(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_180),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_190),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_164),
.A2(n_175),
.B1(n_187),
.B2(n_173),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_182),
.A2(n_102),
.B1(n_83),
.B2(n_147),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_24),
.B1(n_22),
.B2(n_129),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_162),
.A2(n_22),
.B1(n_129),
.B2(n_147),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_173),
.B(n_0),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_168),
.B1(n_169),
.B2(n_176),
.Y(n_249)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_174),
.B(n_1),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_192),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_233),
.A2(n_179),
.B(n_160),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_186),
.A2(n_13),
.B1(n_12),
.B2(n_4),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_193),
.B(n_194),
.Y(n_264)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_223),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_250),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_188),
.B(n_195),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_242),
.A2(n_265),
.B(n_235),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_232),
.Y(n_243)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_246),
.C(n_256),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_190),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_247),
.A2(n_257),
.B(n_228),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_199),
.B1(n_234),
.B2(n_198),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_215),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_168),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g300 ( 
.A(n_252),
.B(n_256),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_262),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_197),
.B(n_168),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_223),
.A2(n_169),
.B1(n_176),
.B2(n_160),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_206),
.B1(n_207),
.B2(n_227),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_220),
.A2(n_200),
.B(n_214),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_201),
.B(n_181),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_202),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_269),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_SL g271 ( 
.A(n_254),
.B(n_213),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_271),
.A2(n_273),
.B(n_274),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_250),
.A2(n_200),
.B(n_204),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_267),
.A2(n_198),
.B1(n_217),
.B2(n_203),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_276),
.A2(n_280),
.B1(n_298),
.B2(n_299),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_278),
.A2(n_293),
.B1(n_297),
.B2(n_237),
.Y(n_308)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_240),
.Y(n_279)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_281),
.Y(n_312)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_282),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_236),
.A2(n_231),
.B(n_218),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_283),
.B(n_291),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_267),
.A2(n_230),
.B1(n_222),
.B2(n_219),
.Y(n_284)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_262),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_237),
.A2(n_205),
.B1(n_208),
.B2(n_193),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_257),
.B(n_247),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_246),
.B(n_194),
.C(n_189),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_292),
.C(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_244),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_290),
.Y(n_302)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_179),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_251),
.A2(n_258),
.B1(n_266),
.B2(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_294),
.B(n_296),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_261),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_249),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_SL g299 ( 
.A1(n_236),
.A2(n_2),
.B(n_5),
.C(n_6),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_270),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_273),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_277),
.B(n_270),
.C(n_247),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_315),
.C(n_318),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_272),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_307),
.B(n_309),
.Y(n_346)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_308),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_272),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_320),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_287),
.A2(n_265),
.B1(n_242),
.B2(n_248),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_316),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_255),
.C(n_260),
.Y(n_315)
);

INVx3_ASAP7_75t_SL g316 ( 
.A(n_293),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_260),
.C(n_259),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_285),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_321),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_295),
.C(n_274),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_304),
.C(n_315),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_259),
.B1(n_239),
.B2(n_263),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_323),
.A2(n_325),
.B1(n_279),
.B2(n_281),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_286),
.B(n_275),
.Y(n_324)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_324),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_283),
.B1(n_278),
.B2(n_291),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_305),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_331),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_316),
.A2(n_297),
.B1(n_288),
.B2(n_294),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_318),
.B(n_299),
.CI(n_290),
.CON(n_334),
.SN(n_334)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_306),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_303),
.A2(n_282),
.B1(n_299),
.B2(n_263),
.Y(n_335)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_238),
.Y(n_336)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_322),
.C(n_313),
.Y(n_354)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_319),
.Y(n_338)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_303),
.A2(n_299),
.B1(n_238),
.B2(n_8),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_339),
.A2(n_317),
.B1(n_312),
.B2(n_326),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_299),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_342),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_325),
.A2(n_2),
.B1(n_6),
.B2(n_8),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_345),
.Y(n_350)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_311),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_310),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_347),
.B(n_348),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_323),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_327),
.A2(n_306),
.B(n_314),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_349),
.A2(n_360),
.B(n_355),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_351),
.A2(n_344),
.B(n_346),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_357),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_332),
.C(n_337),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_356),
.A2(n_329),
.B1(n_343),
.B2(n_345),
.Y(n_376)
);

XOR2x1_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_321),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_330),
.B(n_320),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_359),
.B(n_328),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_360),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_308),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_341),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_371),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_367),
.Y(n_384)
);

INVx6_ASAP7_75t_L g369 ( 
.A(n_358),
.Y(n_369)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_369),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_373),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_350),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_372),
.B(n_352),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_362),
.A2(n_329),
.B1(n_340),
.B2(n_331),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_353),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_363),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_334),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_378),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_344),
.B1(n_342),
.B2(n_334),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_365),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_336),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_354),
.C(n_364),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_385),
.Y(n_400)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_373),
.B(n_349),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_387),
.B(n_388),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_369),
.A2(n_353),
.B1(n_361),
.B2(n_350),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_389),
.B(n_379),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_391),
.B(n_368),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_382),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_393),
.B(n_394),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_384),
.B(n_366),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_390),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_381),
.A2(n_374),
.B1(n_370),
.B2(n_378),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_397),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_383),
.A2(n_368),
.B(n_376),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_398),
.B(n_399),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_402),
.B(n_406),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_400),
.B(n_380),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_404),
.B(n_392),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_380),
.Y(n_406)
);

OAI321xp33_ASAP7_75t_L g407 ( 
.A1(n_397),
.A2(n_386),
.A3(n_357),
.B1(n_341),
.B2(n_10),
.C(n_6),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_407),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_409),
.A2(n_401),
.B(n_405),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_403),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_410),
.A2(n_411),
.B(n_401),
.Y(n_413)
);

OAI21xp33_ASAP7_75t_L g414 ( 
.A1(n_412),
.A2(n_413),
.B(n_408),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_414),
.A2(n_11),
.B(n_8),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_415),
.B(n_9),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_9),
.Y(n_417)
);


endmodule