module fake_jpeg_3816_n_39 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_39);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_10),
.B(n_0),
.C(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_28),
.B(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_4),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_20),
.A2(n_22),
.B1(n_14),
.B2(n_23),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_24),
.B1(n_16),
.B2(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_15),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_31),
.C(n_34),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_30),
.B(n_32),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_30),
.Y(n_39)
);


endmodule