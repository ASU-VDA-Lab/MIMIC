module fake_jpeg_9633_n_60 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

BUFx3_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_4),
.B(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_0),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_19),
.A2(n_23),
.B(n_17),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

BUFx24_ASAP7_75t_SL g24 ( 
.A(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_11),
.B(n_13),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_20),
.B(n_22),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_16),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_15),
.B1(n_16),
.B2(n_14),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_34),
.B1(n_13),
.B2(n_14),
.Y(n_41)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_21),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_13),
.C(n_18),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2x1_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_40),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_32),
.B1(n_33),
.B2(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_39),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_40),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_52),
.Y(n_54)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_30),
.Y(n_52)
);

MAJx2_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_48),
.C(n_50),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_44),
.C(n_47),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.C(n_53),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_2),
.C(n_3),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_55),
.C(n_6),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_6),
.Y(n_60)
);


endmodule