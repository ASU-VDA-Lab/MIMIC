module fake_jpeg_13313_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_5),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_12),
.B(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

NAND2x1_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_21),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_64),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_26),
.B1(n_15),
.B2(n_16),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_61),
.A2(n_31),
.B(n_20),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_30),
.B(n_14),
.C(n_16),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_42),
.C(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_22),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_14),
.B(n_15),
.C(n_22),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_0),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_28),
.A2(n_20),
.B1(n_21),
.B2(n_2),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_36),
.B1(n_41),
.B2(n_3),
.Y(n_77)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_11),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_83),
.B1(n_68),
.B2(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_83),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_40),
.C(n_3),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_61),
.B(n_56),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_11),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_62),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_65),
.B1(n_56),
.B2(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_67),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_71),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_45),
.B1(n_60),
.B2(n_54),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_73),
.B1(n_82),
.B2(n_76),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_78),
.B1(n_80),
.B2(n_79),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_107),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_106),
.B1(n_110),
.B2(n_112),
.Y(n_113)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_108),
.B(n_89),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_111),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_81),
.B1(n_69),
.B2(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_94),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_62),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_89),
.C(n_97),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_100),
.B1(n_90),
.B2(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_1),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_90),
.B(n_95),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_117),
.B(n_87),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_93),
.B(n_94),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_93),
.B1(n_89),
.B2(n_86),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_120),
.B1(n_87),
.B2(n_105),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_109),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_116),
.C(n_113),
.Y(n_128)
);

OAI322xp33_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_105),
.A3(n_86),
.B1(n_98),
.B2(n_46),
.C1(n_87),
.C2(n_3),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_115),
.C(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_126),
.A2(n_127),
.B1(n_49),
.B2(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_130),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_131),
.A2(n_125),
.B1(n_127),
.B2(n_49),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_132),
.B(n_134),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_129),
.C(n_134),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_46),
.C(n_40),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_135),
.B(n_49),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_40),
.Y(n_139)
);


endmodule