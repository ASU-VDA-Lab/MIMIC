module fake_ariane_3282_n_730 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_730);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_730;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_500;
wire n_665;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_672;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_166;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_492;
wire n_234;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_517;
wire n_246;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_33),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_35),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_60),
.Y(n_154)
);

BUFx10_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_36),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_16),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_48),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_10),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_37),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_118),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_62),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_45),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_53),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_72),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_52),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_29),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_40),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_81),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_76),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_79),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_46),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_42),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_39),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_88),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_68),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_28),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_90),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_77),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_111),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_93),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_49),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_29),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_91),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_95),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_63),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_41),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_7),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_143),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_67),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_9),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_43),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_8),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_80),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_98),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_47),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_71),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_117),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_105),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_96),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_26),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_65),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_78),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_86),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_61),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_5),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_11),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_110),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_33),
.Y(n_231)
);

CKINVDCx11_ASAP7_75t_R g232 ( 
.A(n_140),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_50),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_129),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_34),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_112),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_64),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_3),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_82),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_1),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_23),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_97),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_5),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_17),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_54),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_38),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_11),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_101),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_25),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_17),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_139),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_66),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_142),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_51),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_114),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_15),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_58),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_84),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_28),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_8),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_100),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_69),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_25),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_141),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_2),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_9),
.Y(n_266)
);

INVxp33_ASAP7_75t_SL g267 ( 
.A(n_192),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_250),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_157),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_194),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

INVx4_ASAP7_75t_R g275 ( 
.A(n_201),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_212),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_172),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_160),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_172),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_185),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_210),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_155),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_155),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_178),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_233),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_201),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_178),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_180),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_180),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_236),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_198),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_150),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_151),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_152),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_156),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_205),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_209),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_159),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_219),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_162),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_165),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_168),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_264),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_170),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_223),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_228),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_229),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_240),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_174),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_176),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_193),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_179),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_181),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_235),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_183),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_243),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_186),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_187),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_190),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_244),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_191),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_249),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_203),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_204),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_256),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_206),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_207),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_208),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_211),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_214),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_216),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_217),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_263),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_231),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_218),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_219),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_153),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_220),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_221),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_222),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_225),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g351 ( 
.A(n_247),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_242),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_251),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_253),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_254),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_334),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_153),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_281),
.B(n_255),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_351),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_272),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_293),
.B(n_257),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_293),
.B(n_346),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_267),
.A2(n_323),
.B1(n_343),
.B2(n_271),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_202),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_334),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_299),
.B(n_262),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_306),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_333),
.Y(n_369)
);

BUFx12f_ASAP7_75t_L g370 ( 
.A(n_270),
.Y(n_370)
);

OA21x2_ASAP7_75t_L g371 ( 
.A1(n_320),
.A2(n_213),
.B(n_202),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

NAND2xp33_ASAP7_75t_L g373 ( 
.A(n_301),
.B(n_193),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_282),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_302),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_317),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_273),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_276),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_355),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_286),
.A2(n_213),
.B1(n_237),
.B2(n_224),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_298),
.B(n_224),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_307),
.B(n_189),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_269),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_308),
.A2(n_237),
.B(n_188),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_283),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_310),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_289),
.B(n_196),
.Y(n_392)
);

NOR2x1_ASAP7_75t_L g393 ( 
.A(n_290),
.B(n_252),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_284),
.Y(n_394)
);

OA21x2_ASAP7_75t_L g395 ( 
.A1(n_312),
.A2(n_173),
.B(n_199),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_319),
.B(n_239),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_280),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_322),
.B(n_154),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_326),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_291),
.B(n_294),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_303),
.B(n_158),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_328),
.Y(n_406)
);

OAI21x1_ASAP7_75t_L g407 ( 
.A1(n_330),
.A2(n_193),
.B(n_164),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_354),
.B(n_161),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

NOR2x1_ASAP7_75t_L g410 ( 
.A(n_295),
.B(n_296),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_335),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_268),
.A2(n_166),
.B1(n_167),
.B2(n_163),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_336),
.A2(n_171),
.B(n_169),
.Y(n_413)
);

AND2x6_ASAP7_75t_L g414 ( 
.A(n_337),
.B(n_164),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_339),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_340),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_314),
.A2(n_304),
.B1(n_313),
.B2(n_287),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_316),
.B(n_164),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_341),
.B(n_175),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_279),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_344),
.B(n_177),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_347),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_348),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_349),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_350),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_369),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

AO22x2_ASAP7_75t_L g430 ( 
.A1(n_363),
.A2(n_390),
.B1(n_412),
.B2(n_357),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_372),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_386),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_374),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_420),
.B(n_325),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_407),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_420),
.B(n_329),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_368),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_368),
.Y(n_440)
);

NOR2x1p5_ASAP7_75t_L g441 ( 
.A(n_370),
.B(n_331),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_368),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_352),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_375),
.Y(n_445)
);

AND3x2_ASAP7_75t_L g446 ( 
.A(n_377),
.B(n_315),
.C(n_278),
.Y(n_446)
);

CKINVDCx6p67_ASAP7_75t_R g447 ( 
.A(n_367),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_342),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_376),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_405),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_380),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_399),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_391),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_381),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_414),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_411),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_416),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_417),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_417),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_424),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_425),
.Y(n_466)
);

AND3x2_ASAP7_75t_L g467 ( 
.A(n_390),
.B(n_277),
.C(n_274),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_404),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_389),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_394),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_415),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_415),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_415),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_388),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_395),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_401),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_360),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_378),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_396),
.B(n_300),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_409),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_388),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

AND3x2_ASAP7_75t_L g484 ( 
.A(n_356),
.B(n_365),
.C(n_403),
.Y(n_484)
);

AOI21x1_ASAP7_75t_L g485 ( 
.A1(n_361),
.A2(n_366),
.B(n_358),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_361),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_427),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_449),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_486),
.B(n_362),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_444),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_430),
.B(n_286),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_288),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_452),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_480),
.B(n_359),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_452),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_456),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_387),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_441),
.B(n_382),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_431),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_457),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_457),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_362),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_436),
.A2(n_373),
.B(n_413),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_451),
.B(n_292),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_485),
.B(n_364),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_455),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_447),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_460),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_461),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_435),
.B(n_419),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_462),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_435),
.B(n_437),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_364),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_463),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_455),
.Y(n_516)
);

AOI21x1_ASAP7_75t_L g517 ( 
.A1(n_475),
.A2(n_358),
.B(n_400),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_448),
.B(n_288),
.Y(n_518)
);

NAND2x1p5_ASAP7_75t_L g519 ( 
.A(n_459),
.B(n_418),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_466),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_467),
.B(n_422),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_455),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_450),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_446),
.B(n_403),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_443),
.B(n_383),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_464),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_428),
.B(n_297),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_464),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_433),
.B(n_311),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_465),
.B(n_383),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_469),
.Y(n_531)
);

CKINVDCx14_ASAP7_75t_R g532 ( 
.A(n_455),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_433),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_487),
.B(n_392),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_494),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_489),
.B(n_502),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_504),
.B(n_458),
.Y(n_539)
);

A2O1A1Ixp33_ASAP7_75t_L g540 ( 
.A1(n_511),
.A2(n_479),
.B(n_483),
.C(n_477),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_489),
.A2(n_436),
.B(n_434),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_490),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_513),
.B(n_458),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_503),
.A2(n_436),
.B(n_434),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_497),
.B(n_474),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_518),
.B(n_474),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_507),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_476),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_533),
.B(n_478),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_506),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_527),
.A2(n_482),
.B1(n_393),
.B2(n_473),
.Y(n_552)
);

NOR3xp33_ASAP7_75t_L g553 ( 
.A(n_529),
.B(n_410),
.C(n_421),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_526),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_530),
.B(n_481),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_519),
.B(n_459),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_528),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_530),
.B(n_470),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_499),
.Y(n_559)
);

A2O1A1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_505),
.A2(n_514),
.B(n_503),
.C(n_536),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_L g561 ( 
.A(n_506),
.B(n_516),
.Y(n_561)
);

A2O1A1Ixp33_ASAP7_75t_L g562 ( 
.A1(n_488),
.A2(n_423),
.B(n_421),
.C(n_373),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_531),
.B(n_438),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_516),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_493),
.B(n_423),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_524),
.B(n_516),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_495),
.B(n_432),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_496),
.B(n_432),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_521),
.B(n_453),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_500),
.B(n_432),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_501),
.B(n_454),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_537),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_538),
.B(n_491),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_550),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_542),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_543),
.B(n_498),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_543),
.B(n_498),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_547),
.B(n_473),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_546),
.B(n_532),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_539),
.A2(n_492),
.B1(n_468),
.B2(n_472),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_542),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_542),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_554),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_566),
.B(n_522),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_557),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_545),
.B(n_517),
.Y(n_586)
);

AO22x1_ASAP7_75t_L g587 ( 
.A1(n_569),
.A2(n_398),
.B1(n_384),
.B2(n_397),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_564),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_540),
.B(n_471),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_551),
.Y(n_590)
);

INVx5_ASAP7_75t_L g591 ( 
.A(n_559),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_R g592 ( 
.A(n_561),
.B(n_508),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_SL g593 ( 
.A(n_565),
.B(n_549),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_563),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_553),
.A2(n_471),
.B1(n_397),
.B2(n_366),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_548),
.B(n_509),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_567),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_571),
.Y(n_598)
);

AOI21x1_ASAP7_75t_L g599 ( 
.A1(n_587),
.A2(n_544),
.B(n_541),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_597),
.A2(n_568),
.B(n_567),
.Y(n_600)
);

AO31x2_ASAP7_75t_L g601 ( 
.A1(n_586),
.A2(n_560),
.A3(n_562),
.B(n_568),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_593),
.A2(n_556),
.B(n_570),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_575),
.Y(n_603)
);

NOR4xp25_ASAP7_75t_L g604 ( 
.A(n_573),
.B(n_558),
.C(n_555),
.D(n_510),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_575),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_579),
.B(n_552),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_572),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_581),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_576),
.B(n_439),
.Y(n_609)
);

AO21x1_ASAP7_75t_L g610 ( 
.A1(n_589),
.A2(n_515),
.B(n_512),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_583),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_594),
.B(n_598),
.Y(n_613)
);

AO31x2_ASAP7_75t_L g614 ( 
.A1(n_596),
.A2(n_534),
.A3(n_535),
.B(n_520),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_581),
.Y(n_615)
);

OAI21x1_ASAP7_75t_SL g616 ( 
.A1(n_585),
.A2(n_442),
.B(n_440),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_577),
.B(n_0),
.Y(n_617)
);

OA21x2_ASAP7_75t_L g618 ( 
.A1(n_595),
.A2(n_184),
.B(n_182),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_581),
.Y(n_619)
);

OAI21x1_ASAP7_75t_SL g620 ( 
.A1(n_582),
.A2(n_4),
.B(n_6),
.Y(n_620)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_580),
.A2(n_197),
.B(n_195),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_617),
.B(n_578),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_602),
.A2(n_584),
.B(n_591),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_599),
.A2(n_592),
.B(n_591),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_621),
.B(n_604),
.C(n_606),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_600),
.A2(n_590),
.B(n_588),
.Y(n_626)
);

AO31x2_ASAP7_75t_L g627 ( 
.A1(n_610),
.A2(n_275),
.A3(n_590),
.B(n_429),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_603),
.Y(n_628)
);

NOR4xp25_ASAP7_75t_L g629 ( 
.A(n_607),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_629)
);

AOI221xp5_ASAP7_75t_L g630 ( 
.A1(n_611),
.A2(n_612),
.B1(n_620),
.B2(n_613),
.C(n_609),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_603),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_618),
.B(n_227),
.C(n_226),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_618),
.A2(n_234),
.B(n_230),
.Y(n_633)
);

NAND2x1_ASAP7_75t_L g634 ( 
.A(n_616),
.B(n_44),
.Y(n_634)
);

AO31x2_ASAP7_75t_L g635 ( 
.A1(n_614),
.A2(n_89),
.A3(n_148),
.B(n_147),
.Y(n_635)
);

O2A1O1Ixp33_ASAP7_75t_SL g636 ( 
.A1(n_608),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_601),
.A2(n_615),
.B(n_605),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_615),
.A2(n_246),
.B(n_245),
.Y(n_638)
);

INVx6_ASAP7_75t_L g639 ( 
.A(n_631),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_625),
.A2(n_619),
.B1(n_261),
.B2(n_258),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_632),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_637),
.Y(n_642)
);

CKINVDCx11_ASAP7_75t_R g643 ( 
.A(n_631),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_630),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_629),
.B(n_32),
.Y(n_645)
);

CKINVDCx6p67_ASAP7_75t_R g646 ( 
.A(n_622),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_628),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_633),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_638),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_626),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_624),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_635),
.Y(n_652)
);

INVx6_ASAP7_75t_L g653 ( 
.A(n_623),
.Y(n_653)
);

INVx3_ASAP7_75t_SL g654 ( 
.A(n_636),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_634),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_650),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_653),
.B(n_627),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_650),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_642),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_651),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_652),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_639),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_647),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_639),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_643),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_646),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_645),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_654),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_655),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_649),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_659),
.B(n_640),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_660),
.B(n_644),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_661),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_660),
.B(n_641),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_663),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_658),
.B(n_648),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_665),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_656),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_670),
.B(n_146),
.Y(n_679)
);

OR2x2_ASAP7_75t_L g680 ( 
.A(n_667),
.B(n_85),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_677),
.B(n_665),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_677),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_678),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_675),
.B(n_668),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_674),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_673),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_685),
.B(n_671),
.Y(n_687)
);

INVx3_ASAP7_75t_SL g688 ( 
.A(n_684),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_682),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_688),
.B(n_684),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_687),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_689),
.B(n_683),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_692),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_691),
.B(n_683),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_693),
.B(n_692),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_694),
.B(n_690),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_695),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_696),
.B(n_665),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_696),
.B(n_681),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_697),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_699),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_698),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_701),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_702),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_700),
.B(n_666),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_704),
.Y(n_706)
);

AOI221xp5_ASAP7_75t_L g707 ( 
.A1(n_703),
.A2(n_669),
.B1(n_674),
.B2(n_672),
.C(n_680),
.Y(n_707)
);

O2A1O1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_705),
.A2(n_679),
.B(n_676),
.C(n_672),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_708),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_707),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_706),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_709),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_710),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_711),
.Y(n_714)
);

NOR3xp33_ASAP7_75t_L g715 ( 
.A(n_714),
.B(n_712),
.C(n_713),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_715),
.B(n_664),
.Y(n_716)
);

NAND2x1p5_ASAP7_75t_L g717 ( 
.A(n_716),
.B(n_662),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_SL g718 ( 
.A1(n_717),
.A2(n_657),
.B1(n_664),
.B2(n_686),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_718),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_719),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_720),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_721),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_722),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_723),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_724),
.A2(n_145),
.B1(n_103),
.B2(n_104),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_724),
.A2(n_99),
.B1(n_107),
.B2(n_109),
.Y(n_726)
);

AO21x1_ASAP7_75t_L g727 ( 
.A1(n_725),
.A2(n_726),
.B(n_113),
.Y(n_727)
);

OA21x2_ASAP7_75t_L g728 ( 
.A1(n_727),
.A2(n_119),
.B(n_122),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_728),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_729)
);

AOI211xp5_ASAP7_75t_L g730 ( 
.A1(n_729),
.A2(n_127),
.B(n_128),
.C(n_131),
.Y(n_730)
);


endmodule