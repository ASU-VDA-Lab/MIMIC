module fake_netlist_1_697_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_30;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
HB1xp67_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_0), .B(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_5), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
BUFx3_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_6), .B(n_3), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_14), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
BUFx3_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_13), .A2(n_10), .B(n_8), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_19), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
INVx2_ASAP7_75t_SL g25 ( .A(n_21), .Y(n_25) );
OAI22xp33_ASAP7_75t_L g26 ( .A1(n_18), .A2(n_15), .B1(n_11), .B2(n_13), .Y(n_26) );
BUFx3_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_24), .Y(n_28) );
NOR4xp25_ASAP7_75t_SL g29 ( .A(n_24), .B(n_12), .C(n_22), .D(n_3), .Y(n_29) );
INVx5_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_28), .B(n_23), .Y(n_31) );
OAI221xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_28), .B1(n_25), .B2(n_27), .C(n_26), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_28), .Y(n_33) );
OAI221xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_27), .B1(n_22), .B2(n_23), .C(n_17), .Y(n_34) );
XNOR2x1_ASAP7_75t_L g35 ( .A(n_33), .B(n_17), .Y(n_35) );
A2O1A1Ixp33_ASAP7_75t_SL g36 ( .A1(n_32), .A2(n_29), .B(n_27), .C(n_30), .Y(n_36) );
AOI22xp33_ASAP7_75t_SL g37 ( .A1(n_35), .A2(n_30), .B1(n_29), .B2(n_4), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_36), .B(n_29), .Y(n_38) );
NOR2xp33_ASAP7_75t_L g39 ( .A(n_34), .B(n_1), .Y(n_39) );
OR3x2_ASAP7_75t_L g40 ( .A(n_37), .B(n_2), .C(n_4), .Y(n_40) );
AOI322xp5_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_5), .A3(n_7), .B1(n_30), .B2(n_38), .C1(n_37), .C2(n_39), .Y(n_41) );
endmodule