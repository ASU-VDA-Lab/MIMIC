module real_jpeg_24518_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_285;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_240;
wire n_55;
wire n_185;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_128;
wire n_213;
wire n_179;
wire n_295;
wire n_167;
wire n_133;
wire n_202;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_269;
wire n_96;
wire n_273;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_0),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_0),
.B(n_2),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_2),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_2),
.A2(n_20),
.B1(n_48),
.B2(n_49),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_2),
.A2(n_20),
.B1(n_63),
.B2(n_64),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_20),
.B1(n_30),
.B2(n_31),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_2),
.A2(n_28),
.B(n_186),
.C(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_2),
.B(n_29),
.Y(n_202)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_2),
.A2(n_31),
.B(n_44),
.C(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_2),
.B(n_60),
.C(n_63),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_2),
.B(n_73),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_2),
.B(n_62),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_5),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_7),
.A2(n_21),
.B1(n_22),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_7),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_131),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_131),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_131),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_21),
.B1(n_23),
.B2(n_51),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_11),
.A2(n_51),
.B1(n_63),
.B2(n_64),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_111),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_110),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_95),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_15),
.B(n_95),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_71),
.C(n_80),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_16),
.B(n_71),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_38),
.B1(n_69),
.B2(n_70),
.Y(n_16)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_17),
.A2(n_69),
.B1(n_97),
.B2(n_108),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_17),
.B(n_40),
.C(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_33),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_18),
.B(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_19),
.B(n_29),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_20),
.A2(n_27),
.B(n_31),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_20),
.A2(n_46),
.B(n_48),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_21),
.Y(n_187)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_25),
.B(n_34),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_25),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_29),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_29),
.B(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_31),
.B1(n_44),
.B2(n_46),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx6p67_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_33),
.B(n_129),
.Y(n_181)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_50),
.B(n_52),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_41),
.B(n_103),
.Y(n_135)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_42),
.B(n_53),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_42),
.A2(n_47),
.B(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_42),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_102),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_49),
.B(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_52),
.B(n_179),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_54),
.A2(n_55),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_54),
.B(n_168),
.C(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_54),
.A2(n_55),
.B1(n_170),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_66),
.B(n_67),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_57),
.B(n_68),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_57),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_62),
.B(n_217),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_63),
.B(n_253),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_67),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_66),
.A2(n_78),
.B(n_88),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_71),
.A2(n_72),
.B(n_75),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_73),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_74),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_76),
.B(n_215),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_78),
.B(n_227),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_80),
.B(n_302),
.Y(n_301)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_86),
.B(n_90),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_81),
.A2(n_87),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_81),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_90),
.B1(n_91),
.B2(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_81),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_81),
.A2(n_138),
.B1(n_212),
.B2(n_269),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_82),
.B(n_85),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_82),
.B(n_241),
.Y(n_240)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_86),
.B(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_87),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_89),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_89),
.B(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_109),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_101),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_107),
.B(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_298),
.B(n_303),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_160),
.B(n_297),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_152),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_115),
.B(n_152),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_136),
.C(n_139),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_116),
.B(n_136),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_125),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_126),
.C(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_118),
.B(n_124),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_119),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_120),
.B(n_242),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_122),
.A2(n_143),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_122),
.B(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_135),
.B(n_172),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_139),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.C(n_150),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_140),
.A2(n_141),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_147),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_145),
.B(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_148),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_149),
.A2(n_150),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_149),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_150),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_154),
.B(n_158),
.C(n_159),
.Y(n_300)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_292),
.B(n_296),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_205),
.B(n_278),
.C(n_291),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_193),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_163),
.B(n_193),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_176),
.B2(n_192),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_174),
.B2(n_175),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_166),
.B(n_175),
.C(n_192),
.Y(n_279)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_169),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_184),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_178),
.B(n_183),
.C(n_184),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_181),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.C(n_200),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_195),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_200),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.C(n_203),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_203),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_277),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_221),
.B(n_276),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_208),
.B(n_218),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.C(n_214),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_209),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_211),
.B(n_214),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_212),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_271),
.B(n_275),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_262),
.B(n_270),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_244),
.B(n_261),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_231),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_225),
.B(n_231),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_226),
.A2(n_228),
.B1(n_229),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_238),
.B2(n_243),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_234),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_237),
.C(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_235),
.Y(n_237)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_250),
.B(n_260),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_246),
.B(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_256),
.B(n_259),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_264),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_272),
.B(n_273),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_280),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_290),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_288),
.B2(n_289),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_289),
.C(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);


endmodule