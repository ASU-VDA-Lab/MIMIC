module real_jpeg_26660_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_298, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_298;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_288;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_216;
wire n_244;
wire n_128;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

INVx11_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_1),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_130),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_130),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_1),
.A2(n_29),
.B1(n_35),
.B2(n_130),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_2),
.A2(n_41),
.B1(n_62),
.B2(n_63),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_2),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_2),
.A2(n_29),
.B1(n_35),
.B2(n_41),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_5),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_5),
.A2(n_46),
.B(n_50),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_5),
.B(n_48),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_5),
.A2(n_62),
.B(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_62),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_5),
.B(n_101),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_5),
.A2(n_27),
.B1(n_32),
.B2(n_223),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_5),
.A2(n_49),
.B(n_240),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_6),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_141),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_6),
.A2(n_62),
.B1(n_63),
.B2(n_141),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_141),
.Y(n_223)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_8),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_86),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_29),
.B1(n_35),
.B2(n_86),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_9),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_9),
.A2(n_36),
.B1(n_62),
.B2(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_29),
.B1(n_35),
.B2(n_64),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_11),
.A2(n_29),
.B1(n_35),
.B2(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_11),
.A2(n_35),
.A3(n_62),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_12),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_73),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_73),
.Y(n_113)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_14),
.A2(n_49),
.B(n_79),
.C(n_82),
.Y(n_78)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_14),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_14),
.A2(n_62),
.B1(n_63),
.B2(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_15),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_15),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_15),
.A2(n_29),
.B1(n_35),
.B2(n_54),
.Y(n_155)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_17),
.A2(n_42),
.B1(n_43),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_17),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_17),
.A2(n_49),
.B1(n_50),
.B2(n_104),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_17),
.A2(n_29),
.B1(n_35),
.B2(n_104),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_17),
.A2(n_62),
.B1(n_63),
.B2(n_104),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_105),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_22),
.B(n_105),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.C(n_91),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_23),
.B(n_76),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_56),
.B1(n_57),
.B2(n_75),
.Y(n_23)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_25),
.A2(n_38),
.B(n_56),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_25),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_27),
.A2(n_33),
.B1(n_34),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_27),
.A2(n_33),
.B1(n_95),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_27),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_27),
.A2(n_33),
.B1(n_217),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_27),
.A2(n_33),
.B1(n_211),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_28),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_28),
.A2(n_31),
.B1(n_146),
.B2(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_28),
.A2(n_147),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_29),
.B(n_68),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_29),
.B(n_228),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g212 ( 
.A(n_31),
.Y(n_212)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_33),
.Y(n_147)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_53),
.B2(n_55),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_40),
.A2(n_45),
.B1(n_48),
.B2(n_103),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_42),
.A2(n_52),
.B(n_139),
.C(n_144),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_46),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_44),
.A2(n_53),
.B1(n_55),
.B2(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_44),
.A2(n_55),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_45),
.A2(n_48),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_45),
.A2(n_48),
.B1(n_103),
.B2(n_170),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_80),
.Y(n_79)
);

OAI32xp33_ASAP7_75t_L g248 ( 
.A1(n_49),
.A2(n_63),
.A3(n_80),
.B1(n_241),
.B2(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_50),
.B(n_139),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_71),
.B2(n_74),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_66),
.B1(n_67),
.B2(n_97),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_63),
.B1(n_68),
.B2(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_62),
.B(n_250),
.Y(n_249)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_65),
.A2(n_74),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_65),
.A2(n_74),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_67),
.B1(n_72),
.B2(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_67),
.B(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_66),
.A2(n_67),
.B1(n_97),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_66),
.A2(n_67),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_66),
.A2(n_67),
.B1(n_197),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_66),
.A2(n_67),
.B1(n_135),
.B2(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_67),
.B(n_139),
.Y(n_224)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_88),
.B(n_90),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_88),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_82),
.B1(n_128),
.B2(n_131),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_78),
.A2(n_82),
.B1(n_131),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_78),
.A2(n_82),
.B1(n_153),
.B2(n_239),
.Y(n_238)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_80),
.Y(n_250)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_90),
.B(n_106),
.CI(n_118),
.CON(n_105),
.SN(n_105)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_91),
.A2(n_92),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.C(n_102),
.Y(n_92)
);

FAx1_ASAP7_75t_L g278 ( 
.A(n_93),
.B(n_98),
.CI(n_102),
.CON(n_278),
.SN(n_278)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_94),
.B(n_96),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_173),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_101),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_100),
.A2(n_101),
.B1(n_129),
.B2(n_152),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g295 ( 
.A(n_105),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_117),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_114),
.Y(n_116)
);

AOI321xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_276),
.A3(n_284),
.B1(n_289),
.B2(n_294),
.C(n_298),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_175),
.C(n_187),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_157),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_123),
.B(n_157),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_142),
.C(n_149),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_124),
.B(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_137),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_133),
.C(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_139),
.B(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_142),
.A2(n_149),
.B1(n_150),
.B2(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_142),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_156),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_151),
.B(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_154),
.B(n_156),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_155),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_165),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_164),
.C(n_165),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_162),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_174),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_171),
.C(n_174),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_176),
.A2(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_177),
.B(n_178),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_186),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_180),
.B(n_181),
.C(n_186),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_182),
.B(n_184),
.C(n_185),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_270),
.B(n_275),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_256),
.B(n_269),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_234),
.B(n_255),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_213),
.B(n_233),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_202),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_192),
.B(n_202),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_193),
.A2(n_194),
.B1(n_198),
.B2(n_199),
.Y(n_219)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_196),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_209),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_207),
.C(n_209),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_220),
.B(n_232),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_219),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_225),
.B(n_231),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_222),
.B(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_235),
.B(n_236),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_247),
.B1(n_253),
.B2(n_254),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_237)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_246),
.C(n_254),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_244),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_247),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_251),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_258),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_265),
.C(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_268),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_281),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.C(n_280),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_278),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_285),
.A2(n_290),
.B(n_293),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_286),
.B(n_287),
.Y(n_293)
);


endmodule