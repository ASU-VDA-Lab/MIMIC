module fake_jpeg_4005_n_230 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_40),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_24),
.B1(n_14),
.B2(n_16),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_55),
.B1(n_59),
.B2(n_20),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_35),
.A2(n_24),
.B1(n_14),
.B2(n_27),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_19),
.B1(n_15),
.B2(n_22),
.Y(n_70)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_51),
.Y(n_61)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_16),
.B(n_29),
.C(n_24),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_32),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_17),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_17),
.B(n_26),
.C(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_31),
.A2(n_14),
.B1(n_29),
.B2(n_28),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_21),
.B1(n_15),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_76),
.B1(n_55),
.B2(n_52),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_68),
.B(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_49),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_65),
.Y(n_104)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_70),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_74),
.Y(n_93)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_18),
.B1(n_17),
.B2(n_37),
.Y(n_75)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_50),
.B1(n_54),
.B2(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_18),
.B1(n_23),
.B2(n_33),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_50),
.C(n_47),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_23),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_56),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_66),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_103),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_90),
.A2(n_45),
.B1(n_47),
.B2(n_42),
.Y(n_120)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_69),
.B(n_23),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_48),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_96),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_116),
.Y(n_128)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_75),
.B(n_79),
.C(n_37),
.D(n_33),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_89),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_42),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_125),
.C(n_86),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_42),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_72),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_72),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_66),
.B1(n_74),
.B2(n_58),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_102),
.B(n_93),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_78),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_101),
.B(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_134),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_90),
.B1(n_67),
.B2(n_83),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_87),
.Y(n_135)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_137),
.B(n_139),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_98),
.B(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_145),
.Y(n_157)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_90),
.B1(n_99),
.B2(n_92),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_91),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_93),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_125),
.C(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_107),
.C(n_108),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_131),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_149),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_114),
.B1(n_111),
.B2(n_105),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_158),
.B1(n_130),
.B2(n_129),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_107),
.B1(n_113),
.B2(n_121),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_156),
.A2(n_45),
.B1(n_57),
.B2(n_65),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_107),
.B1(n_117),
.B2(n_66),
.Y(n_158)
);

XNOR2x1_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_57),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_45),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_140),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

AOI32xp33_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_137),
.A3(n_136),
.B1(n_128),
.B2(n_141),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_135),
.B(n_131),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_166),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_153),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_144),
.B1(n_130),
.B2(n_143),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_176),
.B1(n_152),
.B2(n_160),
.Y(n_182)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_173),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_172),
.C(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_151),
.A2(n_104),
.B(n_69),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_175),
.A2(n_177),
.B(n_162),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_57),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_189),
.C(n_190),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_182),
.A2(n_188),
.B1(n_185),
.B2(n_183),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

AOI31xp67_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_159),
.A3(n_156),
.B(n_157),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_176),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_162),
.B1(n_147),
.B2(n_148),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_23),
.C(n_26),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_81),
.C(n_26),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_81),
.C(n_26),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_174),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_181),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_192),
.A2(n_5),
.B(n_12),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_4),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_199),
.B1(n_5),
.B2(n_12),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_179),
.A2(n_164),
.B1(n_178),
.B2(n_168),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_0),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_175),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_6),
.Y(n_201)
);

OAI221xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_190),
.B1(n_6),
.B2(n_7),
.C(n_13),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_205),
.A2(n_206),
.B(n_210),
.Y(n_213)
);

OAI221xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_5),
.B1(n_12),
.B2(n_10),
.C(n_8),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_4),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_202),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_215),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_198),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_213),
.B(n_195),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_201),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_4),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_7),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_195),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_220),
.B(n_10),
.Y(n_225)
);

NOR4xp25_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_222),
.C(n_13),
.D(n_1),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_214),
.B(n_213),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_223),
.A2(n_224),
.B(n_225),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_227),
.C(n_0),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_3),
.Y(n_230)
);


endmodule