module fake_jpeg_16378_n_133 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_133);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_133;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_27),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_2),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_59),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_60),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_49),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_66),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_50),
.B1(n_44),
.B2(n_45),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_50),
.B1(n_46),
.B2(n_52),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_49),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_43),
.B1(n_53),
.B2(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_48),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_47),
.B1(n_1),
.B2(n_3),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_7),
.B1(n_9),
.B2(n_39),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_4),
.Y(n_79)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_4),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_5),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_91),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_11),
.B1(n_13),
.B2(n_15),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_10),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_92),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_86),
.B(n_24),
.Y(n_102)
);

XOR2x1_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_89),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_25),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_99),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_111),
.B(n_91),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_112),
.B(n_94),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_114),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_77),
.B1(n_80),
.B2(n_88),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_106),
.B1(n_102),
.B2(n_90),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_122),
.C(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_123),
.B(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_120),
.Y(n_127)
);

AOI21x1_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_118),
.B(n_33),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_93),
.B(n_34),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_31),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_35),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_36),
.Y(n_133)
);


endmodule