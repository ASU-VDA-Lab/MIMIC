module fake_jpeg_14400_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_21),
.Y(n_22)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_13),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_12),
.C(n_9),
.Y(n_33)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_33),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_15),
.B(n_14),
.C(n_12),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_26),
.B(n_9),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_17),
.B1(n_15),
.B2(n_11),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_32),
.B1(n_9),
.B2(n_0),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_21),
.B1(n_18),
.B2(n_14),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_24),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_36),
.C(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_38),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_30),
.B(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_34),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_0),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_47),
.B(n_46),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.C(n_45),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_41),
.B(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_42),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_7),
.Y(n_52)
);


endmodule