module real_jpeg_1110_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_2),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_2),
.A2(n_24),
.B1(n_44),
.B2(n_45),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_2),
.A2(n_24),
.B1(n_55),
.B2(n_56),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_20),
.B1(n_21),
.B2(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_3),
.A2(n_34),
.B1(n_55),
.B2(n_56),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_26),
.C(n_30),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_3),
.B(n_28),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_3),
.B(n_41),
.C(n_45),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_3),
.B(n_94),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_53),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_3),
.B(n_54),
.C(n_56),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_3),
.B(n_47),
.Y(n_234)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_37),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_6),
.A2(n_37),
.B1(n_55),
.B2(n_56),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_113)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_10),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_84),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_82),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_68),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_15),
.B(n_68),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_61),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_35),
.C(n_50),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_17),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_17),
.A2(n_70),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_17),
.A2(n_70),
.B1(n_144),
.B2(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_17),
.B(n_144),
.C(n_154),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g75 ( 
.A1(n_19),
.A2(n_63),
.B(n_65),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_26),
.Y(n_27)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_21),
.B(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_25),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_30),
.B(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_33),
.B(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_35),
.A2(n_50),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_35),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_35)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_38),
.A2(n_47),
.B1(n_105),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_39),
.A2(n_43),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

AOI22x1_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_45),
.B1(n_54),
.B2(n_57),
.Y(n_59)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_45),
.B(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g104 ( 
.A1(n_47),
.A2(n_80),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_75),
.C(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_50),
.A2(n_74),
.B1(n_77),
.B2(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_60),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_58),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_52),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_52),
.A2(n_58),
.B1(n_100),
.B2(n_101),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_52),
.A2(n_58),
.B(n_101),
.Y(n_170)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_53),
.A2(n_60),
.B1(n_116),
.B2(n_143),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_56),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B(n_65),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_63),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_75),
.C(n_76),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_69),
.A2(n_75),
.B1(n_127),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_69),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_70),
.B(n_89),
.C(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_75),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_75),
.A2(n_127),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_75),
.A2(n_126),
.B1(n_127),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_75),
.A2(n_127),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_76),
.B(n_272),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_77),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_258),
.B(n_275),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_148),
.B(n_257),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_128),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_87),
.B(n_128),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_107),
.C(n_118),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_88),
.B(n_107),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_102),
.B2(n_103),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_98),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_91),
.A2(n_98),
.B1(n_99),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_91),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_93),
.A2(n_94),
.B1(n_123),
.B2(n_160),
.Y(n_159)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_95),
.A2(n_96),
.B(n_122),
.Y(n_121)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_96),
.A2(n_122),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_98),
.A2(n_99),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_98),
.A2(n_99),
.B1(n_207),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_99),
.B(n_202),
.C(n_207),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_99),
.B(n_159),
.C(n_234),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_104),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_127),
.C(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_104),
.A2(n_106),
.B1(n_170),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_104),
.A2(n_106),
.B1(n_124),
.B2(n_125),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_104),
.B(n_124),
.C(n_241),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_117),
.Y(n_107)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_117),
.B1(n_136),
.B2(n_139),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_110),
.B(n_123),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_117),
.A2(n_132),
.B(n_139),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_118),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.C(n_127),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_119),
.A2(n_120),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_167),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_121),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_124),
.A2(n_125),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_124),
.B(n_228),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_147),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_140),
.B2(n_141),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_131),
.B(n_140),
.C(n_147),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_144),
.B(n_146),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_144),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_178),
.C(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_144),
.A2(n_162),
.B1(n_203),
.B2(n_206),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_146),
.A2(n_262),
.B1(n_266),
.B2(n_267),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_146),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_252),
.B(n_256),
.Y(n_148)
);

OAI211xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_181),
.B(n_195),
.C(n_251),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_171),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_171),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_163),
.B2(n_164),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_166),
.C(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_161),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_158),
.A2(n_159),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_159),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_159),
.B(n_222),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_170),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_177),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_177),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_179),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_SL g195 ( 
.A(n_182),
.B(n_196),
.C(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_183),
.B(n_184),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_185),
.B(n_187),
.C(n_193),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_193),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_213),
.B(n_250),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_199),
.B(n_201),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_244),
.B(n_249),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_238),
.B(n_243),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_230),
.B(n_237),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_224),
.B(n_229),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_221),
.B(n_223),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_236),
.Y(n_237)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_248),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_254),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_270),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_269),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_269),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_274),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_274),
.Y(n_277)
);


endmodule