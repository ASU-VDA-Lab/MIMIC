module real_jpeg_14210_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx10_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_2),
.A2(n_22),
.B1(n_29),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_3),
.A2(n_37),
.B1(n_43),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_61),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_3),
.A2(n_22),
.B1(n_29),
.B2(n_61),
.Y(n_110)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_5),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_5),
.A2(n_28),
.B1(n_37),
.B2(n_43),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_7),
.A2(n_37),
.B1(n_43),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_22),
.B1(n_29),
.B2(n_63),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_9),
.A2(n_22),
.B1(n_29),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_10),
.A2(n_34),
.B(n_49),
.C(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_10),
.B(n_73),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_10),
.A2(n_43),
.B(n_56),
.C(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_10),
.B(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_10),
.B(n_26),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_10),
.B(n_85),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_11),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_11),
.A2(n_22),
.B1(n_29),
.B2(n_46),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_12),
.Y(n_76)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_90),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_88),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_64),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_17),
.B(n_64),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_44),
.C(n_52),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_18),
.B(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_32),
.B2(n_33),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_20),
.B(n_32),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_21),
.A2(n_26),
.B1(n_30),
.B2(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_21),
.A2(n_26),
.B1(n_27),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_21),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_21),
.A2(n_26),
.B1(n_40),
.B2(n_118),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_21),
.A2(n_26),
.B1(n_110),
.B2(n_118),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_22),
.A2(n_29),
.B1(n_56),
.B2(n_57),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_22),
.B(n_120),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_25),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_29),
.A2(n_40),
.B(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI32xp33_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.A3(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_42),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_34),
.A2(n_35),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_40),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_44),
.B(n_52),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_48),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_58),
.B1(n_59),
.B2(n_62),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_85),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_54),
.A2(n_60),
.B1(n_85),
.B2(n_97),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_80),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_127),
.B(n_131),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_106),
.B(n_126),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_100),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_93),
.B(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_98),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_103),
.C(n_104),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_115),
.B(n_125),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_113),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_121),
.B(n_124),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_122),
.B(n_123),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_129),
.Y(n_131)
);


endmodule