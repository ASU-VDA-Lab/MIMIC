module fake_jpeg_29712_n_57 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_57);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_57;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_7),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_22),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_21),
.C(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_15),
.B1(n_14),
.B2(n_2),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_33),
.B1(n_27),
.B2(n_28),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_24),
.B1(n_1),
.B2(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_24),
.B1(n_4),
.B2(n_5),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_11),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_12),
.Y(n_47)
);

OAI322xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_29),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_6),
.C2(n_12),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_46),
.B1(n_39),
.B2(n_40),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_48),
.B(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_13),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_44),
.B1(n_47),
.B2(n_43),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_49),
.C(n_51),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_53),
.Y(n_57)
);


endmodule