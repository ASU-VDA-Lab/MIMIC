module real_jpeg_22425_n_17 (n_8, n_0, n_2, n_10, n_9, n_350, n_12, n_349, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_350;
input n_12;
input n_349;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_46),
.B1(n_49),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_1),
.A2(n_65),
.B1(n_66),
.B2(n_89),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_89),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_89),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_2),
.A2(n_22),
.B1(n_31),
.B2(n_32),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_2),
.A2(n_22),
.B1(n_65),
.B2(n_66),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_2),
.A2(n_22),
.B1(n_46),
.B2(n_49),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_3),
.A2(n_46),
.B1(n_49),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_3),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_101),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_101),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_3),
.A2(n_23),
.B1(n_25),
.B2(n_101),
.Y(n_216)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_5),
.A2(n_23),
.B1(n_25),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_5),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_5),
.A2(n_46),
.B1(n_49),
.B2(n_56),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_56),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_6),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_6),
.A2(n_46),
.B1(n_49),
.B2(n_106),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_106),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_106),
.Y(n_247)
);

A2O1A1O1Ixp25_ASAP7_75t_L g85 ( 
.A1(n_7),
.A2(n_49),
.B(n_61),
.C(n_86),
.D(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_7),
.B(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_45),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_7),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_7),
.A2(n_107),
.B(n_109),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_7),
.A2(n_31),
.B(n_42),
.C(n_145),
.D(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_7),
.B(n_31),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_7),
.B(n_35),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_7),
.A2(n_32),
.B(n_189),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_125),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_8),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_8),
.A2(n_46),
.B1(n_49),
.B2(n_58),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_58),
.Y(n_282)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_10),
.B(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_10),
.A2(n_129),
.B(n_155),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_11),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_11),
.A2(n_46),
.B1(n_49),
.B2(n_157),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_157),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_157),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_13),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_14),
.A2(n_23),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_34),
.B1(n_46),
.B2(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_14),
.A2(n_34),
.B1(n_65),
.B2(n_66),
.Y(n_236)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

AO21x1_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_342),
.B(n_345),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_75),
.B(n_341),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_20),
.B(n_36),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_20),
.B(n_343),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_20),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_33),
.B2(n_35),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_21),
.A2(n_26),
.B1(n_35),
.B2(n_71),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_23),
.A2(n_28),
.B(n_125),
.C(n_188),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_26),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_26),
.B(n_208),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_26),
.A2(n_33),
.B(n_35),
.Y(n_344)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_27),
.A2(n_30),
.B1(n_55),
.B2(n_57),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_27),
.A2(n_30),
.B1(n_216),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_27),
.A2(n_207),
.B(n_247),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_27),
.A2(n_30),
.B1(n_55),
.B2(n_291),
.Y(n_311)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_28),
.Y(n_189)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_30),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_30),
.A2(n_217),
.B(n_291),
.Y(n_290)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_35),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_70),
.C(n_72),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_37),
.A2(n_38),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_53),
.C(n_59),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_39),
.A2(n_40),
.B1(n_59),
.B2(n_316),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_41),
.A2(n_51),
.B1(n_166),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_41),
.A2(n_202),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_41),
.A2(n_50),
.B1(n_51),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_45),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_42),
.B(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_42),
.A2(n_45),
.B1(n_244),
.B2(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_42),
.A2(n_45),
.B1(n_263),
.B2(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_44),
.Y(n_153)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_46),
.B(n_48),
.Y(n_152)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_49),
.A2(n_145),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_51),
.B(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_51),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_51),
.A2(n_167),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_53),
.A2(n_54),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_59),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_59),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_68),
.B(n_69),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_60),
.A2(n_68),
.B1(n_100),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_60),
.A2(n_143),
.B(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_60),
.A2(n_68),
.B1(n_199),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_60),
.A2(n_68),
.B1(n_229),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_60),
.A2(n_68),
.B1(n_238),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_61),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_61),
.A2(n_64),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_65),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_66),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_68),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_68),
.A2(n_102),
.B(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_69),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_70),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_334),
.B(n_340),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_307),
.A3(n_327),
.B1(n_332),
.B2(n_333),
.C(n_349),
.Y(n_76)
);

AOI321xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_255),
.A3(n_295),
.B1(n_301),
.B2(n_306),
.C(n_350),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_210),
.C(n_251),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_181),
.B(n_209),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_160),
.B(n_180),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_137),
.B(n_159),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_112),
.B(n_136),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_94),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_84),
.B(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_85),
.A2(n_90),
.B1(n_91),
.B2(n_121),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_87),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_99),
.C(n_104),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_107),
.B(n_109),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_105),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_107),
.A2(n_108),
.B1(n_156),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_107),
.A2(n_127),
.B1(n_171),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_107),
.A2(n_192),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_107),
.A2(n_108),
.B1(n_227),
.B2(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_107),
.A2(n_108),
.B(n_236),
.Y(n_268)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_122),
.B(n_135),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_120),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_120),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_130),
.B(n_134),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_126),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_127),
.Y(n_133)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_127),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_139),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_150),
.B2(n_158),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_142),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_144),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_149),
.C(n_158),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_150),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_161),
.B(n_162),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_176),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_177),
.C(n_178),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_169),
.B2(n_175),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_172),
.C(n_173),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_172),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_182),
.B(n_183),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_196),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_185),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_185),
.B(n_195),
.C(n_196),
.Y(n_252)
);

AOI22x1_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_191),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_204),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_198),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_200),
.B(n_203),
.C(n_204),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_211),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_231),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_212),
.B(n_231),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_223),
.C(n_230),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_222),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_215),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_230),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_228),
.Y(n_240)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_249),
.B2(n_250),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_239),
.C(n_250),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_237),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_245),
.C(n_248),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_245),
.B1(n_246),
.B2(n_248),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_242),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_253),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_273),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_256),
.B(n_273),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.C(n_272),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_257),
.A2(n_258),
.B1(n_266),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_262),
.C(n_264),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_271),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_268),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_286),
.B(n_290),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_269),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_269),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_270),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_293),
.B2(n_294),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_284),
.B2(n_285),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_285),
.C(n_294),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_281),
.B(n_283),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_281),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_282),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_283),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_283),
.A2(n_309),
.B1(n_318),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_292),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_288),
.Y(n_292)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_302),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_320),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_320),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_318),
.C(n_319),
.Y(n_308)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_311),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_316),
.C(n_317),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_311),
.B(n_322),
.C(n_326),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_314),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_339),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_336),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_344),
.B(n_347),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_346),
.Y(n_345)
);


endmodule