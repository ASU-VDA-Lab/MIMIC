module fake_ariane_1394_n_734 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_734);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_734;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_672;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_658;
wire n_705;
wire n_630;
wire n_617;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_708;
wire n_308;
wire n_551;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_664;
wire n_629;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_29),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_49),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_93),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_18),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

BUFx8_ASAP7_75t_SL g164 ( 
.A(n_113),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_13),
.B(n_3),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_119),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_22),
.Y(n_167)
);

INVxp33_ASAP7_75t_SL g168 ( 
.A(n_90),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_52),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_102),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_149),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_3),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_36),
.Y(n_173)
);

NOR2xp67_ASAP7_75t_L g174 ( 
.A(n_73),
.B(n_136),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_74),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_115),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_11),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_30),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_55),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_59),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_80),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_13),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_128),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_28),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_122),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_14),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_127),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_131),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_91),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_100),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_67),
.Y(n_195)
);

BUFx8_ASAP7_75t_SL g196 ( 
.A(n_110),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_61),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_85),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_33),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_89),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_17),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_27),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_56),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_81),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_160),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_0),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_0),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

CKINVDCx6p67_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_180),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_1),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_156),
.B(n_1),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_2),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_182),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_4),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_5),
.Y(n_232)
);

NOR2x1_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_19),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_6),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_165),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_174),
.B(n_20),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_6),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_154),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_179),
.B(n_7),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_161),
.Y(n_246)
);

OAI21x1_ASAP7_75t_L g247 ( 
.A1(n_181),
.A2(n_77),
.B(n_151),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_169),
.B(n_7),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

AND2x4_ASAP7_75t_L g250 ( 
.A(n_181),
.B(n_8),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_181),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_220),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_214),
.B(n_168),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_248),
.B(n_166),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_195),
.B1(n_199),
.B2(n_196),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_224),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_230),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_214),
.B(n_248),
.Y(n_266)
);

NAND2xp33_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_202),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_245),
.B(n_167),
.Y(n_268)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_202),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_245),
.B(n_170),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_238),
.A2(n_191),
.B1(n_207),
.B2(n_171),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_175),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g279 ( 
.A(n_250),
.B(n_202),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_219),
.Y(n_280)
);

OR2x6_ASAP7_75t_L g281 ( 
.A(n_227),
.B(n_164),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_211),
.B(n_8),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_225),
.A2(n_208),
.B1(n_202),
.B2(n_201),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_212),
.Y(n_285)
);

BUFx4f_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_178),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_219),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_L g289 ( 
.A(n_216),
.B(n_208),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_225),
.A2(n_208),
.B1(n_200),
.B2(n_197),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_243),
.B(n_183),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_213),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_208),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_209),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_229),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_235),
.B(n_184),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_186),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g298 ( 
.A(n_213),
.B(n_240),
.Y(n_298)
);

NOR2x1p5_ASAP7_75t_L g299 ( 
.A(n_220),
.B(n_192),
.Y(n_299)
);

NAND3xp33_ASAP7_75t_L g300 ( 
.A(n_228),
.B(n_193),
.C(n_10),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_286),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_241),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_217),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_265),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_221),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_SL g306 ( 
.A(n_259),
.B(n_223),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_232),
.B1(n_226),
.B2(n_234),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_229),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_295),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_255),
.Y(n_312)
);

OAI221xp5_ASAP7_75t_L g313 ( 
.A1(n_290),
.A2(n_221),
.B1(n_236),
.B2(n_222),
.C(n_233),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_236),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_236),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_292),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_252),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_252),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_269),
.B(n_215),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_288),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_290),
.A2(n_239),
.B1(n_222),
.B2(n_215),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_257),
.B(n_215),
.Y(n_322)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_269),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_296),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_237),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_287),
.Y(n_329)
);

BUFx12f_ASAP7_75t_SL g330 ( 
.A(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_237),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_297),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_257),
.B(n_222),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_212),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_274),
.B(n_212),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_259),
.B(n_231),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_284),
.B(n_212),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_242),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_284),
.B(n_247),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_268),
.B(n_231),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_268),
.B(n_231),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_253),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_242),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_254),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_254),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_293),
.B(n_242),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_258),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_293),
.B(n_242),
.Y(n_351)
);

O2A1O1Ixp33_ASAP7_75t_L g352 ( 
.A1(n_272),
.A2(n_9),
.B(n_12),
.C(n_14),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_258),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_261),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_272),
.B(n_251),
.Y(n_355)
);

AOI221xp5_ASAP7_75t_L g356 ( 
.A1(n_298),
.A2(n_251),
.B1(n_12),
.B2(n_15),
.C(n_16),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_266),
.B(n_247),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_261),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_256),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_262),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_262),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_21),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_263),
.B(n_251),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_263),
.B(n_251),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_329),
.A2(n_281),
.B1(n_231),
.B2(n_277),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g367 ( 
.A1(n_306),
.A2(n_289),
.B(n_267),
.C(n_282),
.Y(n_367)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

AOI21x1_ASAP7_75t_L g369 ( 
.A1(n_342),
.A2(n_282),
.B(n_275),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_317),
.Y(n_370)
);

O2A1O1Ixp5_ASAP7_75t_L g371 ( 
.A1(n_303),
.A2(n_277),
.B(n_276),
.C(n_275),
.Y(n_371)
);

O2A1O1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_308),
.A2(n_281),
.B(n_270),
.C(n_271),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_331),
.A2(n_285),
.B(n_264),
.Y(n_373)
);

O2A1O1Ixp33_ASAP7_75t_L g374 ( 
.A1(n_352),
.A2(n_276),
.B(n_271),
.C(n_270),
.Y(n_374)
);

NAND2x1p5_ASAP7_75t_L g375 ( 
.A(n_305),
.B(n_251),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_336),
.A2(n_83),
.B(n_148),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_333),
.A2(n_82),
.B(n_147),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_326),
.B(n_9),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_322),
.A2(n_78),
.B(n_145),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_312),
.B(n_152),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_324),
.A2(n_76),
.B(n_143),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_301),
.A2(n_75),
.B(n_142),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_301),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_383)
);

O2A1O1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_304),
.A2(n_18),
.B(n_23),
.C(n_24),
.Y(n_384)
);

O2A1O1Ixp5_ASAP7_75t_L g385 ( 
.A1(n_357),
.A2(n_25),
.B(n_26),
.C(n_31),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_302),
.A2(n_326),
.B1(n_310),
.B2(n_335),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_310),
.B(n_144),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_357),
.A2(n_355),
.B(n_309),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_320),
.B(n_32),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_314),
.B(n_140),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_355),
.A2(n_34),
.B(n_35),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_319),
.A2(n_37),
.B(n_38),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_338),
.B(n_39),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_319),
.A2(n_40),
.B(n_41),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_307),
.B(n_139),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_327),
.B(n_314),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_328),
.A2(n_43),
.B(n_44),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_327),
.B(n_45),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_328),
.A2(n_46),
.B(n_47),
.Y(n_403)
);

OR2x6_ASAP7_75t_L g404 ( 
.A(n_330),
.B(n_48),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_315),
.B(n_50),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_L g406 ( 
.A1(n_313),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_311),
.B(n_57),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_359),
.B(n_137),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_343),
.B(n_58),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_356),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_321),
.B(n_64),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_344),
.B(n_341),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_337),
.B(n_323),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_323),
.B(n_135),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_346),
.A2(n_65),
.B(n_66),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

AOI21x1_ASAP7_75t_L g418 ( 
.A1(n_349),
.A2(n_68),
.B(n_69),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_334),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_334),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_351),
.A2(n_71),
.B(n_72),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_345),
.B(n_84),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_339),
.A2(n_86),
.B(n_87),
.Y(n_425)
);

AOI21x1_ASAP7_75t_L g426 ( 
.A1(n_353),
.A2(n_88),
.B(n_92),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_354),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_332),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_360),
.A2(n_94),
.B(n_96),
.Y(n_429)
);

NAND3xp33_ASAP7_75t_SL g430 ( 
.A(n_347),
.B(n_97),
.C(n_98),
.Y(n_430)
);

AO21x1_ASAP7_75t_L g431 ( 
.A1(n_348),
.A2(n_99),
.B(n_101),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_386),
.B(n_358),
.Y(n_432)
);

AO32x2_ASAP7_75t_L g433 ( 
.A1(n_383),
.A2(n_362),
.A3(n_361),
.B1(n_340),
.B2(n_350),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_361),
.B1(n_364),
.B2(n_363),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_369),
.A2(n_103),
.B(n_104),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_371),
.A2(n_105),
.B(n_106),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_397),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_378),
.B(n_107),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_412),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_112),
.Y(n_440)
);

AOI31xp67_ASAP7_75t_L g441 ( 
.A1(n_424),
.A2(n_116),
.A3(n_118),
.B(n_120),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_387),
.A2(n_408),
.B(n_393),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_400),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_129),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_419),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_404),
.B(n_133),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_399),
.A2(n_130),
.B1(n_132),
.B2(n_365),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_372),
.Y(n_449)
);

AO31x2_ASAP7_75t_L g450 ( 
.A1(n_431),
.A2(n_398),
.A3(n_410),
.B(n_406),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_422),
.Y(n_451)
);

NOR2xp67_ASAP7_75t_L g452 ( 
.A(n_368),
.B(n_391),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g453 ( 
.A1(n_392),
.A2(n_405),
.B(n_379),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_377),
.A2(n_389),
.B(n_411),
.C(n_380),
.Y(n_454)
);

AO21x1_ASAP7_75t_L g455 ( 
.A1(n_416),
.A2(n_402),
.B(n_382),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_391),
.B(n_413),
.Y(n_456)
);

OAI21x1_ASAP7_75t_SL g457 ( 
.A1(n_384),
.A2(n_374),
.B(n_381),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_370),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_407),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_426),
.A2(n_425),
.B(n_376),
.Y(n_460)
);

AO31x2_ASAP7_75t_L g461 ( 
.A1(n_367),
.A2(n_428),
.A3(n_414),
.B(n_403),
.Y(n_461)
);

NAND2x1p5_ASAP7_75t_L g462 ( 
.A(n_368),
.B(n_366),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_368),
.B(n_366),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_373),
.A2(n_385),
.B(n_396),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_423),
.B(n_366),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_390),
.A2(n_423),
.B1(n_415),
.B2(n_375),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_390),
.A2(n_423),
.B1(n_394),
.B2(n_401),
.Y(n_467)
);

AO31x2_ASAP7_75t_L g468 ( 
.A1(n_429),
.A2(n_421),
.A3(n_418),
.B(n_430),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_371),
.A2(n_342),
.B(n_388),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_397),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

AOI21x1_ASAP7_75t_L g472 ( 
.A1(n_387),
.A2(n_342),
.B(n_369),
.Y(n_472)
);

A2O1A1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_372),
.A2(n_306),
.B(n_386),
.C(n_377),
.Y(n_473)
);

AOI21x1_ASAP7_75t_L g474 ( 
.A1(n_387),
.A2(n_342),
.B(n_369),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_397),
.Y(n_475)
);

NAND3xp33_ASAP7_75t_L g476 ( 
.A(n_386),
.B(n_329),
.C(n_259),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_369),
.A2(n_388),
.B(n_371),
.Y(n_477)
);

OAI21x1_ASAP7_75t_L g478 ( 
.A1(n_369),
.A2(n_388),
.B(n_371),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_397),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_386),
.B(n_305),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_369),
.A2(n_388),
.B(n_371),
.Y(n_481)
);

AOI211x1_ASAP7_75t_L g482 ( 
.A1(n_383),
.A2(n_308),
.B(n_388),
.C(n_216),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_371),
.A2(n_342),
.B(n_388),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_369),
.A2(n_388),
.B(n_371),
.Y(n_484)
);

AOI211x1_ASAP7_75t_L g485 ( 
.A1(n_383),
.A2(n_308),
.B(n_388),
.C(n_216),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_447),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_480),
.B(n_476),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_471),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_472),
.A2(n_474),
.B(n_484),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_458),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_459),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_477),
.A2(n_481),
.B(n_478),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_451),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_437),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_469),
.A2(n_483),
.B(n_460),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_432),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_456),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_454),
.A2(n_442),
.B(n_455),
.Y(n_498)
);

OAI221xp5_ASAP7_75t_L g499 ( 
.A1(n_473),
.A2(n_470),
.B1(n_475),
.B2(n_448),
.C(n_449),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_453),
.A2(n_435),
.B(n_464),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_444),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_440),
.A2(n_446),
.B1(n_448),
.B2(n_439),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_463),
.B(n_452),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_479),
.B(n_445),
.Y(n_504)
);

AOI221xp5_ASAP7_75t_L g505 ( 
.A1(n_482),
.A2(n_485),
.B1(n_479),
.B2(n_443),
.C(n_438),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_467),
.A2(n_457),
.B(n_436),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_482),
.B(n_485),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_466),
.A2(n_434),
.B(n_439),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_465),
.Y(n_510)
);

AO32x2_ASAP7_75t_L g511 ( 
.A1(n_433),
.A2(n_450),
.A3(n_441),
.B1(n_468),
.B2(n_452),
.Y(n_511)
);

AO21x2_ASAP7_75t_L g512 ( 
.A1(n_433),
.A2(n_450),
.B(n_468),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_462),
.A2(n_463),
.B(n_450),
.Y(n_513)
);

AO21x2_ASAP7_75t_L g514 ( 
.A1(n_433),
.A2(n_474),
.B(n_472),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_468),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_470),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_472),
.A2(n_474),
.B(n_477),
.Y(n_517)
);

CKINVDCx6p67_ASAP7_75t_R g518 ( 
.A(n_479),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_463),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_480),
.B(n_386),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_473),
.B(n_329),
.C(n_482),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_447),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_454),
.A2(n_473),
.B(n_469),
.Y(n_523)
);

AO21x2_ASAP7_75t_L g524 ( 
.A1(n_472),
.A2(n_474),
.B(n_442),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_451),
.Y(n_525)
);

A2O1A1Ixp33_ASAP7_75t_SL g526 ( 
.A1(n_464),
.A2(n_389),
.B(n_384),
.C(n_377),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_463),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_472),
.A2(n_474),
.B(n_442),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_L g529 ( 
.A1(n_473),
.A2(n_476),
.B(n_372),
.C(n_454),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_480),
.B(n_329),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_463),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_520),
.B(n_487),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_507),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_503),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_496),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_502),
.A2(n_530),
.B(n_529),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_509),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_527),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_503),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_513),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_487),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_486),
.Y(n_542)
);

BUFx5_ASAP7_75t_L g543 ( 
.A(n_497),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_519),
.Y(n_544)
);

AOI21x1_ASAP7_75t_L g545 ( 
.A1(n_498),
.A2(n_506),
.B(n_500),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_488),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_522),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_494),
.Y(n_548)
);

INVx4_ASAP7_75t_SL g549 ( 
.A(n_503),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_516),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_519),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_504),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_523),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_SL g554 ( 
.A(n_502),
.B(n_499),
.C(n_505),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_525),
.B(n_493),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_500),
.A2(n_495),
.B(n_489),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_527),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_521),
.B(n_512),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_490),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_508),
.B(n_531),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_491),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_515),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_529),
.A2(n_501),
.B1(n_518),
.B2(n_510),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_518),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_531),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_531),
.B(n_512),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_508),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_553),
.B(n_511),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_553),
.B(n_511),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_544),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_532),
.B(n_511),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_537),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_532),
.B(n_511),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_541),
.B(n_514),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_537),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_514),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_566),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_566),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_558),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_536),
.B(n_492),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_552),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_544),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_548),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_542),
.B(n_492),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_555),
.B(n_526),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_558),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_562),
.B(n_524),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_542),
.B(n_528),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_560),
.Y(n_589)
);

AO31x2_ASAP7_75t_L g590 ( 
.A1(n_540),
.A2(n_517),
.A3(n_562),
.B(n_533),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_546),
.B(n_547),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_538),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_546),
.B(n_547),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_554),
.B(n_561),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_533),
.B(n_535),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_549),
.B(n_534),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_559),
.B(n_565),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_567),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_564),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_571),
.B(n_567),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_572),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_571),
.B(n_543),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_577),
.B(n_549),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_577),
.B(n_549),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_590),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_543),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_583),
.B(n_595),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_592),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_578),
.B(n_563),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_572),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_575),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_597),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_590),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_575),
.Y(n_614)
);

AND2x4_ASAP7_75t_SL g615 ( 
.A(n_596),
.B(n_534),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_597),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_592),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_578),
.B(n_549),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_595),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_574),
.B(n_556),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_584),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_573),
.B(n_543),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_584),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_573),
.B(n_543),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_591),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_591),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_594),
.A2(n_538),
.B1(n_565),
.B2(n_539),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_588),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_576),
.B(n_543),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_588),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_576),
.B(n_556),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_568),
.B(n_543),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_627),
.B(n_585),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_619),
.B(n_607),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_612),
.B(n_587),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_601),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_606),
.B(n_594),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_601),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_610),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_600),
.B(n_569),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_600),
.B(n_602),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_602),
.B(n_569),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_610),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_622),
.B(n_568),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_603),
.B(n_589),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_622),
.B(n_580),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_616),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_625),
.B(n_593),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_611),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_608),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_626),
.B(n_593),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_613),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_611),
.Y(n_653)
);

AND2x4_ASAP7_75t_SL g654 ( 
.A(n_603),
.B(n_618),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_614),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_620),
.B(n_587),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_614),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_604),
.A2(n_596),
.B1(n_543),
.B2(n_599),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_636),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_638),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_637),
.B(n_630),
.Y(n_661)
);

NAND2x1p5_ASAP7_75t_L g662 ( 
.A(n_633),
.B(n_582),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_656),
.B(n_631),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_637),
.B(n_647),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_639),
.Y(n_665)
);

AND3x2_ASAP7_75t_L g666 ( 
.A(n_645),
.B(n_550),
.C(n_605),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_643),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_649),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_656),
.B(n_620),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_634),
.B(n_628),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_653),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_655),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_635),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_642),
.B(n_628),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_657),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_641),
.B(n_582),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_641),
.B(n_624),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_659),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_677),
.B(n_642),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_663),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_660),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_669),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_665),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_661),
.B(n_644),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_667),
.Y(n_685)
);

AOI222xp33_ASAP7_75t_L g686 ( 
.A1(n_673),
.A2(n_633),
.B1(n_605),
.B2(n_580),
.C1(n_579),
.C2(n_586),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_668),
.Y(n_687)
);

NOR2x1_ASAP7_75t_L g688 ( 
.A(n_683),
.B(n_664),
.Y(n_688)
);

NAND2x1_ASAP7_75t_L g689 ( 
.A(n_683),
.B(n_676),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_678),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_686),
.A2(n_662),
.B(n_684),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_686),
.A2(n_613),
.B1(n_618),
.B2(n_604),
.Y(n_692)
);

OAI21xp33_ASAP7_75t_SL g693 ( 
.A1(n_679),
.A2(n_674),
.B(n_673),
.Y(n_693)
);

OAI32xp33_ASAP7_75t_L g694 ( 
.A1(n_684),
.A2(n_662),
.A3(n_670),
.B1(n_609),
.B2(n_672),
.Y(n_694)
);

OAI211xp5_ASAP7_75t_L g695 ( 
.A1(n_691),
.A2(n_687),
.B(n_685),
.C(n_681),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_690),
.B(n_680),
.Y(n_696)
);

AOI221x1_ASAP7_75t_L g697 ( 
.A1(n_693),
.A2(n_675),
.B1(n_671),
.B2(n_682),
.C(n_613),
.Y(n_697)
);

OAI221xp5_ASAP7_75t_L g698 ( 
.A1(n_692),
.A2(n_658),
.B1(n_609),
.B2(n_651),
.C(n_648),
.Y(n_698)
);

NAND4xp25_ASAP7_75t_L g699 ( 
.A(n_694),
.B(n_650),
.C(n_623),
.D(n_621),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_689),
.Y(n_700)
);

NOR3xp33_ASAP7_75t_L g701 ( 
.A(n_695),
.B(n_688),
.C(n_652),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_696),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_700),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_699),
.B(n_644),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_702),
.B(n_698),
.Y(n_705)
);

AND4x1_ASAP7_75t_L g706 ( 
.A(n_701),
.B(n_697),
.C(n_640),
.D(n_646),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_703),
.B(n_646),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_707),
.B(n_705),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_706),
.B(n_704),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_706),
.B(n_570),
.C(n_617),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_708),
.B(n_631),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_710),
.B(n_650),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_709),
.B(n_640),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_708),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_708),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_714),
.Y(n_716)
);

OA22x2_ASAP7_75t_L g717 ( 
.A1(n_715),
.A2(n_666),
.B1(n_654),
.B2(n_650),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_713),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_711),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_712),
.Y(n_720)
);

OAI22xp5_ASAP7_75t_L g721 ( 
.A1(n_716),
.A2(n_621),
.B1(n_623),
.B2(n_654),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_719),
.B(n_624),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_718),
.B(n_632),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_717),
.Y(n_724)
);

AOI22x1_ASAP7_75t_L g725 ( 
.A1(n_724),
.A2(n_720),
.B1(n_617),
.B2(n_608),
.Y(n_725)
);

XNOR2xp5_ASAP7_75t_L g726 ( 
.A(n_723),
.B(n_551),
.Y(n_726)
);

OAI21xp5_ASAP7_75t_SL g727 ( 
.A1(n_722),
.A2(n_592),
.B(n_615),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_726),
.A2(n_721),
.B1(n_570),
.B2(n_598),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_727),
.A2(n_551),
.B1(n_632),
.B2(n_629),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_725),
.Y(n_730)
);

OAI21x1_ASAP7_75t_L g731 ( 
.A1(n_730),
.A2(n_565),
.B(n_545),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_731),
.B(n_728),
.Y(n_732)
);

OR2x6_ASAP7_75t_L g733 ( 
.A(n_732),
.B(n_729),
.Y(n_733)
);

OAI21xp5_ASAP7_75t_SL g734 ( 
.A1(n_733),
.A2(n_615),
.B(n_557),
.Y(n_734)
);


endmodule