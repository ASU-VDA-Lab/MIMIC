module fake_ariane_2501_n_1701 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1701);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1701;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_89),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_32),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_45),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_15),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_62),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_86),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_63),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_11),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_49),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_56),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_39),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_128),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_36),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_65),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_47),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_57),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_76),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_25),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_44),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_28),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_122),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_93),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_38),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_41),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_110),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_71),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_108),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_69),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_73),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_138),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_99),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_120),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_132),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_97),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_22),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_52),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_61),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_95),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_94),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_55),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_12),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_28),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_106),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_67),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_123),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_16),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_12),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_66),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_96),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_22),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_21),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_6),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_136),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_84),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_113),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_36),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_103),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_44),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_24),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_125),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_109),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_24),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_114),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_18),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_129),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_79),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_75),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_19),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_70),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_115),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_111),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_80),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_143),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_0),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_23),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_34),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_139),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_1),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_41),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_74),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_51),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_30),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_15),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_19),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_4),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_8),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_8),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_27),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_127),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_92),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_20),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_53),
.Y(n_260)
);

BUFx2_ASAP7_75t_SL g261 ( 
.A(n_26),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_11),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_17),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_141),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_43),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_85),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_4),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_10),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_100),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_37),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_1),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_39),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_23),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_40),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_82),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_30),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_144),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_43),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_42),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_149),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_17),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_5),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_104),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_45),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_116),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_121),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_98),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_20),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_101),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_25),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_38),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_107),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_7),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_34),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_10),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_102),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_59),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_64),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_126),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_37),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_68),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_140),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_46),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_152),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_29),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_160),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_160),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_262),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_153),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_158),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_271),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_227),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_189),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_179),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_221),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_168),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_161),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_161),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_192),
.B(n_0),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_182),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_173),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_183),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_183),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_178),
.B(n_2),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_173),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_211),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_184),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_213),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_184),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_224),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_229),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_235),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_226),
.B(n_2),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_242),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_230),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_246),
.B(n_3),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_250),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_183),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_251),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_230),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_178),
.B(n_249),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_174),
.B(n_3),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_252),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_254),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_255),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_263),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_285),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_185),
.B(n_6),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_285),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_223),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_183),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_177),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_183),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_223),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_272),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_223),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_186),
.B(n_9),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_278),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_273),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_R g365 ( 
.A(n_155),
.B(n_54),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_164),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_164),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_163),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_279),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_163),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_177),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_170),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_165),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_165),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_293),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_278),
.Y(n_376)
);

NOR2xp67_ASAP7_75t_L g377 ( 
.A(n_249),
.B(n_9),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_166),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_166),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_190),
.B(n_13),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_261),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_295),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_278),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_167),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_170),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_167),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_326),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_383),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_326),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_171),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_330),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_R g393 ( 
.A(n_368),
.B(n_187),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_330),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_308),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_383),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_352),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_327),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_328),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_328),
.B(n_175),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_352),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_343),
.B(n_197),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_354),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g404 ( 
.A1(n_347),
.A2(n_214),
.B(n_200),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_R g405 ( 
.A(n_370),
.B(n_188),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_354),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_312),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_314),
.B(n_259),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_306),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_376),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_376),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_307),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_313),
.B(n_259),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_321),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_322),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_317),
.B(n_288),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_320),
.B(n_288),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_358),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_370),
.B(n_373),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_323),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_332),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_325),
.B(n_201),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_334),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_318),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_SL g429 ( 
.A(n_316),
.B(n_256),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_333),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_340),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_381),
.B(n_175),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_345),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_336),
.B(n_291),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_339),
.B(n_291),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_342),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_344),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_373),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_348),
.B(n_278),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_350),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_R g446 ( 
.A(n_374),
.B(n_191),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_311),
.A2(n_256),
.B1(n_300),
.B2(n_294),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_351),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_374),
.Y(n_449)
);

CKINVDCx8_ASAP7_75t_R g450 ( 
.A(n_309),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_360),
.B(n_202),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_366),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_364),
.B(n_290),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_369),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_382),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_324),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_378),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_378),
.Y(n_458)
);

CKINVDCx8_ASAP7_75t_R g459 ( 
.A(n_309),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_346),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_456),
.B(n_355),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_310),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_402),
.Y(n_463)
);

INVx4_ASAP7_75t_SL g464 ( 
.A(n_399),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_456),
.B(n_379),
.Y(n_465)
);

INVx5_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_329),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_441),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_357),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_411),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_426),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_377),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_456),
.B(n_379),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_409),
.B(n_355),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_410),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_409),
.B(n_359),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_420),
.Y(n_478)
);

OR2x6_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_338),
.Y(n_479)
);

INVx4_ASAP7_75t_L g480 ( 
.A(n_441),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_441),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_410),
.Y(n_482)
);

NAND3xp33_ASAP7_75t_L g483 ( 
.A(n_422),
.B(n_386),
.C(n_384),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_456),
.B(n_384),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_426),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_393),
.B(n_386),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_430),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_405),
.B(n_310),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_410),
.Y(n_490)
);

NAND2x1p5_ASAP7_75t_L g491 ( 
.A(n_409),
.B(n_194),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_430),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_391),
.A2(n_319),
.B1(n_316),
.B2(n_341),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_421),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_440),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_440),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_428),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_437),
.B(n_428),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_421),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_447),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_441),
.B(n_359),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_446),
.B(n_442),
.Y(n_507)
);

BUFx10_ASAP7_75t_L g508 ( 
.A(n_449),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_457),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_443),
.B(n_200),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_396),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_458),
.B(n_315),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_448),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_417),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_416),
.B(n_315),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_395),
.B(n_361),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_387),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_396),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_396),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_423),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_433),
.B(n_319),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_448),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_395),
.B(n_375),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_395),
.B(n_353),
.Y(n_525)
);

BUFx4f_ASAP7_75t_L g526 ( 
.A(n_416),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_416),
.B(n_206),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_407),
.B(n_362),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_399),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_448),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_424),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_455),
.A2(n_380),
.B1(n_305),
.B2(n_300),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_407),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_455),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_452),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_435),
.B(n_438),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_455),
.A2(n_157),
.B1(n_268),
.B2(n_214),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_408),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_443),
.B(n_236),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_436),
.B(n_290),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_450),
.B(n_459),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_438),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_444),
.B(n_208),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_444),
.B(n_169),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_445),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_445),
.B(n_169),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_SL g547 ( 
.A(n_450),
.B(n_293),
.C(n_294),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_425),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_454),
.B(n_280),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_425),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_450),
.B(n_459),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_454),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_451),
.B(n_299),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_408),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_436),
.B(n_236),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_436),
.B(n_280),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_388),
.B(n_398),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_439),
.B(n_289),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_439),
.B(n_289),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_388),
.Y(n_560)
);

BUFx10_ASAP7_75t_L g561 ( 
.A(n_390),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_392),
.B(n_154),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_439),
.B(n_290),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_459),
.B(n_367),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_398),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_412),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_404),
.B(n_209),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_408),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_412),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_394),
.B(n_156),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_397),
.B(n_198),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_400),
.B(n_172),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_415),
.A2(n_278),
.B1(n_212),
.B2(n_304),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_413),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_415),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_415),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_400),
.B(n_172),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_418),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_418),
.B(n_176),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_418),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_401),
.Y(n_581)
);

BUFx10_ASAP7_75t_L g582 ( 
.A(n_403),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_427),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_404),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_404),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_460),
.B(n_419),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_419),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_419),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_406),
.B(n_232),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_460),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_R g591 ( 
.A(n_434),
.B(n_365),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_429),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_414),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_431),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_411),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_432),
.B(n_372),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_505),
.A2(n_385),
.B1(n_301),
.B2(n_297),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_465),
.B(n_205),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_468),
.B(n_480),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_548),
.B(n_176),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_550),
.B(n_180),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_499),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g603 ( 
.A(n_596),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_478),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_517),
.B(n_207),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_465),
.B(n_216),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_474),
.B(n_217),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_478),
.Y(n_609)
);

AND2x6_ASAP7_75t_SL g610 ( 
.A(n_479),
.B(n_234),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_529),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_553),
.A2(n_474),
.B1(n_477),
.B2(n_475),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_493),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_516),
.B(n_180),
.Y(n_614)
);

OAI22xp33_ASAP7_75t_L g615 ( 
.A1(n_505),
.A2(n_218),
.B1(n_303),
.B2(n_231),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_508),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_516),
.B(n_475),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_463),
.B(n_553),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_471),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_493),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_496),
.B(n_181),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_475),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_532),
.A2(n_258),
.B1(n_296),
.B2(n_244),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_468),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_496),
.B(n_238),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_504),
.Y(n_626)
);

BUFx5_ASAP7_75t_L g627 ( 
.A(n_555),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_480),
.B(n_238),
.Y(n_628)
);

AND2x2_ASAP7_75t_SL g629 ( 
.A(n_532),
.B(n_237),
.Y(n_629)
);

INVxp33_ASAP7_75t_L g630 ( 
.A(n_462),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_479),
.A2(n_264),
.B1(n_248),
.B2(n_257),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_479),
.A2(n_275),
.B1(n_239),
.B2(n_225),
.Y(n_632)
);

OAI221xp5_ASAP7_75t_L g633 ( 
.A1(n_537),
.A2(n_270),
.B1(n_241),
.B2(n_243),
.C(n_253),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_502),
.B(n_222),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_503),
.B(n_265),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_500),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_477),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_542),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_576),
.B(n_240),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_576),
.B(n_286),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_502),
.B(n_267),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_555),
.A2(n_282),
.B1(n_274),
.B2(n_276),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_506),
.B(n_286),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_470),
.B(n_284),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_481),
.B(n_287),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_545),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_461),
.A2(n_495),
.B1(n_484),
.B2(n_481),
.Y(n_647)
);

NOR2x1p5_ASAP7_75t_L g648 ( 
.A(n_531),
.B(n_292),
.Y(n_648)
);

NOR2xp67_ASAP7_75t_L g649 ( 
.A(n_483),
.B(n_298),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_501),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_508),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_511),
.Y(n_652)
);

AND2x6_ASAP7_75t_SL g653 ( 
.A(n_514),
.B(n_14),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_511),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_559),
.B(n_516),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_585),
.B(n_159),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_518),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_585),
.B(n_159),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_484),
.B(n_14),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_552),
.Y(n_660)
);

OAI221xp5_ASAP7_75t_L g661 ( 
.A1(n_537),
.A2(n_302),
.B1(n_283),
.B2(n_277),
.C(n_269),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_525),
.B(n_266),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_518),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_519),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_491),
.B(n_16),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_528),
.B(n_260),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_529),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_491),
.B(n_18),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_533),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_560),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_519),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_585),
.B(n_159),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_SL g673 ( 
.A1(n_514),
.A2(n_247),
.B1(n_233),
.B2(n_228),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_585),
.B(n_159),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_592),
.B(n_21),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_535),
.B(n_26),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_476),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_587),
.B(n_543),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_515),
.B(n_27),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_524),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_515),
.B(n_29),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_587),
.B(n_220),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_469),
.B(n_31),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_540),
.B(n_31),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_476),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_526),
.B(n_529),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_529),
.Y(n_687)
);

NOR3xp33_ASAP7_75t_L g688 ( 
.A(n_547),
.B(n_219),
.C(n_215),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_521),
.B(n_32),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_563),
.B(n_210),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_526),
.B(n_159),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_541),
.B(n_159),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_593),
.B(n_33),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_565),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_482),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_566),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_589),
.B(n_33),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_595),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_555),
.A2(n_159),
.B1(n_162),
.B2(n_199),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_555),
.A2(n_162),
.B1(n_203),
.B2(n_196),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_510),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_556),
.B(n_558),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_556),
.B(n_204),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_556),
.B(n_195),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_520),
.B(n_35),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_589),
.B(n_35),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_593),
.B(n_40),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_574),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_524),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_558),
.B(n_536),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_486),
.B(n_193),
.Y(n_711)
);

BUFx6f_ASAP7_75t_SL g712 ( 
.A(n_561),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_509),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_524),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_482),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_509),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_486),
.B(n_162),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_590),
.B(n_162),
.Y(n_718)
);

AND2x6_ASAP7_75t_SL g719 ( 
.A(n_595),
.B(n_162),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_569),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_561),
.B(n_48),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_581),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_490),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_549),
.B(n_50),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_564),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_541),
.A2(n_58),
.B1(n_60),
.B2(n_72),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_549),
.B(n_147),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_549),
.B(n_77),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_510),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_575),
.B(n_145),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_578),
.B(n_81),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_551),
.B(n_83),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_559),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_580),
.B(n_87),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_551),
.B(n_90),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_588),
.B(n_91),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_591),
.Y(n_737)
);

NOR3xp33_ASAP7_75t_L g738 ( 
.A(n_512),
.B(n_105),
.C(n_118),
.Y(n_738)
);

NOR3xp33_ASAP7_75t_L g739 ( 
.A(n_512),
.B(n_124),
.C(n_135),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_510),
.A2(n_137),
.B1(n_539),
.B2(n_467),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_581),
.B(n_582),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_569),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_567),
.A2(n_557),
.B(n_538),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_559),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_490),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_467),
.B(n_473),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_467),
.B(n_473),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_473),
.B(n_586),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_472),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_611),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_618),
.B(n_598),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_737),
.B(n_583),
.Y(n_752)
);

AOI21x1_ASAP7_75t_L g753 ( 
.A1(n_656),
.A2(n_584),
.B(n_534),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_598),
.B(n_507),
.C(n_557),
.Y(n_754)
);

AO32x1_ASAP7_75t_L g755 ( 
.A1(n_647),
.A2(n_584),
.A3(n_530),
.B1(n_485),
.B2(n_487),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_629),
.A2(n_573),
.B1(n_510),
.B2(n_539),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_607),
.B(n_586),
.Y(n_757)
);

O2A1O1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_607),
.A2(n_507),
.B(n_579),
.C(n_544),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_608),
.B(n_612),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_638),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_608),
.A2(n_546),
.B(n_489),
.C(n_570),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_646),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_660),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_630),
.B(n_562),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_602),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_658),
.A2(n_674),
.B(n_743),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_670),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_714),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_604),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_658),
.A2(n_522),
.B(n_568),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_748),
.B(n_539),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_678),
.B(n_539),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_611),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_694),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_659),
.A2(n_513),
.B(n_523),
.C(n_488),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_674),
.A2(n_522),
.B(n_554),
.Y(n_776)
);

AND2x6_ASAP7_75t_L g777 ( 
.A(n_740),
.B(n_498),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_701),
.Y(n_778)
);

AO21x1_ASAP7_75t_L g779 ( 
.A1(n_726),
.A2(n_497),
.B(n_494),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_SL g780 ( 
.A(n_729),
.B(n_582),
.Y(n_780)
);

CKINVDCx10_ASAP7_75t_R g781 ( 
.A(n_712),
.Y(n_781)
);

O2A1O1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_615),
.A2(n_489),
.B(n_571),
.C(n_492),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_710),
.B(n_573),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_603),
.B(n_594),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_679),
.A2(n_527),
.B(n_572),
.Y(n_785)
);

OAI21xp33_ASAP7_75t_L g786 ( 
.A1(n_606),
.A2(n_577),
.B(n_591),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_679),
.A2(n_466),
.B(n_464),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_629),
.A2(n_464),
.B1(n_466),
.B2(n_623),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_684),
.B(n_464),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_730),
.A2(n_466),
.B(n_731),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_628),
.A2(n_645),
.B(n_672),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_702),
.B(n_605),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_659),
.A2(n_706),
.B(n_697),
.C(n_681),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_696),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_636),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_623),
.A2(n_597),
.B1(n_631),
.B2(n_632),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_650),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_681),
.A2(n_720),
.B(n_742),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_655),
.B(n_680),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_714),
.B(n_709),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_611),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_619),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_698),
.B(n_617),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_SL g804 ( 
.A1(n_734),
.A2(n_736),
.B(n_726),
.C(n_686),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_609),
.B(n_613),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_620),
.B(n_626),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_615),
.A2(n_697),
.B(n_706),
.C(n_601),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_631),
.B(n_711),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_655),
.B(n_622),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_624),
.A2(n_691),
.B(n_662),
.Y(n_810)
);

AOI21x1_ASAP7_75t_L g811 ( 
.A1(n_691),
.A2(n_735),
.B(n_692),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_597),
.A2(n_632),
.B1(n_747),
.B2(n_746),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_666),
.A2(n_686),
.B(n_643),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_676),
.Y(n_814)
);

NOR2xp67_ASAP7_75t_L g815 ( 
.A(n_716),
.B(n_741),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_600),
.A2(n_682),
.B(n_717),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_711),
.B(n_708),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_637),
.B(n_690),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_642),
.B(n_729),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_749),
.Y(n_820)
);

INVx11_ASAP7_75t_L g821 ( 
.A(n_712),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_621),
.A2(n_625),
.B(n_640),
.Y(n_822)
);

INVx11_ASAP7_75t_L g823 ( 
.A(n_616),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_639),
.A2(n_689),
.B(n_633),
.C(n_614),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_725),
.B(n_733),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_689),
.A2(n_683),
.B(n_635),
.C(n_644),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_733),
.B(n_744),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_675),
.B(n_665),
.Y(n_828)
);

AO21x1_ASAP7_75t_L g829 ( 
.A1(n_735),
.A2(n_692),
.B(n_732),
.Y(n_829)
);

OAI321xp33_ASAP7_75t_L g830 ( 
.A1(n_665),
.A2(n_668),
.A3(n_705),
.B1(n_642),
.B2(n_700),
.C(n_699),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_616),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_744),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_675),
.B(n_668),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_705),
.A2(n_661),
.B(n_641),
.C(n_634),
.Y(n_834)
);

AO21x1_ASAP7_75t_L g835 ( 
.A1(n_738),
.A2(n_739),
.B(n_718),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_651),
.B(n_722),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_627),
.B(n_669),
.Y(n_837)
);

AO21x1_ASAP7_75t_L g838 ( 
.A1(n_724),
.A2(n_727),
.B(n_728),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_651),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_677),
.A2(n_745),
.B(n_723),
.Y(n_840)
);

AO21x1_ASAP7_75t_L g841 ( 
.A1(n_685),
.A2(n_715),
.B(n_695),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_611),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_669),
.A2(n_704),
.B(n_703),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_705),
.A2(n_688),
.B(n_693),
.C(n_707),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_SL g845 ( 
.A(n_722),
.B(n_713),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_699),
.A2(n_700),
.B(n_649),
.C(n_721),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_652),
.A2(n_664),
.B(n_671),
.Y(n_847)
);

NOR2x1_ASAP7_75t_L g848 ( 
.A(n_713),
.B(n_648),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_654),
.A2(n_663),
.B(n_657),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_701),
.B(n_627),
.Y(n_850)
);

NOR2xp67_ASAP7_75t_L g851 ( 
.A(n_667),
.B(n_687),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_627),
.B(n_667),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_701),
.B(n_627),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_667),
.A2(n_687),
.B1(n_673),
.B2(n_627),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_610),
.B(n_719),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_687),
.A2(n_584),
.B(n_743),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_653),
.B(n_326),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_598),
.A2(n_607),
.B1(n_608),
.B2(n_631),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_602),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_638),
.Y(n_860)
);

OAI21xp33_ASAP7_75t_L g861 ( 
.A1(n_598),
.A2(n_608),
.B(n_607),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_638),
.Y(n_862)
);

AND2x6_ASAP7_75t_L g863 ( 
.A(n_740),
.B(n_655),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_612),
.B(n_618),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_714),
.B(n_505),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_714),
.Y(n_866)
);

AOI21x1_ASAP7_75t_L g867 ( 
.A1(n_656),
.A2(n_674),
.B(n_658),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_714),
.Y(n_868)
);

AO21x1_ASAP7_75t_L g869 ( 
.A1(n_726),
.A2(n_735),
.B(n_681),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_599),
.A2(n_618),
.B(n_656),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_618),
.B(n_548),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_599),
.A2(n_618),
.B(n_656),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_612),
.B(n_618),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_743),
.A2(n_584),
.B(n_567),
.Y(n_874)
);

O2A1O1Ixp5_ASAP7_75t_L g875 ( 
.A1(n_598),
.A2(n_608),
.B(n_607),
.C(n_656),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_618),
.B(n_548),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_598),
.A2(n_607),
.B1(n_608),
.B2(n_631),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_618),
.B(n_548),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_612),
.B(n_618),
.Y(n_879)
);

AO22x1_ASAP7_75t_L g880 ( 
.A1(n_698),
.A2(n_505),
.B1(n_330),
.B2(n_352),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_619),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_598),
.A2(n_608),
.B(n_607),
.C(n_659),
.Y(n_882)
);

BUFx4f_ASAP7_75t_L g883 ( 
.A(n_655),
.Y(n_883)
);

OAI21x1_ASAP7_75t_L g884 ( 
.A1(n_743),
.A2(n_584),
.B(n_656),
.Y(n_884)
);

BUFx8_ASAP7_75t_L g885 ( 
.A(n_712),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_618),
.B(n_548),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_714),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_599),
.A2(n_618),
.B(n_656),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_612),
.A2(n_618),
.B1(n_607),
.B2(n_608),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_618),
.B(n_548),
.Y(n_890)
);

O2A1O1Ixp5_ASAP7_75t_L g891 ( 
.A1(n_598),
.A2(n_608),
.B(n_607),
.C(n_656),
.Y(n_891)
);

AOI21x1_ASAP7_75t_L g892 ( 
.A1(n_656),
.A2(n_674),
.B(n_658),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_598),
.A2(n_608),
.B(n_607),
.C(n_659),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_618),
.B(n_548),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_618),
.B(n_548),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_599),
.A2(n_618),
.B(n_656),
.Y(n_896)
);

NAND2x1p5_ASAP7_75t_L g897 ( 
.A(n_729),
.B(n_655),
.Y(n_897)
);

CKINVDCx8_ASAP7_75t_R g898 ( 
.A(n_619),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_599),
.A2(n_618),
.B(n_656),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_714),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_737),
.B(n_326),
.Y(n_901)
);

OAI21xp33_ASAP7_75t_L g902 ( 
.A1(n_598),
.A2(n_608),
.B(n_607),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_701),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_737),
.B(n_326),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_618),
.B(n_548),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_598),
.A2(n_607),
.B1(n_608),
.B2(n_631),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_737),
.B(n_326),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_618),
.B(n_548),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_598),
.A2(n_608),
.B(n_607),
.C(n_659),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_618),
.B(n_548),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_599),
.A2(n_618),
.B(n_656),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_655),
.B(n_701),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_618),
.B(n_548),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_599),
.A2(n_618),
.B(n_656),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_737),
.B(n_326),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_638),
.Y(n_916)
);

AO21x1_ASAP7_75t_L g917 ( 
.A1(n_889),
.A2(n_877),
.B(n_858),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_856),
.A2(n_884),
.B(n_874),
.Y(n_918)
);

OA21x2_ASAP7_75t_L g919 ( 
.A1(n_874),
.A2(n_838),
.B(n_766),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_865),
.B(n_900),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_760),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_861),
.A2(n_902),
.B(n_893),
.Y(n_922)
);

NOR2x1_ASAP7_75t_L g923 ( 
.A(n_881),
.B(n_831),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_751),
.B(n_757),
.Y(n_924)
);

AOI221xp5_ASAP7_75t_L g925 ( 
.A1(n_796),
.A2(n_826),
.B1(n_793),
.B2(n_807),
.C(n_880),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_900),
.B(n_768),
.Y(n_926)
);

BUFx4_ASAP7_75t_SL g927 ( 
.A(n_839),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_759),
.B(n_864),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_882),
.A2(n_909),
.B(n_906),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_875),
.A2(n_891),
.B(n_872),
.Y(n_930)
);

OAI21x1_ASAP7_75t_L g931 ( 
.A1(n_753),
.A2(n_892),
.B(n_867),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_814),
.B(n_866),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_873),
.B(n_879),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_770),
.A2(n_776),
.B(n_811),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_762),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_871),
.A2(n_878),
.B(n_876),
.Y(n_936)
);

AOI21x1_ASAP7_75t_L g937 ( 
.A1(n_779),
.A2(n_869),
.B(n_791),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_763),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_886),
.A2(n_894),
.B(n_890),
.Y(n_939)
);

NOR2x1_ASAP7_75t_SL g940 ( 
.A(n_778),
.B(n_903),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_778),
.Y(n_941)
);

AO21x2_ASAP7_75t_L g942 ( 
.A1(n_798),
.A2(n_790),
.B(n_841),
.Y(n_942)
);

BUFx4f_ASAP7_75t_L g943 ( 
.A(n_836),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_SL g944 ( 
.A(n_828),
.B(n_833),
.C(n_834),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_SL g945 ( 
.A1(n_855),
.A2(n_754),
.B(n_761),
.Y(n_945)
);

NAND2x1_ASAP7_75t_L g946 ( 
.A(n_903),
.B(n_750),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_912),
.B(n_836),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_812),
.B(n_808),
.Y(n_948)
);

INVx3_ASAP7_75t_SL g949 ( 
.A(n_802),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_895),
.B(n_905),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_799),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_870),
.A2(n_888),
.B(n_911),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_908),
.A2(n_910),
.B(n_913),
.Y(n_953)
);

AOI21xp33_ASAP7_75t_L g954 ( 
.A1(n_830),
.A2(n_754),
.B(n_824),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_817),
.B(n_783),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_767),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_774),
.B(n_794),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_896),
.A2(n_899),
.B(n_914),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_799),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_804),
.A2(n_813),
.B(n_810),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_860),
.B(n_862),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_814),
.B(n_868),
.Y(n_962)
);

AOI21xp33_ASAP7_75t_L g963 ( 
.A1(n_830),
.A2(n_844),
.B(n_758),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_782),
.A2(n_786),
.B(n_846),
.C(n_798),
.Y(n_964)
);

AO31x2_ASAP7_75t_L g965 ( 
.A1(n_829),
.A2(n_775),
.A3(n_835),
.B(n_822),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_823),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_901),
.B(n_904),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_756),
.A2(n_916),
.B1(n_788),
.B2(n_818),
.Y(n_968)
);

BUFx4_ASAP7_75t_SL g969 ( 
.A(n_781),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_816),
.A2(n_843),
.B(n_787),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_SL g971 ( 
.A1(n_857),
.A2(n_803),
.B(n_907),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_883),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_800),
.B(n_764),
.Y(n_973)
);

OAI21x1_ASAP7_75t_L g974 ( 
.A1(n_840),
.A2(n_849),
.B(n_847),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_897),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_852),
.A2(n_854),
.B(n_837),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_785),
.A2(n_789),
.B(n_819),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_820),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_863),
.B(n_792),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_771),
.A2(n_772),
.B(n_755),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_805),
.Y(n_981)
);

NOR3xp33_ASAP7_75t_L g982 ( 
.A(n_915),
.B(n_752),
.C(n_784),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_780),
.B(n_883),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_850),
.A2(n_853),
.B(n_851),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_780),
.B(n_809),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_806),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_821),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_897),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_863),
.B(n_859),
.Y(n_989)
);

OAI21xp33_ASAP7_75t_L g990 ( 
.A1(n_887),
.A2(n_848),
.B(n_845),
.Y(n_990)
);

OAI21x1_ASAP7_75t_SL g991 ( 
.A1(n_769),
.A2(n_797),
.B(n_795),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_809),
.B(n_898),
.Y(n_992)
);

OAI21x1_ASAP7_75t_SL g993 ( 
.A1(n_863),
.A2(n_777),
.B(n_773),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_825),
.B(n_827),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_777),
.A2(n_815),
.B(n_832),
.Y(n_995)
);

AOI21xp33_ASAP7_75t_L g996 ( 
.A1(n_912),
.A2(n_750),
.B(n_773),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_777),
.A2(n_863),
.B(n_912),
.Y(n_997)
);

INVx6_ASAP7_75t_L g998 ( 
.A(n_885),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_885),
.Y(n_999)
);

NAND3xp33_ASAP7_75t_SL g1000 ( 
.A(n_777),
.B(n_773),
.C(n_801),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_801),
.A2(n_856),
.B(n_884),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_842),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_842),
.A2(n_877),
.B(n_906),
.C(n_858),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_842),
.A2(n_893),
.B(n_882),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_856),
.A2(n_884),
.B(n_874),
.Y(n_1005)
);

AOI21x1_ASAP7_75t_L g1006 ( 
.A1(n_753),
.A2(n_779),
.B(n_766),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_856),
.A2(n_884),
.B(n_874),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_900),
.Y(n_1008)
);

AOI221xp5_ASAP7_75t_SL g1009 ( 
.A1(n_882),
.A2(n_893),
.B1(n_909),
.B2(n_889),
.C(n_902),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_778),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_858),
.A2(n_906),
.B(n_877),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_900),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_901),
.B(n_326),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_757),
.B(n_759),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_751),
.B(n_757),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_901),
.B(n_326),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_757),
.B(n_759),
.Y(n_1017)
);

NAND2x1p5_ASAP7_75t_L g1018 ( 
.A(n_778),
.B(n_903),
.Y(n_1018)
);

BUFx10_ASAP7_75t_L g1019 ( 
.A(n_752),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_757),
.B(n_759),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_856),
.A2(n_884),
.B(n_874),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_856),
.A2(n_884),
.B(n_874),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_861),
.A2(n_902),
.B(n_893),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_L g1024 ( 
.A1(n_753),
.A2(n_779),
.B(n_766),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_865),
.B(n_505),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_856),
.A2(n_884),
.B(n_874),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_882),
.A2(n_909),
.B(n_893),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_760),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_865),
.B(n_505),
.Y(n_1029)
);

OAI22x1_ASAP7_75t_L g1030 ( 
.A1(n_858),
.A2(n_330),
.B1(n_352),
.B2(n_326),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_858),
.B(n_877),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_861),
.A2(n_902),
.B(n_893),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_757),
.B(n_759),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_778),
.Y(n_1034)
);

NAND2xp33_ASAP7_75t_L g1035 ( 
.A(n_861),
.B(n_902),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_L g1036 ( 
.A1(n_882),
.A2(n_909),
.B(n_893),
.C(n_889),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_858),
.A2(n_877),
.B(n_906),
.C(n_902),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_856),
.A2(n_884),
.B(n_874),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_881),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_858),
.A2(n_877),
.B1(n_906),
.B2(n_759),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_861),
.A2(n_902),
.B(n_893),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_856),
.A2(n_884),
.B(n_874),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_823),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_858),
.A2(n_877),
.B1(n_906),
.B2(n_759),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_765),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_858),
.A2(n_877),
.B1(n_906),
.B2(n_759),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_L g1047 ( 
.A1(n_753),
.A2(n_779),
.B(n_766),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_757),
.B(n_759),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_SL g1049 ( 
.A1(n_858),
.A2(n_906),
.B(n_877),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_778),
.B(n_903),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_865),
.B(n_505),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_856),
.A2(n_884),
.B(n_874),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_760),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_883),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_881),
.B(n_619),
.Y(n_1055)
);

CKINVDCx11_ASAP7_75t_R g1056 ( 
.A(n_949),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_966),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_966),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_L g1059 ( 
.A(n_1037),
.B(n_1011),
.Y(n_1059)
);

OR2x6_ASAP7_75t_L g1060 ( 
.A(n_972),
.B(n_998),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_967),
.B(n_1013),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_1055),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1016),
.A2(n_1031),
.B1(n_1040),
.B2(n_1044),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_924),
.B(n_1015),
.Y(n_1064)
);

NOR2x1_ASAP7_75t_SL g1065 ( 
.A(n_1000),
.B(n_983),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_957),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_932),
.B(n_962),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_L g1068 ( 
.A(n_1040),
.B(n_1044),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_1014),
.B(n_1017),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_925),
.A2(n_1046),
.B(n_1003),
.C(n_945),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_SL g1071 ( 
.A1(n_1027),
.A2(n_929),
.B(n_930),
.C(n_1032),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1014),
.B(n_1017),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_978),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_972),
.B(n_947),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_1046),
.A2(n_917),
.B1(n_971),
.B2(n_1030),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_969),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_982),
.A2(n_1033),
.B1(n_1048),
.B2(n_1020),
.Y(n_1077)
);

OA21x2_ASAP7_75t_L g1078 ( 
.A1(n_930),
.A2(n_952),
.B(n_970),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_972),
.B(n_947),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_1036),
.A2(n_954),
.B(n_1048),
.C(n_1020),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_957),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_927),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_943),
.Y(n_1083)
);

OR2x6_ASAP7_75t_SL g1084 ( 
.A(n_994),
.B(n_973),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_943),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_961),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_L g1087 ( 
.A(n_1033),
.B(n_1027),
.Y(n_1087)
);

AND2x6_ASAP7_75t_L g1088 ( 
.A(n_979),
.B(n_975),
.Y(n_1088)
);

BUFx12f_ASAP7_75t_L g1089 ( 
.A(n_998),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_1054),
.B(n_997),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_961),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_997),
.B(n_959),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_959),
.B(n_975),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1023),
.A2(n_1041),
.B(n_1035),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_920),
.B(n_1025),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1029),
.B(n_1051),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_928),
.B(n_1008),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_1002),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_921),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1008),
.B(n_926),
.Y(n_1100)
);

OA21x2_ASAP7_75t_L g1101 ( 
.A1(n_952),
.A2(n_960),
.B(n_958),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_1039),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_988),
.B(n_951),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_928),
.B(n_981),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_954),
.A2(n_963),
.B(n_944),
.C(n_1009),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_1043),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_936),
.A2(n_953),
.B(n_939),
.Y(n_1107)
);

INVx6_ASAP7_75t_L g1108 ( 
.A(n_1019),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_963),
.A2(n_1009),
.B(n_964),
.C(n_950),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_950),
.A2(n_955),
.B(n_933),
.C(n_979),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_933),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_988),
.B(n_985),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_1012),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_935),
.Y(n_1114)
);

INVx5_ASAP7_75t_L g1115 ( 
.A(n_987),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_938),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_999),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_956),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1028),
.Y(n_1119)
);

AND2x6_ASAP7_75t_L g1120 ( 
.A(n_989),
.B(n_1010),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_946),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1019),
.B(n_1053),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_923),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_992),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1018),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_986),
.B(n_955),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1004),
.A2(n_948),
.B(n_968),
.C(n_977),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_989),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_990),
.B(n_995),
.Y(n_1129)
);

CKINVDCx20_ASAP7_75t_R g1130 ( 
.A(n_996),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_940),
.B(n_1034),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1018),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1045),
.B(n_968),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_991),
.A2(n_993),
.B1(n_996),
.B2(n_942),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1050),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_941),
.B(n_1034),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_941),
.A2(n_1010),
.B(n_919),
.C(n_942),
.Y(n_1137)
);

NOR2x1_ASAP7_75t_L g1138 ( 
.A(n_919),
.B(n_1050),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_976),
.B(n_984),
.Y(n_1139)
);

BUFx12f_ASAP7_75t_L g1140 ( 
.A(n_965),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_965),
.Y(n_1141)
);

OAI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_937),
.A2(n_1047),
.B1(n_1024),
.B2(n_1006),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_931),
.B(n_1001),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_918),
.B(n_1052),
.Y(n_1144)
);

AND2x2_ASAP7_75t_SL g1145 ( 
.A(n_974),
.B(n_1021),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_934),
.A2(n_1005),
.B(n_1007),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_L g1147 ( 
.A1(n_1022),
.A2(n_1026),
.B(n_1038),
.C(n_1042),
.Y(n_1147)
);

HAxp5_ASAP7_75t_L g1148 ( 
.A(n_967),
.B(n_648),
.CON(n_1148),
.SN(n_1148)
);

INVxp67_ASAP7_75t_SL g1149 ( 
.A(n_1012),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_972),
.B(n_912),
.Y(n_1150)
);

INVx5_ASAP7_75t_L g1151 ( 
.A(n_972),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_967),
.B(n_326),
.Y(n_1152)
);

BUFx2_ASAP7_75t_R g1153 ( 
.A(n_999),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_924),
.B(n_1015),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_SL g1155 ( 
.A1(n_1027),
.A2(n_929),
.B(n_930),
.C(n_922),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1037),
.A2(n_902),
.B(n_861),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_924),
.B(n_1015),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_924),
.B(n_1015),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_972),
.B(n_912),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_1055),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_972),
.B(n_912),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_932),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_957),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1037),
.A2(n_902),
.B(n_861),
.Y(n_1164)
);

CKINVDCx11_ASAP7_75t_R g1165 ( 
.A(n_949),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_924),
.B(n_1015),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_924),
.B(n_1015),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_924),
.B(n_1015),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1055),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1013),
.A2(n_629),
.B1(n_796),
.B2(n_505),
.Y(n_1170)
);

BUFx2_ASAP7_75t_L g1171 ( 
.A(n_1055),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_924),
.B(n_1015),
.Y(n_1172)
);

OR2x2_ASAP7_75t_SL g1173 ( 
.A(n_998),
.B(n_179),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1037),
.A2(n_902),
.B(n_861),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_SL g1175 ( 
.A1(n_1027),
.A2(n_929),
.B(n_930),
.C(n_922),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_967),
.B(n_326),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_957),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_924),
.B(n_1015),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1037),
.A2(n_793),
.B(n_882),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_932),
.B(n_962),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_978),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_969),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1037),
.A2(n_893),
.B(n_909),
.C(n_882),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_969),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_924),
.B(n_1015),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1055),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_957),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_967),
.A2(n_877),
.B1(n_906),
.B2(n_858),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1055),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_932),
.B(n_962),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_924),
.B(n_1015),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1037),
.A2(n_893),
.B(n_909),
.C(n_882),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_967),
.B(n_326),
.Y(n_1193)
);

INVxp67_ASAP7_75t_L g1194 ( 
.A(n_932),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_924),
.B(n_1015),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_926),
.B(n_973),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1013),
.A2(n_629),
.B1(n_796),
.B2(n_505),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1055),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_932),
.B(n_962),
.Y(n_1199)
);

INVx3_ASAP7_75t_SL g1200 ( 
.A(n_998),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1061),
.A2(n_1059),
.B1(n_1193),
.B2(n_1176),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1090),
.B(n_1092),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1073),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1152),
.A2(n_1068),
.B1(n_1164),
.B2(n_1156),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1070),
.B(n_1063),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1067),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1122),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1162),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1181),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1099),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1057),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1111),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1170),
.A2(n_1197),
.B1(n_1188),
.B2(n_1075),
.Y(n_1213)
);

BUFx8_ASAP7_75t_L g1214 ( 
.A(n_1089),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1077),
.A2(n_1179),
.B1(n_1174),
.B2(n_1192),
.Y(n_1215)
);

NAND2x1p5_ASAP7_75t_L g1216 ( 
.A(n_1151),
.B(n_1083),
.Y(n_1216)
);

BUFx10_ASAP7_75t_L g1217 ( 
.A(n_1076),
.Y(n_1217)
);

AO21x2_ASAP7_75t_L g1218 ( 
.A1(n_1107),
.A2(n_1142),
.B(n_1133),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1090),
.Y(n_1219)
);

NAND2x1p5_ASAP7_75t_L g1220 ( 
.A(n_1151),
.B(n_1083),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1151),
.B(n_1083),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1180),
.B(n_1190),
.Y(n_1222)
);

OAI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1084),
.A2(n_1172),
.B1(n_1168),
.B2(n_1154),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1114),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1116),
.Y(n_1225)
);

BUFx2_ASAP7_75t_R g1226 ( 
.A(n_1182),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1092),
.A2(n_1130),
.B1(n_1140),
.B2(n_1065),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1120),
.Y(n_1228)
);

AO21x2_ASAP7_75t_L g1229 ( 
.A1(n_1129),
.A2(n_1127),
.B(n_1110),
.Y(n_1229)
);

NAND2x1p5_ASAP7_75t_L g1230 ( 
.A(n_1085),
.B(n_1150),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1118),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1112),
.B(n_1093),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1147),
.A2(n_1101),
.B(n_1078),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1119),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1087),
.A2(n_1096),
.B1(n_1072),
.B2(n_1069),
.Y(n_1235)
);

CKINVDCx11_ASAP7_75t_R g1236 ( 
.A(n_1200),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1120),
.Y(n_1237)
);

NAND2x1p5_ASAP7_75t_L g1238 ( 
.A(n_1085),
.B(n_1150),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1097),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1125),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1199),
.A2(n_1095),
.B1(n_1185),
.B2(n_1158),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1137),
.B(n_1183),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1064),
.A2(n_1166),
.B1(n_1178),
.B2(n_1167),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1184),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1157),
.A2(n_1191),
.B1(n_1195),
.B2(n_1126),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1143),
.A2(n_1144),
.B(n_1138),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1066),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1081),
.A2(n_1091),
.B1(n_1086),
.B2(n_1177),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1102),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1105),
.A2(n_1141),
.B(n_1109),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1128),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1163),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1120),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1187),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1104),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1194),
.A2(n_1100),
.B1(n_1196),
.B2(n_1112),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1149),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1123),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1124),
.A2(n_1093),
.B1(n_1113),
.B2(n_1088),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1080),
.B(n_1134),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1088),
.A2(n_1103),
.B1(n_1079),
.B2(n_1074),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1101),
.A2(n_1132),
.B(n_1145),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1085),
.B(n_1108),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1103),
.Y(n_1264)
);

INVx5_ASAP7_75t_L g1265 ( 
.A(n_1088),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1088),
.B(n_1074),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1079),
.A2(n_1159),
.B1(n_1161),
.B2(n_1060),
.Y(n_1267)
);

OAI22x1_ASAP7_75t_L g1268 ( 
.A1(n_1139),
.A2(n_1155),
.B1(n_1175),
.B2(n_1071),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1098),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1060),
.A2(n_1117),
.B1(n_1108),
.B2(n_1062),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1136),
.B(n_1169),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1139),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1143),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1131),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1121),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1121),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1135),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1131),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1171),
.B(n_1186),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1121),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1160),
.A2(n_1198),
.B1(n_1189),
.B2(n_1115),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1056),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1173),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1115),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1115),
.A2(n_1058),
.B1(n_1106),
.B2(n_1148),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1082),
.B(n_1153),
.Y(n_1286)
);

BUFx2_ASAP7_75t_R g1287 ( 
.A(n_1165),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1077),
.B(n_1069),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1170),
.A2(n_629),
.B1(n_1197),
.B2(n_796),
.Y(n_1289)
);

AO21x1_ASAP7_75t_L g1290 ( 
.A1(n_1059),
.A2(n_1049),
.B(n_1031),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1152),
.A2(n_1193),
.B1(n_1176),
.B2(n_1061),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1061),
.B(n_1063),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1120),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1162),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1073),
.Y(n_1295)
);

AOI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1146),
.A2(n_937),
.B(n_1094),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1070),
.B(n_1063),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1073),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1061),
.A2(n_877),
.B1(n_906),
.B2(n_858),
.Y(n_1299)
);

INVxp67_ASAP7_75t_SL g1300 ( 
.A(n_1100),
.Y(n_1300)
);

AO21x2_ASAP7_75t_L g1301 ( 
.A1(n_1107),
.A2(n_980),
.B(n_1142),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1073),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1120),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1120),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1061),
.A2(n_334),
.B1(n_307),
.B2(n_322),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1067),
.B(n_1180),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1146),
.A2(n_937),
.B(n_1094),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1057),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1162),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1073),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1073),
.Y(n_1311)
);

BUFx12f_ASAP7_75t_L g1312 ( 
.A(n_1076),
.Y(n_1312)
);

INVx8_ASAP7_75t_L g1313 ( 
.A(n_1089),
.Y(n_1313)
);

BUFx2_ASAP7_75t_SL g1314 ( 
.A(n_1117),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1073),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1212),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1246),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1265),
.Y(n_1318)
);

BUFx8_ASAP7_75t_SL g1319 ( 
.A(n_1312),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1262),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1265),
.B(n_1228),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_1208),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1201),
.A2(n_1292),
.B(n_1299),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1262),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1219),
.B(n_1294),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1228),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1202),
.B(n_1205),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1309),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1247),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_1257),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1202),
.B(n_1205),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1252),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1314),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1297),
.B(n_1272),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1250),
.B(n_1210),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1292),
.A2(n_1291),
.B1(n_1204),
.B2(n_1213),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1250),
.B(n_1224),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_1250),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1215),
.A2(n_1213),
.B(n_1235),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_L g1340 ( 
.A(n_1254),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1249),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1265),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1288),
.B(n_1245),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_L g1344 ( 
.A(n_1223),
.B(n_1243),
.C(n_1260),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1225),
.Y(n_1345)
);

OAI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1260),
.A2(n_1242),
.B(n_1243),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1233),
.A2(n_1307),
.B(n_1296),
.Y(n_1347)
);

INVx5_ASAP7_75t_SL g1348 ( 
.A(n_1242),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1231),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1234),
.Y(n_1350)
);

INVxp33_ASAP7_75t_L g1351 ( 
.A(n_1263),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1218),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1242),
.Y(n_1353)
);

OR2x6_ASAP7_75t_L g1354 ( 
.A(n_1242),
.B(n_1273),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1218),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1237),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1229),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1207),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1229),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1222),
.B(n_1306),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1264),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1245),
.A2(n_1289),
.B(n_1285),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1301),
.B(n_1274),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1206),
.B(n_1300),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1203),
.Y(n_1365)
);

AOI21xp33_ASAP7_75t_L g1366 ( 
.A1(n_1290),
.A2(n_1289),
.B(n_1239),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1268),
.A2(n_1284),
.B(n_1277),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1209),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1274),
.B(n_1237),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1253),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1253),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1274),
.B(n_1253),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1312),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1293),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1295),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1303),
.B(n_1304),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1255),
.B(n_1241),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1298),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1302),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1275),
.A2(n_1280),
.B(n_1259),
.Y(n_1380)
);

OR2x6_ASAP7_75t_L g1381 ( 
.A(n_1266),
.B(n_1232),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1258),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1278),
.Y(n_1383)
);

OR2x6_ASAP7_75t_L g1384 ( 
.A(n_1266),
.B(n_1232),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1284),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1310),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_1282),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1311),
.A2(n_1315),
.B(n_1251),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1363),
.B(n_1268),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1363),
.B(n_1248),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1322),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1328),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1321),
.B(n_1232),
.Y(n_1393)
);

AND2x2_ASAP7_75t_SL g1394 ( 
.A(n_1353),
.B(n_1261),
.Y(n_1394)
);

INVxp33_ASAP7_75t_L g1395 ( 
.A(n_1358),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1330),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1340),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1335),
.B(n_1241),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1343),
.B(n_1256),
.Y(n_1399)
);

NAND2xp33_ASAP7_75t_SL g1400 ( 
.A(n_1336),
.B(n_1282),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1337),
.B(n_1271),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1357),
.B(n_1269),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1325),
.B(n_1279),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1355),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1382),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1320),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1320),
.B(n_1286),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1316),
.Y(n_1408)
);

OAI221xp5_ASAP7_75t_L g1409 ( 
.A1(n_1323),
.A2(n_1305),
.B1(n_1270),
.B2(n_1227),
.C(n_1283),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1324),
.B(n_1286),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1324),
.B(n_1286),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1334),
.B(n_1211),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1347),
.B(n_1308),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1325),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1352),
.A2(n_1281),
.B(n_1263),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1347),
.B(n_1276),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1339),
.A2(n_1221),
.B(n_1216),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1356),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1345),
.B(n_1349),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1349),
.B(n_1240),
.Y(n_1420)
);

INVx4_ASAP7_75t_L g1421 ( 
.A(n_1318),
.Y(n_1421)
);

OAI221xp5_ASAP7_75t_L g1422 ( 
.A1(n_1344),
.A2(n_1267),
.B1(n_1238),
.B2(n_1230),
.C(n_1220),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_R g1423 ( 
.A(n_1373),
.B(n_1236),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1396),
.B(n_1341),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1396),
.B(n_1361),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1397),
.B(n_1364),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1397),
.B(n_1364),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1391),
.B(n_1360),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1389),
.B(n_1327),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1409),
.A2(n_1344),
.B(n_1362),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1409),
.A2(n_1346),
.B1(n_1348),
.B2(n_1353),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1409),
.A2(n_1366),
.B1(n_1377),
.B2(n_1353),
.Y(n_1432)
);

OAI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1400),
.A2(n_1338),
.B1(n_1359),
.B2(n_1350),
.C(n_1329),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1389),
.B(n_1407),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1422),
.A2(n_1348),
.B1(n_1353),
.B2(n_1333),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1391),
.B(n_1360),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1400),
.B(n_1329),
.C(n_1332),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1399),
.A2(n_1388),
.B1(n_1354),
.B2(n_1378),
.Y(n_1438)
);

OAI21xp33_ASAP7_75t_L g1439 ( 
.A1(n_1390),
.A2(n_1332),
.B(n_1367),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1407),
.B(n_1331),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1419),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1417),
.B(n_1348),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1392),
.B(n_1401),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1392),
.B(n_1385),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_SL g1445 ( 
.A(n_1417),
.B(n_1348),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1401),
.B(n_1385),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1407),
.B(n_1356),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1406),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1401),
.B(n_1385),
.Y(n_1449)
);

NAND3xp33_ASAP7_75t_SL g1450 ( 
.A(n_1423),
.B(n_1387),
.C(n_1351),
.Y(n_1450)
);

NAND4xp25_ASAP7_75t_L g1451 ( 
.A(n_1405),
.B(n_1370),
.C(n_1374),
.D(n_1352),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_L g1452 ( 
.A(n_1405),
.B(n_1385),
.C(n_1386),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1401),
.B(n_1383),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_L g1454 ( 
.A(n_1402),
.B(n_1375),
.C(n_1386),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1417),
.A2(n_1422),
.B(n_1402),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1414),
.B(n_1419),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1410),
.B(n_1369),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1393),
.B(n_1371),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1399),
.A2(n_1390),
.B1(n_1394),
.B2(n_1422),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1411),
.B(n_1372),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1414),
.B(n_1383),
.Y(n_1461)
);

OAI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1390),
.A2(n_1367),
.B(n_1380),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1419),
.B(n_1326),
.Y(n_1463)
);

OAI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1402),
.A2(n_1317),
.B1(n_1368),
.B2(n_1379),
.C(n_1365),
.Y(n_1464)
);

OAI221xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1390),
.A2(n_1384),
.B1(n_1381),
.B2(n_1354),
.C(n_1376),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1441),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1441),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1434),
.B(n_1413),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1434),
.B(n_1413),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1448),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1454),
.B(n_1456),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1443),
.B(n_1403),
.Y(n_1472)
);

NAND2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1442),
.B(n_1342),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1448),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1426),
.B(n_1403),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1454),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1453),
.B(n_1419),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1452),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1452),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1429),
.B(n_1413),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1427),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1464),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1446),
.B(n_1413),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1449),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1445),
.B(n_1342),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1429),
.B(n_1416),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1425),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1461),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1424),
.B(n_1418),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1447),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1428),
.B(n_1395),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1463),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1455),
.B(n_1408),
.Y(n_1493)
);

INVx4_ASAP7_75t_L g1494 ( 
.A(n_1447),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_SL g1495 ( 
.A(n_1430),
.B(n_1421),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1440),
.B(n_1416),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1444),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1436),
.B(n_1418),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1451),
.B(n_1418),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1494),
.B(n_1437),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1482),
.B(n_1395),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1491),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1475),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1494),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1475),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1476),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1472),
.B(n_1451),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1482),
.B(n_1420),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1472),
.B(n_1412),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1491),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1476),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1494),
.B(n_1457),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1481),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1467),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1467),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1472),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1487),
.B(n_1420),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1493),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1498),
.B(n_1412),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1480),
.B(n_1460),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1493),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1480),
.B(n_1437),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1487),
.B(n_1420),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1471),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1471),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1488),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1478),
.B(n_1450),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1498),
.B(n_1412),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1488),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1468),
.B(n_1411),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1478),
.B(n_1430),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1466),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1479),
.B(n_1420),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1501),
.B(n_1313),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1531),
.B(n_1479),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1530),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1531),
.B(n_1492),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1518),
.B(n_1492),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1506),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1511),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1500),
.B(n_1458),
.Y(n_1541)
);

OAI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1527),
.A2(n_1495),
.B1(n_1433),
.B2(n_1431),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1527),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1526),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1529),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1521),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1522),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1503),
.B(n_1489),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1507),
.A2(n_1499),
.B1(n_1495),
.B2(n_1431),
.Y(n_1549)
);

A2O1A1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1500),
.A2(n_1439),
.B(n_1432),
.C(n_1522),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1512),
.Y(n_1551)
);

OAI22xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1524),
.A2(n_1499),
.B1(n_1465),
.B2(n_1462),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1502),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1525),
.B(n_1484),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1505),
.B(n_1489),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1510),
.B(n_1484),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1508),
.B(n_1287),
.Y(n_1557)
);

NOR2xp67_ASAP7_75t_L g1558 ( 
.A(n_1500),
.B(n_1499),
.Y(n_1558)
);

OAI21xp33_ASAP7_75t_L g1559 ( 
.A1(n_1522),
.A2(n_1497),
.B(n_1489),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1520),
.B(n_1490),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1520),
.B(n_1496),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1504),
.B(n_1236),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1516),
.B(n_1498),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1519),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1504),
.B(n_1319),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1533),
.B(n_1477),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1514),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1517),
.B(n_1483),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1523),
.B(n_1486),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1509),
.B(n_1477),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1528),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1504),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1543),
.A2(n_1439),
.B1(n_1459),
.B2(n_1394),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1539),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1543),
.A2(n_1535),
.B1(n_1550),
.B2(n_1542),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1541),
.B(n_1562),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1547),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1539),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1546),
.B(n_1515),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1552),
.A2(n_1394),
.B1(n_1462),
.B2(n_1398),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1542),
.A2(n_1394),
.B1(n_1398),
.B2(n_1415),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1568),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1548),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1540),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1553),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1555),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1561),
.B(n_1530),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1546),
.B(n_1537),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1544),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1573),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1564),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1536),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1545),
.Y(n_1594)
);

INVx1_ASAP7_75t_SL g1595 ( 
.A(n_1563),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1538),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1536),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1534),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1558),
.B(n_1530),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1554),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1556),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1551),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1560),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1579),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1586),
.B(n_1557),
.Y(n_1605)
);

AOI32xp33_ASAP7_75t_L g1606 ( 
.A1(n_1576),
.A2(n_1557),
.A3(n_1559),
.B1(n_1550),
.B2(n_1549),
.Y(n_1606)
);

OAI31xp33_ASAP7_75t_L g1607 ( 
.A1(n_1576),
.A2(n_1581),
.A3(n_1582),
.B(n_1574),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1581),
.A2(n_1534),
.B1(n_1415),
.B2(n_1394),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1579),
.Y(n_1609)
);

NAND2xp33_ASAP7_75t_L g1610 ( 
.A(n_1586),
.B(n_1423),
.Y(n_1610)
);

OAI311xp33_ASAP7_75t_L g1611 ( 
.A1(n_1582),
.A2(n_1567),
.A3(n_1570),
.B1(n_1569),
.C1(n_1571),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1596),
.B(n_1572),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1575),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1575),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1596),
.B(n_1572),
.Y(n_1615)
);

AOI21xp33_ASAP7_75t_L g1616 ( 
.A1(n_1578),
.A2(n_1563),
.B(n_1534),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1574),
.A2(n_1566),
.B1(n_1435),
.B2(n_1411),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1591),
.B(n_1565),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1583),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1583),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1588),
.B(n_1496),
.Y(n_1621)
);

OAI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1601),
.A2(n_1532),
.B1(n_1485),
.B2(n_1473),
.C(n_1438),
.Y(n_1622)
);

AOI21xp33_ASAP7_75t_L g1623 ( 
.A1(n_1578),
.A2(n_1415),
.B(n_1404),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1585),
.Y(n_1624)
);

OAI21xp33_ASAP7_75t_L g1625 ( 
.A1(n_1589),
.A2(n_1497),
.B(n_1474),
.Y(n_1625)
);

AOI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1578),
.A2(n_1470),
.B(n_1469),
.Y(n_1626)
);

INVx1_ASAP7_75t_SL g1627 ( 
.A(n_1591),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1589),
.A2(n_1474),
.B(n_1470),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1595),
.Y(n_1629)
);

NOR2x1_ASAP7_75t_L g1630 ( 
.A(n_1627),
.B(n_1597),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1629),
.B(n_1587),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1605),
.B(n_1588),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1604),
.Y(n_1633)
);

NOR2x1_ASAP7_75t_L g1634 ( 
.A(n_1610),
.B(n_1597),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1609),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1619),
.Y(n_1636)
);

NAND2xp33_ASAP7_75t_SL g1637 ( 
.A(n_1618),
.B(n_1599),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1610),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1626),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1605),
.B(n_1588),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1620),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1612),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1624),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1613),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1621),
.B(n_1598),
.Y(n_1645)
);

INVxp67_ASAP7_75t_SL g1646 ( 
.A(n_1615),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1616),
.B(n_1595),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1614),
.Y(n_1648)
);

NAND2xp33_ASAP7_75t_L g1649 ( 
.A(n_1606),
.B(n_1244),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1625),
.B(n_1577),
.Y(n_1650)
);

AOI32xp33_ASAP7_75t_L g1651 ( 
.A1(n_1649),
.A2(n_1611),
.A3(n_1608),
.B1(n_1584),
.B2(n_1587),
.Y(n_1651)
);

AND3x1_ASAP7_75t_L g1652 ( 
.A(n_1634),
.B(n_1607),
.C(n_1598),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1630),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1630),
.A2(n_1617),
.B(n_1608),
.C(n_1622),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1631),
.A2(n_1580),
.B(n_1598),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1638),
.A2(n_1587),
.B1(n_1592),
.B2(n_1584),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_SL g1657 ( 
.A(n_1637),
.B(n_1244),
.C(n_1628),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1632),
.B(n_1592),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1642),
.A2(n_1646),
.B1(n_1639),
.B2(n_1647),
.C(n_1644),
.Y(n_1659)
);

AO22x2_ASAP7_75t_SL g1660 ( 
.A1(n_1647),
.A2(n_1226),
.B1(n_1602),
.B2(n_1592),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1639),
.A2(n_1623),
.B1(n_1601),
.B2(n_1600),
.C(n_1584),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1652),
.B(n_1635),
.C(n_1633),
.Y(n_1662)
);

NOR2x1_ASAP7_75t_L g1663 ( 
.A(n_1658),
.B(n_1633),
.Y(n_1663)
);

NOR2x1_ASAP7_75t_L g1664 ( 
.A(n_1656),
.B(n_1635),
.Y(n_1664)
);

BUFx8_ASAP7_75t_SL g1665 ( 
.A(n_1660),
.Y(n_1665)
);

AOI211x1_ASAP7_75t_L g1666 ( 
.A1(n_1655),
.A2(n_1632),
.B(n_1640),
.C(n_1650),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1653),
.B(n_1640),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1657),
.B(n_1645),
.Y(n_1668)
);

NOR2x1_ASAP7_75t_L g1669 ( 
.A(n_1659),
.B(n_1644),
.Y(n_1669)
);

NAND3x1_ASAP7_75t_L g1670 ( 
.A(n_1661),
.B(n_1648),
.C(n_1643),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1669),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1666),
.B(n_1645),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1662),
.A2(n_1651),
.B(n_1641),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1663),
.Y(n_1674)
);

AND3x1_ASAP7_75t_L g1675 ( 
.A(n_1664),
.B(n_1641),
.C(n_1650),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1671),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1675),
.A2(n_1670),
.B1(n_1667),
.B2(n_1645),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1674),
.B(n_1636),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1672),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1673),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1671),
.Y(n_1681)
);

NOR2x1p5_ASAP7_75t_L g1682 ( 
.A(n_1676),
.B(n_1668),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1677),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1679),
.A2(n_1654),
.B1(n_1578),
.B2(n_1648),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1681),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1680),
.A2(n_1665),
.B1(n_1584),
.B2(n_1593),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1685),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1682),
.Y(n_1688)
);

NAND2x1p5_ASAP7_75t_L g1689 ( 
.A(n_1684),
.B(n_1678),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1687),
.Y(n_1690)
);

AND4x1_ASAP7_75t_L g1691 ( 
.A(n_1690),
.B(n_1686),
.C(n_1678),
.D(n_1687),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1691),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1691),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_SL g1694 ( 
.A1(n_1692),
.A2(n_1689),
.B(n_1688),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1693),
.B(n_1683),
.Y(n_1695)
);

OAI21x1_ASAP7_75t_L g1696 ( 
.A1(n_1695),
.A2(n_1643),
.B(n_1636),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1694),
.Y(n_1697)
);

AO21x2_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1593),
.B(n_1580),
.Y(n_1698)
);

AOI322xp5_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1696),
.A3(n_1593),
.B1(n_1600),
.B2(n_1603),
.C1(n_1597),
.C2(n_1594),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1594),
.B1(n_1590),
.B2(n_1585),
.C(n_1603),
.Y(n_1700)
);

AOI211xp5_ASAP7_75t_L g1701 ( 
.A1(n_1700),
.A2(n_1214),
.B(n_1217),
.C(n_1313),
.Y(n_1701)
);


endmodule