module fake_ariane_1246_n_106 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_106);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_106;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_81;
wire n_43;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_19),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVxp67_ASAP7_75t_SL g33 ( 
.A(n_3),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_R g39 ( 
.A(n_21),
.B(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_1),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OR2x6_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_28),
.Y(n_50)
);

OAI221xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_26),
.B1(n_30),
.B2(n_35),
.C(n_28),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_33),
.B1(n_34),
.B2(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

OAI221xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_35),
.B1(n_30),
.B2(n_26),
.C(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_56),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_54),
.B(n_29),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_47),
.B(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

OAI21x1_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_52),
.B(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_57),
.B1(n_47),
.B2(n_41),
.Y(n_66)
);

OA21x2_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_57),
.B(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_38),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_63),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_R g73 ( 
.A(n_69),
.B(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_71),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_76),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_75),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_88)
);

INVxp67_ASAP7_75t_SL g89 ( 
.A(n_83),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_4),
.Y(n_90)
);

AOI222xp33_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_43),
.B1(n_64),
.B2(n_85),
.C1(n_86),
.C2(n_72),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_90),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_87),
.B(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_73),
.A3(n_39),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_93),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_5),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_74),
.B(n_67),
.Y(n_99)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_94),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_100),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_98),
.Y(n_102)
);

OAI21x1_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_99),
.B(n_96),
.Y(n_103)
);

NAND5xp2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_6),
.C(n_8),
.D(n_67),
.E(n_64),
.Y(n_104)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_67),
.C(n_6),
.Y(n_105)
);

AO22x2_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_74),
.B1(n_10),
.B2(n_16),
.Y(n_106)
);


endmodule