module fake_netlist_6_2583_n_966 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_966);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_966;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_873;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_603;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_842;
wire n_720;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_624;
wire n_451;
wire n_824;
wire n_962;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_735;
wire n_483;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_386;
wire n_249;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_817;
wire n_701;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_262;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_949;
wire n_678;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_40),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_200),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_182),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_58),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_171),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_178),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_104),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_68),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_114),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_80),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_90),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_101),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_127),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_92),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g240 ( 
.A(n_132),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_149),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_55),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_91),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_157),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_108),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_105),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_147),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_174),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_95),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_172),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_117),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_204),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_209),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_144),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_137),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_151),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_23),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_94),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_141),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_179),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_199),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_201),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_67),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_153),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_121),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_183),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_152),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_111),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_73),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_11),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_62),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_37),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_155),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_72),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_116),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_41),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_110),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_85),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_112),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_202),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_168),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_74),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_170),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_142),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_186),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_206),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_129),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_113),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_164),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_102),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_97),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_225),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_134),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_109),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_49),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_140),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_221),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_219),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_10),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_100),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_222),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_78),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_9),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_133),
.Y(n_309)
);

HB1xp67_ASAP7_75t_SL g310 ( 
.A(n_184),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_130),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_1),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_223),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_135),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_32),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_197),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_47),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_193),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_99),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_47),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_124),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_32),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_181),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_175),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_180),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_208),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_131),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_42),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_162),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_148),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_88),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_191),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_20),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_195),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_54),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_145),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_158),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_138),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_82),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_163),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_12),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_55),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_119),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_79),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_122),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_118),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_22),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_70),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_34),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_81),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_48),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_212),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_70),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_98),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_120),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_30),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_125),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_63),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_14),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_139),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_8),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_187),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_103),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_59),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_128),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_3),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_73),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_37),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_26),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_59),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_45),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_74),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_28),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_51),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_25),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_31),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_75),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_77),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_10),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_16),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_75),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_36),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_161),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_136),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_194),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_166),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_29),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_67),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_169),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_123),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_203),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_205),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_160),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_377),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_259),
.B(n_0),
.Y(n_395)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_241),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_241),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_227),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_259),
.B(n_0),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_1),
.Y(n_401)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_241),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_239),
.B(n_2),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_241),
.Y(n_405)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_252),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_371),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_252),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_252),
.Y(n_410)
);

BUFx8_ASAP7_75t_L g411 ( 
.A(n_383),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_344),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_285),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_2),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_240),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_240),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_311),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_311),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_250),
.B(n_4),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_228),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_239),
.B(n_5),
.Y(n_421)
);

CKINVDCx6p67_ASAP7_75t_R g422 ( 
.A(n_275),
.Y(n_422)
);

BUFx8_ASAP7_75t_SL g423 ( 
.A(n_308),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_240),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_269),
.B(n_6),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_278),
.Y(n_426)
);

BUFx12f_ASAP7_75t_L g427 ( 
.A(n_344),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_231),
.Y(n_428)
);

INVx5_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_278),
.B(n_7),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_229),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_365),
.Y(n_432)
);

BUFx12f_ASAP7_75t_L g433 ( 
.A(n_226),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_282),
.B(n_7),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_327),
.B(n_8),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_282),
.B(n_11),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_269),
.B(n_13),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_289),
.B(n_13),
.Y(n_438)
);

INVx5_ASAP7_75t_L g439 ( 
.A(n_365),
.Y(n_439)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_365),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_365),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_294),
.B(n_14),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_240),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_289),
.B(n_15),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_294),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_313),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_313),
.B(n_15),
.Y(n_447)
);

AND2x4_ASAP7_75t_L g448 ( 
.A(n_316),
.B(n_17),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_367),
.B(n_17),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_374),
.B(n_18),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_316),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_321),
.B(n_18),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_233),
.B(n_19),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_320),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_321),
.B(n_21),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_240),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_332),
.B(n_21),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_355),
.B(n_23),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_245),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_341),
.B(n_347),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_391),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_24),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_232),
.B(n_234),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_281),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_237),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_304),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_328),
.B(n_26),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_333),
.B(n_342),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_366),
.B(n_27),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_235),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_359),
.B(n_27),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_361),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_261),
.B(n_29),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_356),
.B(n_31),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_369),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_372),
.B(n_33),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_380),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

INVx5_ASAP7_75t_L g479 ( 
.A(n_246),
.Y(n_479)
);

BUFx8_ASAP7_75t_L g480 ( 
.A(n_382),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_238),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_242),
.B(n_33),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_243),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_244),
.B(n_34),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_267),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_273),
.B(n_35),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_274),
.B(n_35),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_253),
.B(n_36),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_378),
.B(n_38),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_276),
.B(n_39),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_248),
.B(n_39),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_254),
.B(n_41),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_301),
.B(n_42),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_258),
.B(n_43),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_264),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_287),
.B(n_44),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_265),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_280),
.B(n_83),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_284),
.B(n_45),
.Y(n_499)
);

INVxp33_ASAP7_75t_SL g500 ( 
.A(n_300),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_310),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_291),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_295),
.B(n_46),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_307),
.B(n_46),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_309),
.B(n_50),
.Y(n_505)
);

NOR2x1p5_ASAP7_75t_L g506 ( 
.A(n_403),
.B(n_312),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_399),
.Y(n_507)
);

OAI22xp33_ASAP7_75t_L g508 ( 
.A1(n_490),
.A2(n_317),
.B1(n_322),
.B2(n_315),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_247),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_401),
.A2(n_236),
.B1(n_268),
.B2(n_230),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_SL g512 ( 
.A1(n_490),
.A2(n_348),
.B1(n_349),
.B2(n_335),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_414),
.A2(n_286),
.B1(n_288),
.B2(n_272),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_L g514 ( 
.A1(n_460),
.A2(n_353),
.B1(n_358),
.B2(n_351),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_412),
.B(n_364),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_398),
.B(n_318),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_404),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_L g519 ( 
.A1(n_460),
.A2(n_394),
.B1(n_488),
.B2(n_484),
.Y(n_519)
);

AO22x2_ASAP7_75t_L g520 ( 
.A1(n_395),
.A2(n_325),
.B1(n_326),
.B2(n_319),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_500),
.B(n_329),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_482),
.A2(n_493),
.B1(n_491),
.B2(n_433),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_397),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_397),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_496),
.A2(n_370),
.B1(n_373),
.B2(n_368),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_397),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_453),
.A2(n_386),
.B1(n_375),
.B2(n_376),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_485),
.B(n_249),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_485),
.B(n_251),
.Y(n_529)
);

CKINVDCx6p67_ASAP7_75t_R g530 ( 
.A(n_427),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_405),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_405),
.Y(n_532)
);

AND2x2_ASAP7_75t_SL g533 ( 
.A(n_469),
.B(n_330),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_473),
.A2(n_387),
.B1(n_388),
.B2(n_379),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_486),
.A2(n_256),
.B1(n_257),
.B2(n_255),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_487),
.A2(n_262),
.B1(n_263),
.B2(n_260),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_405),
.Y(n_537)
);

OAI22xp33_ASAP7_75t_L g538 ( 
.A1(n_484),
.A2(n_345),
.B1(n_346),
.B2(n_339),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_504),
.A2(n_270),
.B1(n_271),
.B2(n_266),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_420),
.B(n_277),
.Y(n_540)
);

AO22x2_ASAP7_75t_L g541 ( 
.A1(n_400),
.A2(n_392),
.B1(n_52),
.B2(n_50),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_409),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_409),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_409),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_413),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_435),
.A2(n_283),
.B1(n_290),
.B2(n_279),
.Y(n_546)
);

OAI22xp33_ASAP7_75t_L g547 ( 
.A1(n_488),
.A2(n_293),
.B1(n_296),
.B2(n_292),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_428),
.B(n_297),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_400),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_549)
);

OAI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_419),
.A2(n_299),
.B1(n_302),
.B2(n_298),
.Y(n_550)
);

AO22x2_ASAP7_75t_L g551 ( 
.A1(n_436),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_449),
.A2(n_393),
.B1(n_389),
.B2(n_385),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_470),
.B(n_384),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_413),
.Y(n_555)
);

AO22x2_ASAP7_75t_L g556 ( 
.A1(n_436),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_450),
.A2(n_362),
.B1(n_360),
.B2(n_357),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_417),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_417),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_492),
.A2(n_421),
.B1(n_425),
.B2(n_403),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_421),
.A2(n_354),
.B1(n_352),
.B2(n_350),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_417),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_408),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_494),
.A2(n_324),
.B1(n_340),
.B2(n_338),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_418),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_503),
.A2(n_343),
.B1(n_337),
.B2(n_336),
.Y(n_567)
);

INVx8_ASAP7_75t_L g568 ( 
.A(n_423),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_442),
.B(n_303),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_470),
.B(n_305),
.Y(n_570)
);

AO22x2_ASAP7_75t_L g571 ( 
.A1(n_442),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_426),
.B(n_306),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_505),
.A2(n_323),
.B1(n_334),
.B2(n_331),
.Y(n_573)
);

AND2x2_ASAP7_75t_SL g574 ( 
.A(n_434),
.B(n_447),
.Y(n_574)
);

OAI22xp33_ASAP7_75t_L g575 ( 
.A1(n_467),
.A2(n_314),
.B1(n_63),
.B2(n_64),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_422),
.B(n_84),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_445),
.B(n_86),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_445),
.B(n_463),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_447),
.B(n_87),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_R g580 ( 
.A1(n_474),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_578),
.B(n_463),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_560),
.A2(n_574),
.B(n_533),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_579),
.Y(n_583)
);

CKINVDCx14_ASAP7_75t_R g584 ( 
.A(n_530),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_524),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_526),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_526),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_537),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_528),
.A2(n_498),
.B(n_444),
.Y(n_589)
);

XOR2x2_ASAP7_75t_L g590 ( 
.A(n_512),
.B(n_489),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_507),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_523),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_572),
.B(n_430),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_531),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_532),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_542),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_543),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_507),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_544),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_545),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_529),
.B(n_396),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_555),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_579),
.B(n_448),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_562),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_563),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_566),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_516),
.B(n_497),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_559),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_579),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_511),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_540),
.B(n_548),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_521),
.B(n_502),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_517),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_517),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_518),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_518),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_553),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_579),
.B(n_448),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_467),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_553),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_570),
.B(n_464),
.Y(n_622)
);

AOI21x1_ASAP7_75t_L g623 ( 
.A1(n_577),
.A2(n_416),
.B(n_415),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_564),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_569),
.B(n_452),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_568),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_569),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_514),
.B(n_438),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_508),
.B(n_455),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_510),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_513),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_509),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_547),
.B(n_465),
.Y(n_633)
);

INVxp33_ASAP7_75t_L g634 ( 
.A(n_527),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_520),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_576),
.B(n_411),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_554),
.Y(n_637)
);

XNOR2x2_ASAP7_75t_L g638 ( 
.A(n_549),
.B(n_471),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g639 ( 
.A(n_506),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_541),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_546),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_515),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_549),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_534),
.B(n_565),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_551),
.Y(n_645)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_522),
.B(n_519),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_567),
.B(n_464),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_551),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_593),
.B(n_573),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_613),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_629),
.A2(n_538),
.B1(n_580),
.B2(n_571),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_591),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_625),
.B(n_556),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_591),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_632),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_608),
.B(n_561),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_608),
.B(n_552),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_637),
.B(n_622),
.Y(n_658)
);

AND2x6_ASAP7_75t_L g659 ( 
.A(n_603),
.B(n_452),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_625),
.B(n_556),
.Y(n_660)
);

AND2x2_ASAP7_75t_SL g661 ( 
.A(n_628),
.B(n_462),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_589),
.A2(n_557),
.B(n_536),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_614),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_628),
.A2(n_539),
.B(n_535),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_603),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_625),
.B(n_571),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_614),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_632),
.Y(n_668)
);

AND2x2_ASAP7_75t_SL g669 ( 
.A(n_603),
.B(n_619),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_615),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_637),
.B(n_498),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_619),
.B(n_498),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_610),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_581),
.B(n_462),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_598),
.B(n_477),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_619),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_598),
.B(n_477),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_626),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_582),
.B(n_478),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_610),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_632),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_634),
.B(n_550),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_615),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_647),
.B(n_478),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_616),
.Y(n_685)
);

AND2x2_ASAP7_75t_SL g686 ( 
.A(n_644),
.B(n_471),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_612),
.B(n_459),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_627),
.B(n_466),
.Y(n_688)
);

AND2x2_ASAP7_75t_SL g689 ( 
.A(n_610),
.B(n_476),
.Y(n_689)
);

INVx4_ASAP7_75t_L g690 ( 
.A(n_583),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_616),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_639),
.B(n_472),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_583),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_617),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_633),
.B(n_472),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_635),
.B(n_475),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_634),
.B(n_525),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_640),
.B(n_475),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_618),
.Y(n_699)
);

AND2x2_ASAP7_75t_SL g700 ( 
.A(n_640),
.B(n_476),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_623),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_621),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_642),
.Y(n_703)
);

OAI21xp5_ASAP7_75t_L g704 ( 
.A1(n_601),
.A2(n_499),
.B(n_457),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_624),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_611),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_592),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_594),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_595),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_642),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_643),
.B(n_431),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_641),
.B(n_575),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_596),
.B(n_446),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_597),
.B(n_599),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_645),
.B(n_431),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_642),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_600),
.Y(n_717)
);

OAI21xp5_ASAP7_75t_L g718 ( 
.A1(n_646),
.A2(n_458),
.B(n_437),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_602),
.B(n_446),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_604),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_648),
.B(n_605),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_SL g722 ( 
.A(n_661),
.B(n_641),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_665),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_703),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_695),
.B(n_606),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_654),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_652),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_703),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_663),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_678),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_SL g731 ( 
.A(n_664),
.B(n_636),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_665),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_695),
.B(n_607),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_703),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_650),
.B(n_630),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_679),
.B(n_658),
.Y(n_736)
);

NAND2x1p5_ASAP7_75t_L g737 ( 
.A(n_669),
.B(n_585),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_692),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_652),
.Y(n_739)
);

NAND2x1p5_ASAP7_75t_L g740 ( 
.A(n_669),
.B(n_586),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_657),
.B(n_631),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_663),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_692),
.Y(n_743)
);

INVx5_ASAP7_75t_L g744 ( 
.A(n_710),
.Y(n_744)
);

NAND2x1p5_ASAP7_75t_L g745 ( 
.A(n_676),
.B(n_655),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_667),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_675),
.B(n_587),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_SL g748 ( 
.A(n_662),
.B(n_631),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_667),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_716),
.Y(n_750)
);

NOR2x1_ASAP7_75t_L g751 ( 
.A(n_690),
.B(n_620),
.Y(n_751)
);

NAND2x1p5_ASAP7_75t_L g752 ( 
.A(n_676),
.B(n_655),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_668),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_687),
.B(n_584),
.Y(n_754)
);

NAND2x1p5_ASAP7_75t_L g755 ( 
.A(n_668),
.B(n_609),
.Y(n_755)
);

BUFx12f_ASAP7_75t_L g756 ( 
.A(n_696),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_681),
.Y(n_757)
);

AND2x2_ASAP7_75t_SL g758 ( 
.A(n_712),
.B(n_638),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_681),
.B(n_588),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_677),
.B(n_446),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_687),
.B(n_584),
.Y(n_761)
);

AND2x6_ASAP7_75t_L g762 ( 
.A(n_672),
.B(n_638),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_670),
.Y(n_763)
);

NAND2x1p5_ASAP7_75t_L g764 ( 
.A(n_690),
.B(n_454),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_686),
.B(n_649),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_656),
.B(n_700),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_672),
.B(n_424),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_696),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_685),
.Y(n_769)
);

BUFx4f_ASAP7_75t_L g770 ( 
.A(n_700),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_686),
.B(n_451),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_693),
.B(n_689),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_683),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_691),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_691),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_693),
.B(n_451),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_672),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_773),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_774),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_775),
.Y(n_780)
);

BUFx2_ASAP7_75t_SL g781 ( 
.A(n_744),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_728),
.Y(n_782)
);

BUFx2_ASAP7_75t_SL g783 ( 
.A(n_744),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_777),
.Y(n_784)
);

INVx8_ASAP7_75t_L g785 ( 
.A(n_767),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_727),
.Y(n_786)
);

INVx3_ASAP7_75t_SL g787 ( 
.A(n_730),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_726),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_766),
.B(n_736),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_735),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_729),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_753),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_742),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_777),
.B(n_768),
.Y(n_794)
);

INVx5_ASAP7_75t_L g795 ( 
.A(n_767),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_739),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_738),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_756),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_746),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_753),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_757),
.Y(n_801)
);

CKINVDCx6p67_ASAP7_75t_R g802 ( 
.A(n_754),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_749),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_757),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_762),
.Y(n_805)
);

INVx5_ASAP7_75t_SL g806 ( 
.A(n_728),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_723),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_723),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_763),
.Y(n_809)
);

INVx8_ASAP7_75t_L g810 ( 
.A(n_767),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_766),
.B(n_684),
.Y(n_811)
);

CKINVDCx6p67_ASAP7_75t_R g812 ( 
.A(n_761),
.Y(n_812)
);

INVx5_ASAP7_75t_L g813 ( 
.A(n_767),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_769),
.Y(n_814)
);

NAND2x1p5_ASAP7_75t_L g815 ( 
.A(n_724),
.B(n_673),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_762),
.Y(n_816)
);

BUFx12f_ASAP7_75t_L g817 ( 
.A(n_743),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_770),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_736),
.B(n_674),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_765),
.B(n_674),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_734),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_732),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_751),
.B(n_694),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_782),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_803),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_811),
.A2(n_748),
.B1(n_741),
.B2(n_758),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_814),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_SL g828 ( 
.A1(n_790),
.A2(n_651),
.B(n_697),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_787),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_811),
.A2(n_748),
.B1(n_731),
.B2(n_722),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_789),
.B(n_760),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_820),
.A2(n_731),
.B1(n_722),
.B2(n_718),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_819),
.A2(n_651),
.B(n_682),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_786),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_796),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_799),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_809),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_817),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_805),
.A2(n_733),
.B1(n_725),
.B2(n_772),
.Y(n_839)
);

BUFx10_ASAP7_75t_L g840 ( 
.A(n_797),
.Y(n_840)
);

INVx6_ASAP7_75t_L g841 ( 
.A(n_798),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_802),
.A2(n_590),
.B1(n_688),
.B2(n_771),
.Y(n_842)
);

BUFx10_ASAP7_75t_L g843 ( 
.A(n_823),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_816),
.A2(n_812),
.B1(n_802),
.B2(n_818),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_778),
.B(n_725),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_779),
.A2(n_733),
.B1(n_772),
.B2(n_747),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_812),
.A2(n_660),
.B1(n_666),
.B2(n_653),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_780),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_788),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_780),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_801),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_823),
.A2(n_659),
.B1(n_704),
.B2(n_696),
.Y(n_852)
);

BUFx10_ASAP7_75t_L g853 ( 
.A(n_823),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_791),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_833),
.A2(n_826),
.B1(n_832),
.B2(n_830),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_842),
.A2(n_740),
.B1(n_737),
.B2(n_795),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_839),
.A2(n_699),
.B1(n_705),
.B2(n_702),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_839),
.A2(n_699),
.B1(n_702),
.B2(n_694),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_844),
.A2(n_795),
.B1(n_813),
.B2(n_794),
.Y(n_859)
);

AOI211xp5_ASAP7_75t_L g860 ( 
.A1(n_828),
.A2(n_468),
.B(n_715),
.C(n_711),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_828),
.B(n_698),
.Y(n_861)
);

INVx5_ASAP7_75t_L g862 ( 
.A(n_824),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_825),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_846),
.A2(n_671),
.B(n_706),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_831),
.A2(n_709),
.B1(n_707),
.B2(n_480),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_845),
.A2(n_813),
.B1(n_745),
.B2(n_752),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_848),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_831),
.A2(n_717),
.B1(n_720),
.B2(n_708),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_834),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_835),
.A2(n_717),
.B1(n_720),
.B2(n_708),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_847),
.B(n_721),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_SL g872 ( 
.A1(n_852),
.A2(n_764),
.B(n_759),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_836),
.A2(n_791),
.B1(n_793),
.B2(n_714),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_837),
.A2(n_793),
.B1(n_481),
.B2(n_483),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_827),
.B(n_801),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_829),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_841),
.A2(n_810),
.B1(n_785),
.B2(n_783),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_850),
.Y(n_878)
);

INVx4_ASAP7_75t_SL g879 ( 
.A(n_824),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_SL g880 ( 
.A1(n_838),
.A2(n_804),
.B1(n_792),
.B2(n_800),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_849),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_854),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_851),
.B(n_792),
.Y(n_883)
);

OA21x2_ASAP7_75t_L g884 ( 
.A1(n_864),
.A2(n_776),
.B(n_719),
.Y(n_884)
);

OAI222xp33_ASAP7_75t_L g885 ( 
.A1(n_855),
.A2(n_822),
.B1(n_755),
.B2(n_851),
.C1(n_807),
.C2(n_808),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_SL g886 ( 
.A1(n_861),
.A2(n_856),
.B1(n_871),
.B2(n_880),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_860),
.B(n_713),
.C(n_495),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_875),
.B(n_843),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_865),
.A2(n_853),
.B1(n_840),
.B2(n_784),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_SL g890 ( 
.A1(n_859),
.A2(n_810),
.B1(n_785),
.B2(n_783),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_857),
.A2(n_806),
.B1(n_781),
.B2(n_750),
.Y(n_891)
);

OAI21xp33_ASAP7_75t_SL g892 ( 
.A1(n_858),
.A2(n_821),
.B(n_776),
.Y(n_892)
);

NOR3xp33_ASAP7_75t_L g893 ( 
.A(n_872),
.B(n_701),
.C(n_443),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_873),
.B(n_461),
.C(n_479),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_876),
.B(n_89),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_874),
.A2(n_815),
.B1(n_680),
.B2(n_461),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_874),
.A2(n_815),
.B1(n_680),
.B2(n_402),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_866),
.A2(n_867),
.B1(n_869),
.B2(n_870),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_867),
.A2(n_456),
.B1(n_479),
.B2(n_441),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_868),
.A2(n_402),
.B1(n_406),
.B2(n_440),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_870),
.A2(n_406),
.B1(n_440),
.B2(n_439),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_881),
.A2(n_882),
.B1(n_878),
.B2(n_863),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_877),
.A2(n_410),
.B1(n_439),
.B2(n_432),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_SL g904 ( 
.A1(n_883),
.A2(n_66),
.B(n_69),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_862),
.A2(n_69),
.B1(n_71),
.B2(n_76),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_902),
.B(n_879),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_SL g907 ( 
.A1(n_904),
.A2(n_905),
.B(n_886),
.Y(n_907)
);

NAND3xp33_ASAP7_75t_L g908 ( 
.A(n_887),
.B(n_432),
.C(n_429),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_898),
.B(n_93),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_884),
.B(n_96),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_888),
.B(n_106),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_893),
.B(n_107),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_889),
.B(n_115),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_892),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_895),
.B(n_126),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_890),
.B(n_410),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_891),
.B(n_143),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_885),
.A2(n_146),
.B(n_150),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_SL g919 ( 
.A1(n_894),
.A2(n_154),
.B1(n_156),
.B2(n_159),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_914),
.Y(n_920)
);

AND2x6_ASAP7_75t_L g921 ( 
.A(n_912),
.B(n_903),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_911),
.B(n_910),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_910),
.B(n_899),
.Y(n_923)
);

OR2x2_ASAP7_75t_L g924 ( 
.A(n_906),
.B(n_900),
.Y(n_924)
);

AO21x2_ASAP7_75t_L g925 ( 
.A1(n_916),
.A2(n_897),
.B(n_896),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_918),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_918),
.B(n_901),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_907),
.A2(n_165),
.B(n_167),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_918),
.B(n_173),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_L g930 ( 
.A(n_909),
.B(n_176),
.C(n_177),
.Y(n_930)
);

NAND4xp75_ASAP7_75t_L g931 ( 
.A(n_928),
.B(n_917),
.C(n_913),
.D(n_915),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_920),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_926),
.B(n_917),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_926),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_922),
.B(n_919),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_923),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_927),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_927),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_929),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_924),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_921),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_925),
.B(n_908),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_941),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_934),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_937),
.Y(n_945)
);

XNOR2xp5_ASAP7_75t_L g946 ( 
.A(n_931),
.B(n_930),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_933),
.Y(n_947)
);

AOI22x1_ASAP7_75t_L g948 ( 
.A1(n_946),
.A2(n_942),
.B1(n_939),
.B2(n_935),
.Y(n_948)
);

AO22x2_ASAP7_75t_L g949 ( 
.A1(n_943),
.A2(n_938),
.B1(n_936),
.B2(n_940),
.Y(n_949)
);

AO22x2_ASAP7_75t_L g950 ( 
.A1(n_947),
.A2(n_938),
.B1(n_937),
.B2(n_932),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_945),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_951),
.Y(n_952)
);

AOI22x1_ASAP7_75t_L g953 ( 
.A1(n_952),
.A2(n_949),
.B1(n_950),
.B2(n_948),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_953),
.Y(n_954)
);

NOR2x1_ASAP7_75t_L g955 ( 
.A(n_954),
.B(n_944),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_955),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_956),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_957),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_958),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_959),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_960),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_961),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_962),
.A2(n_192),
.B1(n_196),
.B2(n_198),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_963),
.Y(n_964)
);

AOI221xp5_ASAP7_75t_L g965 ( 
.A1(n_964),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.C(n_214),
.Y(n_965)
);

AOI211xp5_ASAP7_75t_L g966 ( 
.A1(n_965),
.A2(n_216),
.B(n_217),
.C(n_218),
.Y(n_966)
);


endmodule