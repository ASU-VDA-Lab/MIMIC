module real_jpeg_29755_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_0),
.B(n_58),
.Y(n_57)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_1),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_1),
.A2(n_29),
.B(n_33),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_1),
.B(n_31),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_1),
.A2(n_47),
.B(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_1),
.B(n_47),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_1),
.B(n_53),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_1),
.A2(n_56),
.B1(n_66),
.B2(n_226),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_1),
.A2(n_32),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_2),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_185)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_4),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_4),
.A2(n_25),
.B1(n_58),
.B2(n_59),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_4),
.A2(n_25),
.B1(n_47),
.B2(n_48),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_68),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_8),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_77),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_9),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_10),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_136),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_136),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_136),
.Y(n_226)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_11),
.A2(n_47),
.A3(n_59),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_12),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_99),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_99),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_99),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_13),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_13),
.A2(n_37),
.B1(n_58),
.B2(n_59),
.Y(n_215)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_15),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_46)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_16),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_16),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_63),
.Y(n_84)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_17),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_127),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_102),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_21),
.B(n_102),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_78),
.C(n_89),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_22),
.B(n_78),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_22),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_38),
.CI(n_54),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_23),
.B(n_38),
.C(n_54),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_24),
.A2(n_28),
.B1(n_31),
.B2(n_98),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_26),
.A2(n_35),
.B(n_140),
.C(n_141),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_28),
.A2(n_31),
.B1(n_135),
.B2(n_165),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_31),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_43),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g250 ( 
.A1(n_32),
.A2(n_43),
.A3(n_48),
.B1(n_243),
.B2(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_33),
.B(n_140),
.Y(n_243)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_36),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_51),
.B2(n_53),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_39),
.A2(n_41),
.B1(n_53),
.B2(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_41),
.A2(n_53),
.B1(n_163),
.B2(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_46),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_42),
.A2(n_46),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_42),
.A2(n_46),
.B1(n_146),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_42),
.A2(n_46),
.B1(n_183),
.B2(n_241),
.Y(n_240)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_43),
.Y(n_252)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_48),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_47),
.B(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_51),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_69),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_55),
.B(n_69),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B1(n_64),
.B2(n_67),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_67),
.B(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_56),
.A2(n_62),
.B1(n_64),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_56),
.A2(n_88),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_56),
.A2(n_88),
.B1(n_220),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_56),
.A2(n_64),
.B1(n_215),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_57),
.A2(n_93),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_57),
.A2(n_65),
.B1(n_143),
.B2(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_57),
.A2(n_65),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_59),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_58),
.B(n_74),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_58),
.B(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g88 ( 
.A(n_65),
.Y(n_88)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_76),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_72),
.B1(n_84),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_71),
.A2(n_72),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_71),
.A2(n_72),
.B1(n_201),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_71),
.A2(n_72),
.B1(n_168),
.B2(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_72),
.B(n_140),
.Y(n_227)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_76),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_86),
.B2(n_87),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_87),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_82),
.A2(n_85),
.B1(n_96),
.B2(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_82),
.A2(n_85),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_87),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_89),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_97),
.C(n_100),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_90),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_91),
.B(n_94),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_98),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_101),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_123),
.B2(n_124),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_112),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_111),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_109),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_119),
.B1(n_134),
.B2(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_123),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_151),
.B(n_278),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_149),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_129),
.B(n_149),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_148),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_148),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.C(n_145),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_145),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_142),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_140),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_188),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_171),
.B(n_187),
.Y(n_153)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_169),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_169),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_159),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.C(n_166),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_161),
.B1(n_166),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_174),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_175),
.B(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_276),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_178),
.Y(n_276)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.C(n_186),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_181),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_184),
.B(n_186),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_185),
.Y(n_254)
);

NOR3xp33_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.C(n_191),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_272),
.B(n_277),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_258),
.B(n_271),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_236),
.B(n_257),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_216),
.B(n_235),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_196),
.B(n_206),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_202),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_197),
.A2(n_198),
.B1(n_202),
.B2(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_212),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_214),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_223),
.B(n_234),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_222),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_228),
.B(n_233),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_227),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_237),
.B(n_238),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_249),
.B1(n_255),
.B2(n_256),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_244),
.B1(n_247),
.B2(n_248),
.Y(n_239)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_244),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_248),
.C(n_256),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_246),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_249),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_253),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_260),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_267),
.C(n_269),
.Y(n_273)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);


endmodule