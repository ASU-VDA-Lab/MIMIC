module fake_jpeg_8628_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_5),
.B(n_2),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_6),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_13),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_19),
.C(n_15),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_27),
.C(n_24),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_19),
.C(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_25),
.B(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_28),
.B(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_31),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_34),
.B(n_22),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_21),
.C(n_16),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_13),
.B(n_11),
.Y(n_35)
);

AOI322xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_36),
.A3(n_7),
.B1(n_34),
.B2(n_12),
.C1(n_9),
.C2(n_10),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_10),
.C(n_8),
.Y(n_38)
);


endmodule