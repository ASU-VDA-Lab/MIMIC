module fake_jpeg_3211_n_503 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_434;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_51),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_52),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx12f_ASAP7_75t_SL g59 ( 
.A(n_28),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_7),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_94),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_65),
.Y(n_146)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_80),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_86),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_15),
.B(n_14),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_87),
.B(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_15),
.B(n_7),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_20),
.B(n_6),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_13),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_9),
.Y(n_109)
);

BUFx24_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_99),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_109),
.B(n_137),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_56),
.A2(n_44),
.B1(n_42),
.B2(n_30),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_112),
.A2(n_113),
.B1(n_154),
.B2(n_38),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_46),
.B1(n_47),
.B2(n_45),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_18),
.B1(n_40),
.B2(n_28),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_149),
.B1(n_82),
.B2(n_68),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_64),
.A2(n_46),
.B1(n_31),
.B2(n_28),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_46),
.B1(n_31),
.B2(n_40),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_58),
.B(n_20),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_55),
.B(n_44),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_53),
.B(n_43),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_98),
.A2(n_28),
.B1(n_40),
.B2(n_42),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_71),
.B(n_30),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_40),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_81),
.A2(n_46),
.B1(n_45),
.B2(n_41),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_79),
.B(n_31),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_69),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_103),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_166),
.Y(n_212)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_175),
.Y(n_208)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_164),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_103),
.A2(n_41),
.B(n_86),
.C(n_96),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_165),
.A2(n_192),
.B(n_195),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_67),
.C(n_73),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_167),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_109),
.B(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_173),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_83),
.B1(n_70),
.B2(n_51),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_172),
.A2(n_180),
.B1(n_205),
.B2(n_159),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_106),
.B(n_19),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_106),
.A2(n_43),
.B1(n_19),
.B2(n_74),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_174),
.A2(n_181),
.B1(n_188),
.B2(n_189),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_65),
.B1(n_50),
.B2(n_52),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_176),
.A2(n_145),
.B1(n_151),
.B2(n_131),
.Y(n_225)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_177),
.Y(n_233)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_178),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_184),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_110),
.A2(n_40),
.B1(n_84),
.B2(n_55),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_182),
.B(n_183),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_129),
.B(n_100),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_123),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_185),
.B(n_186),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_114),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_104),
.B(n_99),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_136),
.A2(n_38),
.B1(n_39),
.B2(n_8),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_139),
.A2(n_38),
.B1(n_39),
.B2(n_8),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_193),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_38),
.B(n_39),
.C(n_8),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_0),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_123),
.B(n_9),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_116),
.Y(n_196)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_130),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_198),
.Y(n_214)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_201),
.Y(n_215)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_115),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_118),
.Y(n_204)
);

INVx11_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_167),
.A2(n_160),
.B1(n_111),
.B2(n_125),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_221),
.B1(n_232),
.B2(n_185),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_163),
.A2(n_159),
.B1(n_134),
.B2(n_142),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_225),
.B1(n_198),
.B2(n_192),
.Y(n_255)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_180),
.B1(n_178),
.B2(n_183),
.Y(n_232)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_231),
.A2(n_175),
.B(n_182),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_243),
.A2(n_214),
.B(n_207),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_173),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_245),
.C(n_253),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_171),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_209),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_246),
.B(n_248),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_193),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_247),
.B(n_251),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_254),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_233),
.Y(n_250)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_169),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_166),
.C(n_184),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_238),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_255),
.A2(n_239),
.B1(n_220),
.B2(n_213),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_161),
.C(n_165),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_263),
.C(n_213),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_215),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_257),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_241),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_258),
.B(n_260),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_187),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_169),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_241),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_265),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_219),
.B(n_187),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_195),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_268),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_215),
.B(n_186),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_231),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_266),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_226),
.A2(n_121),
.B(n_196),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_269),
.B(n_218),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_162),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_211),
.A2(n_203),
.B(n_199),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_194),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_237),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_177),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_232),
.A2(n_200),
.B1(n_197),
.B2(n_142),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_214),
.B1(n_233),
.B2(n_223),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_273),
.A2(n_279),
.B(n_285),
.Y(n_307)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_274),
.Y(n_306)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

OAI32xp33_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_260),
.A3(n_257),
.B1(n_270),
.B2(n_247),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_278),
.B(n_298),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_226),
.B(n_219),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_224),
.B1(n_207),
.B2(n_217),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_292),
.B1(n_301),
.B2(n_272),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_284),
.B(n_283),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_207),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_289),
.A2(n_294),
.B1(n_303),
.B2(n_235),
.Y(n_330)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_250),
.Y(n_290)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_290),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_258),
.A2(n_145),
.B1(n_223),
.B2(n_222),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_261),
.A2(n_222),
.B1(n_239),
.B2(n_209),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_252),
.B(n_227),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_291),
.Y(n_315)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_256),
.A2(n_237),
.B(n_235),
.C(n_220),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_263),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_264),
.A2(n_223),
.B1(n_134),
.B2(n_146),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_248),
.A2(n_240),
.B1(n_230),
.B2(n_233),
.Y(n_303)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_304),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_302),
.A2(n_268),
.B1(n_267),
.B2(n_245),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_305),
.B(n_314),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_245),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_281),
.C(n_282),
.Y(n_350)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_263),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_313),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_276),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_302),
.A2(n_243),
.B1(n_244),
.B2(n_259),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_318),
.C(n_326),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_316),
.Y(n_356)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_276),
.Y(n_317)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_317),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_253),
.C(n_244),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_302),
.A2(n_259),
.B1(n_269),
.B2(n_253),
.Y(n_320)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_280),
.A2(n_302),
.B1(n_273),
.B2(n_286),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_321),
.A2(n_322),
.B1(n_287),
.B2(n_294),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_286),
.A2(n_269),
.B1(n_271),
.B2(n_265),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_297),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_283),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_285),
.A2(n_259),
.B1(n_246),
.B2(n_254),
.Y(n_324)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_249),
.Y(n_325)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_325),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_246),
.C(n_227),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_277),
.B(n_234),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_332),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_277),
.B(n_252),
.C(n_262),
.Y(n_328)
);

MAJx2_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_298),
.C(n_293),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_329),
.Y(n_364)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_288),
.B(n_228),
.Y(n_331)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_331),
.Y(n_365)
);

OAI32xp33_ASAP7_75t_L g332 ( 
.A1(n_288),
.A2(n_228),
.A3(n_234),
.B1(n_164),
.B2(n_201),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_191),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_315),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_338),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_318),
.B(n_278),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_341),
.B(n_346),
.Y(n_366)
);

AO22x1_ASAP7_75t_L g342 ( 
.A1(n_324),
.A2(n_284),
.B1(n_289),
.B2(n_292),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_342),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_325),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_344),
.B(n_351),
.Y(n_381)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_345),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_285),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_327),
.C(n_333),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_362),
.C(n_307),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_309),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_307),
.C(n_322),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_287),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_353),
.B(n_332),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_216),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_358),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_321),
.A2(n_303),
.B1(n_300),
.B2(n_298),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_329),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_359),
.B(n_361),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_304),
.A2(n_300),
.B1(n_290),
.B2(n_274),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_319),
.A2(n_299),
.B1(n_275),
.B2(n_296),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_314),
.B(n_301),
.C(n_157),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_328),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_367),
.B(n_369),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_375),
.B1(n_362),
.B2(n_365),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_373),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_356),
.B(n_355),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_372),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_343),
.A2(n_320),
.B(n_305),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_310),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_376),
.B(n_378),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_306),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_380),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_334),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_216),
.Y(n_379)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_379),
.Y(n_417)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_383),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_346),
.B(n_334),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_387),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_311),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_390),
.Y(n_401)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_386),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_337),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_388),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_311),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_235),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_342),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_354),
.B(n_216),
.C(n_108),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_364),
.C(n_336),
.Y(n_398)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_368),
.Y(n_394)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_206),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_366),
.C(n_377),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_402),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_348),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_354),
.C(n_340),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_408),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_382),
.A2(n_335),
.B1(n_340),
.B2(n_363),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_406),
.A2(n_389),
.B1(n_299),
.B2(n_240),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_407),
.A2(n_370),
.B1(n_393),
.B2(n_380),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_361),
.C(n_358),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_410),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_363),
.C(n_335),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_411),
.B(n_413),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_342),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_389),
.Y(n_426)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_392),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_416),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_384),
.C(n_391),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_424),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_405),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_423),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_411),
.Y(n_422)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_428),
.C(n_434),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_408),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_373),
.Y(n_424)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_425),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_140),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_404),
.Y(n_428)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_429),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_299),
.C(n_190),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_433),
.B(n_395),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_435),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_202),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_415),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_230),
.Y(n_437)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_437),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_403),
.C(n_398),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_447),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_454),
.Y(n_466)
);

OAI321xp33_ASAP7_75t_L g445 ( 
.A1(n_419),
.A2(n_413),
.A3(n_397),
.B1(n_409),
.B2(n_406),
.C(n_417),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_445),
.A2(n_120),
.B1(n_10),
.B2(n_11),
.Y(n_468)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_446),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_412),
.C(n_395),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_431),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_450),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_420),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_412),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_451),
.B(n_455),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_146),
.C(n_127),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_452),
.B(n_440),
.Y(n_457)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_458),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_448),
.B(n_418),
.C(n_436),
.Y(n_458)
);

AND2x2_ASAP7_75t_SL g459 ( 
.A(n_438),
.B(n_434),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_462),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_R g462 ( 
.A(n_449),
.B(n_426),
.C(n_433),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_442),
.A2(n_126),
.B1(n_119),
.B2(n_155),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_465),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_450),
.A2(n_119),
.B1(n_155),
.B2(n_101),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_148),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_470),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_441),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_0),
.C(n_1),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_469),
.A2(n_1),
.B(n_2),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_453),
.B(n_443),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_454),
.Y(n_472)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_472),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_461),
.A2(n_444),
.B(n_452),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_473),
.B(n_481),
.Y(n_487)
);

INVx6_ASAP7_75t_L g476 ( 
.A(n_460),
.Y(n_476)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_476),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_479),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_456),
.B(n_6),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_462),
.A2(n_10),
.B(n_13),
.Y(n_480)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_480),
.A2(n_468),
.B(n_469),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_12),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_459),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_484),
.B(n_485),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_475),
.A2(n_467),
.B(n_458),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_488),
.A2(n_471),
.B(n_477),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_466),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_490),
.A2(n_480),
.B(n_466),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_489),
.B(n_476),
.Y(n_491)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_491),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_492),
.A2(n_493),
.B(n_495),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_486),
.A2(n_487),
.B(n_483),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_494),
.A2(n_483),
.B(n_478),
.Y(n_497)
);

OAI321xp33_ASAP7_75t_L g499 ( 
.A1(n_497),
.A2(n_118),
.A3(n_39),
.B1(n_12),
.B2(n_10),
.C(n_1),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_499),
.A2(n_500),
.B(n_2),
.Y(n_501)
);

OAI321xp33_ASAP7_75t_L g500 ( 
.A1(n_496),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_498),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_501),
.B(n_3),
.Y(n_502)
);

OAI21xp33_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_5),
.B(n_185),
.Y(n_503)
);


endmodule