module real_jpeg_19868_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_1),
.A2(n_5),
.B1(n_40),
.B2(n_44),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_2),
.A2(n_3),
.B1(n_34),
.B2(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_2),
.A2(n_5),
.B1(n_34),
.B2(n_40),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_25),
.B(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_2),
.B(n_81),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_2),
.A2(n_5),
.B(n_10),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_83),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_2),
.A2(n_22),
.B(n_29),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_3),
.A2(n_8),
.B1(n_32),
.B2(n_59),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_3),
.A2(n_34),
.B(n_64),
.C(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_5),
.A2(n_10),
.B1(n_38),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_53),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_5),
.A2(n_7),
.B1(n_40),
.B2(n_42),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_5),
.A2(n_8),
.B1(n_32),
.B2(n_40),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_9),
.A2(n_59),
.B(n_62),
.C(n_65),
.Y(n_61)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_64),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_112),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_111),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_86),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_16),
.B(n_86),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_72),
.B2(n_85),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_35),
.B(n_45),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_20),
.A2(n_78),
.B1(n_91),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_20),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_20),
.B(n_141),
.C(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_20),
.A2(n_125),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_24),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_23),
.A2(n_25),
.B(n_34),
.C(n_180),
.Y(n_179)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_29),
.A2(n_34),
.B(n_38),
.C(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_31),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_33),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_34),
.B(n_54),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_34),
.B(n_39),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_36),
.A2(n_39),
.B1(n_71),
.B2(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_36),
.B(n_39),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_41),
.B(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_40),
.B(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_67),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_56),
.B2(n_66),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_49),
.B1(n_68),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_51),
.B(n_98),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_54),
.B1(n_55),
.B2(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_52),
.A2(n_53),
.B1(n_99),
.B2(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_75),
.B(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_54),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.C(n_82),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_74),
.A2(n_76),
.B1(n_173),
.B2(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_74),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_76),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_76),
.B(n_130),
.C(n_171),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_76),
.A2(n_173),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_76),
.B(n_189),
.C(n_196),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_82),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_78),
.B(n_125),
.C(n_126),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_81),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_109),
.C(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_90),
.B1(n_120),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_82),
.A2(n_90),
.B1(n_101),
.B2(n_102),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_82),
.B(n_102),
.C(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_94),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_92),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_94),
.B(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_105),
.C(n_109),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_95),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_101),
.B1(n_102),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_131),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_101),
.A2(n_102),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_102),
.B(n_156),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_134),
.Y(n_214)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_218),
.B(n_223),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_146),
.B(n_204),
.C(n_217),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_132),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_115),
.B(n_132),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_117),
.B(n_119),
.C(n_123),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_163),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_139),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.C(n_140),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_133),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_135),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_138),
.B(n_140),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_153),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_203),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_198),
.B(n_202),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_186),
.B(n_197),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_175),
.B(n_185),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_166),
.B(n_174),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_158),
.B(n_165),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_154),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B(n_164),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_177),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_183),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_187),
.B(n_188),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_195),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_205),
.B(n_206),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_215),
.B2(n_216),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_213),
.C(n_216),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_215),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_220),
.Y(n_223)
);


endmodule