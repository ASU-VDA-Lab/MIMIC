module fake_jpeg_13315_n_110 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_110);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_1),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_42),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_53),
.B(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_43),
.B1(n_42),
.B2(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_57),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_60),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_43),
.B1(n_35),
.B2(n_44),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_40),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_35),
.A3(n_16),
.B1(n_17),
.B2(n_33),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_18),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_64),
.C(n_57),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_72),
.B(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_70),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_4),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_77),
.B(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_51),
.B1(n_5),
.B2(n_6),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_4),
.B(n_5),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_6),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_63),
.B(n_20),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_76),
.B(n_77),
.C(n_74),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_7),
.B(n_8),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_88),
.B(n_22),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_26),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_89),
.B1(n_27),
.B2(n_28),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_31),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_13),
.B1(n_14),
.B2(n_19),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_97),
.B1(n_98),
.B2(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_96),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_29),
.B(n_30),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

AO221x1_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_81),
.B1(n_91),
.B2(n_82),
.C(n_83),
.Y(n_104)
);

OAI321xp33_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_91),
.A3(n_79),
.B1(n_85),
.B2(n_98),
.C(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_88),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_99),
.B(n_101),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_102),
.B(n_100),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_86),
.Y(n_110)
);


endmodule