module fake_netlist_5_2567_n_2388 (n_137, n_676, n_294, n_431, n_318, n_380, n_419, n_653, n_611, n_444, n_642, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_684, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_61, n_678, n_664, n_376, n_697, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_667, n_515, n_57, n_353, n_351, n_367, n_620, n_643, n_452, n_397, n_493, n_111, n_525, n_703, n_698, n_483, n_544, n_683, n_155, n_649, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_672, n_4, n_378, n_551, n_17, n_581, n_688, n_382, n_554, n_254, n_690, n_33, n_23, n_583, n_671, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_674, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_689, n_606, n_559, n_275, n_640, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_692, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_668, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_659, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_650, n_320, n_694, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_658, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_654, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_138, n_264, n_109, n_669, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_696, n_215, n_350, n_196, n_662, n_459, n_646, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_670, n_15, n_336, n_584, n_681, n_591, n_145, n_48, n_521, n_614, n_663, n_50, n_337, n_430, n_313, n_631, n_673, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_675, n_296, n_613, n_241, n_637, n_357, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_691, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_638, n_700, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_652, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_648, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_641, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_695, n_180, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_702, n_285, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_159, n_334, n_599, n_541, n_391, n_701, n_434, n_645, n_539, n_175, n_538, n_666, n_262, n_238, n_639, n_99, n_687, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_706, n_256, n_305, n_533, n_52, n_278, n_110, n_2388);

input n_137;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_684;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_61;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_667;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_703;
input n_698;
input n_483;
input n_544;
input n_683;
input n_155;
input n_649;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_672;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_674;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_689;
input n_606;
input n_559;
input n_275;
input n_640;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_692;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_668;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_659;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_650;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_658;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_654;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_215;
input n_350;
input n_196;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_670;
input n_15;
input n_336;
input n_584;
input n_681;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_675;
input n_296;
input n_613;
input n_241;
input n_637;
input n_357;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_691;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_638;
input n_700;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_648;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_641;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_695;
input n_180;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_702;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_175;
input n_538;
input n_666;
input n_262;
input n_238;
input n_639;
input n_99;
input n_687;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_706;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2388;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_880;
wire n_1007;
wire n_2369;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_1939;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2085;
wire n_1669;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_897;
wire n_798;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_1513;
wire n_1600;
wire n_845;
wire n_2235;
wire n_1862;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_1473;
wire n_1587;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_793;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_1884;
wire n_1038;
wire n_1369;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_809;
wire n_870;
wire n_931;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_868;
wire n_914;
wire n_2120;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_913;
wire n_1537;
wire n_865;
wire n_2227;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_1333;
wire n_1121;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_738;
wire n_1624;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_1760;
wire n_936;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_959;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_1079;
wire n_2093;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_1431;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_1800;
wire n_1548;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_1237;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_1552;
wire n_1435;
wire n_879;
wire n_2088;
wire n_824;
wire n_1645;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_1553;
wire n_1811;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_912;
wire n_968;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_1974;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_984;
wire n_2082;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_1671;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_1802;
wire n_849;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_1174;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_710;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2003;
wire n_766;
wire n_1457;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_2103;
wire n_2160;
wire n_2228;
wire n_1602;
wire n_1178;
wire n_855;
wire n_1461;
wire n_850;
wire n_2286;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_1273;
wire n_1822;
wire n_2363;
wire n_916;
wire n_1081;
wire n_2332;
wire n_1235;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_1172;
wire n_1341;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_1589;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_1337;
wire n_1495;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2083;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_2044;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_78),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_422),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_437),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_332),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_96),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_60),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_555),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_404),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_312),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_347),
.Y(n_718)
);

CKINVDCx16_ASAP7_75t_R g719 ( 
.A(n_698),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_492),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_226),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_309),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_287),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_353),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_398),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_602),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_379),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_355),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_502),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_659),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_536),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_252),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_37),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_110),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_702),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_238),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_212),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_159),
.Y(n_738)
);

CKINVDCx16_ASAP7_75t_R g739 ( 
.A(n_630),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_393),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_188),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_662),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_663),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_157),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_586),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_436),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_186),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_304),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_680),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_119),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_504),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_417),
.Y(n_752)
);

CKINVDCx14_ASAP7_75t_R g753 ( 
.A(n_6),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_72),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_20),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_669),
.Y(n_756)
);

INVx1_ASAP7_75t_SL g757 ( 
.A(n_391),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_518),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_59),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_122),
.Y(n_760)
);

BUFx8_ASAP7_75t_SL g761 ( 
.A(n_627),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_650),
.Y(n_762)
);

BUFx10_ASAP7_75t_L g763 ( 
.A(n_32),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_89),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_263),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_138),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_449),
.Y(n_767)
);

CKINVDCx11_ASAP7_75t_R g768 ( 
.A(n_479),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_52),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_666),
.Y(n_770)
);

BUFx10_ASAP7_75t_L g771 ( 
.A(n_448),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_656),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_647),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_668),
.Y(n_774)
);

CKINVDCx14_ASAP7_75t_R g775 ( 
.A(n_316),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_313),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_511),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_507),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_503),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_204),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_164),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_168),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_397),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_472),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_661),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_544),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_658),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_657),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_0),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_477),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_588),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_185),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_6),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_221),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_200),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_311),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_127),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_361),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_249),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_665),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_107),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_257),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_653),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_86),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_350),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_297),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_368),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_413),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_346),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_75),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_468),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_380),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_505),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_143),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_703),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_629),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_23),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_673),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_648),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_426),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_187),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_396),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_651),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_655),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_539),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_258),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_371),
.Y(n_827)
);

BUFx10_ASAP7_75t_L g828 ( 
.A(n_352),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_581),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_300),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_687),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_101),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_522),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_45),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_452),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_93),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_369),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_646),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_310),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_642),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_55),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_438),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_27),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_402),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_667),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_575),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_14),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_245),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_670),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_675),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_556),
.Y(n_851)
);

BUFx8_ASAP7_75t_SL g852 ( 
.A(n_35),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_184),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_128),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_654),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_314),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_88),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_14),
.Y(n_858)
);

BUFx8_ASAP7_75t_SL g859 ( 
.A(n_491),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_547),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_557),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_455),
.Y(n_862)
);

CKINVDCx14_ASAP7_75t_R g863 ( 
.A(n_645),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_315),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_94),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_490),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_61),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_652),
.Y(n_868)
);

CKINVDCx14_ASAP7_75t_R g869 ( 
.A(n_381),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_672),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_664),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_321),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_563),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_660),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_498),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_36),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_390),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_306),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_644),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_649),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_420),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_388),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_251),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_593),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_832),
.Y(n_885)
);

INVxp33_ASAP7_75t_SL g886 ( 
.A(n_843),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_832),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_832),
.Y(n_888)
);

NOR2xp67_ASAP7_75t_L g889 ( 
.A(n_713),
.B(n_0),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_734),
.Y(n_890)
);

CKINVDCx16_ASAP7_75t_R g891 ( 
.A(n_719),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_750),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_759),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_789),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_801),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_804),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_867),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_876),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_733),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_761),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_710),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_771),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_717),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_814),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_720),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_725),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_729),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_731),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_735),
.Y(n_909)
);

CKINVDCx14_ASAP7_75t_R g910 ( 
.A(n_753),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_736),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_742),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_749),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_762),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_859),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_774),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_765),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_780),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_852),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_768),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_795),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_763),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_799),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_763),
.Y(n_924)
);

CKINVDCx16_ASAP7_75t_R g925 ( 
.A(n_739),
.Y(n_925)
);

NOR2xp67_ASAP7_75t_L g926 ( 
.A(n_817),
.B(n_1),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_808),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_805),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_818),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_822),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_709),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_771),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_837),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_839),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_844),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_850),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_853),
.Y(n_937)
);

INVxp33_ASAP7_75t_SL g938 ( 
.A(n_714),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_860),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_861),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_754),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_836),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_858),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_862),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_870),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_711),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_879),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_715),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_882),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_728),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_884),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_774),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_783),
.Y(n_953)
);

CKINVDCx16_ASAP7_75t_R g954 ( 
.A(n_775),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_820),
.Y(n_955)
);

INVxp67_ASAP7_75t_SL g956 ( 
.A(n_830),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_824),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_774),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_873),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_755),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_877),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_716),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_712),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_840),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_760),
.B(n_1),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_740),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_792),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_803),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_833),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_868),
.Y(n_970)
);

NOR2xp67_ASAP7_75t_L g971 ( 
.A(n_764),
.B(n_2),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_769),
.Y(n_972)
);

INVxp67_ASAP7_75t_L g973 ( 
.A(n_793),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_718),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_806),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_810),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_834),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_841),
.B(n_2),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_847),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_854),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_825),
.Y(n_981)
);

INVxp67_ASAP7_75t_SL g982 ( 
.A(n_871),
.Y(n_982)
);

CKINVDCx16_ASAP7_75t_R g983 ( 
.A(n_863),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_857),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_865),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_916),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_916),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_985),
.B(n_878),
.Y(n_988)
);

AND2x6_ASAP7_75t_L g989 ( 
.A(n_975),
.B(n_757),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_885),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_886),
.A2(n_869),
.B1(n_849),
.B2(n_766),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_938),
.B(n_777),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_887),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_902),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_916),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_932),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_981),
.A2(n_797),
.B1(n_767),
.B2(n_782),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_946),
.B(n_948),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_954),
.B(n_806),
.Y(n_999)
);

INVx5_ASAP7_75t_L g1000 ( 
.A(n_952),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_972),
.B(n_748),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_888),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_952),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_900),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_952),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_962),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_984),
.B(n_721),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_974),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_958),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_958),
.Y(n_1010)
);

CKINVDCx11_ASAP7_75t_R g1011 ( 
.A(n_928),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_976),
.B(n_722),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_941),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_950),
.Y(n_1014)
);

BUFx8_ASAP7_75t_L g1015 ( 
.A(n_979),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_982),
.A2(n_724),
.B1(n_726),
.B2(n_723),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_958),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_898),
.Y(n_1018)
);

OA21x2_ASAP7_75t_L g1019 ( 
.A1(n_968),
.A2(n_730),
.B(n_727),
.Y(n_1019)
);

BUFx12f_ASAP7_75t_L g1020 ( 
.A(n_915),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_899),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_942),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_943),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_890),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_892),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_980),
.B(n_732),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_901),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_903),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_905),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_893),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_931),
.B(n_737),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_894),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_960),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_895),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_973),
.B(n_738),
.Y(n_1035)
);

AND2x6_ASAP7_75t_L g1036 ( 
.A(n_953),
.B(n_828),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_955),
.Y(n_1037)
);

BUFx12f_ASAP7_75t_L g1038 ( 
.A(n_920),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_956),
.B(n_741),
.Y(n_1039)
);

INVx6_ASAP7_75t_L g1040 ( 
.A(n_891),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_896),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_957),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_897),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_910),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_963),
.Y(n_1045)
);

CKINVDCx8_ASAP7_75t_R g1046 ( 
.A(n_925),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_977),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_922),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_966),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_983),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_SL g1051 ( 
.A(n_924),
.B(n_828),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_967),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_906),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_907),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_959),
.B(n_866),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_961),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_978),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_908),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_909),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_911),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_912),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_969),
.Y(n_1062)
);

INVx6_ASAP7_75t_L g1063 ( 
.A(n_904),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_913),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_964),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_914),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_970),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_917),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_918),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_919),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_921),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_987),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1014),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_987),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1021),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1027),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1021),
.Y(n_1077)
);

NAND2xp33_ASAP7_75t_SL g1078 ( 
.A(n_1057),
.B(n_743),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_SL g1079 ( 
.A(n_1033),
.B(n_744),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1028),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1022),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1029),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1022),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1023),
.B(n_923),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1054),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1068),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_992),
.B(n_965),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_995),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1053),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_986),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1005),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1053),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1009),
.Y(n_1093)
);

INVxp33_ASAP7_75t_SL g1094 ( 
.A(n_1051),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_1063),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1058),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_1013),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1001),
.B(n_971),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1058),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1059),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1059),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_998),
.B(n_927),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_1007),
.B(n_889),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1055),
.B(n_929),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1060),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_995),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1006),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_1050),
.B(n_949),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_1003),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1060),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_1061),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_1061),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1010),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_1039),
.B(n_752),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1045),
.B(n_930),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1024),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1018),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_1024),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1017),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_1008),
.Y(n_1120)
);

INVx3_ASAP7_75t_L g1121 ( 
.A(n_1025),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_1040),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1066),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1025),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1012),
.B(n_933),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1030),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1026),
.B(n_934),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1047),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1016),
.B(n_756),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1030),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_990),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1034),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_993),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1034),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1041),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1048),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1041),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1019),
.B(n_935),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1000),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1071),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1000),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_994),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_996),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1031),
.B(n_936),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1037),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_1042),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1032),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1043),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_989),
.Y(n_1149)
);

NAND2xp33_ASAP7_75t_L g1150 ( 
.A(n_1036),
.B(n_745),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1002),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1035),
.B(n_926),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1049),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1064),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1056),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1052),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1069),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1062),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1067),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_988),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_997),
.B(n_937),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1044),
.B(n_939),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_989),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1070),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_999),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1102),
.B(n_991),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_1122),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1136),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1098),
.B(n_1046),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1104),
.B(n_1036),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1161),
.A2(n_944),
.B1(n_945),
.B2(n_940),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_1095),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1163),
.B(n_883),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1138),
.A2(n_951),
.B1(n_947),
.B2(n_747),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1084),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_1162),
.Y(n_1176)
);

BUFx10_ASAP7_75t_L g1177 ( 
.A(n_1164),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1076),
.B(n_1080),
.Y(n_1178)
);

OR2x6_ASAP7_75t_L g1179 ( 
.A(n_1163),
.B(n_1038),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1082),
.B(n_746),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1165),
.B(n_751),
.Y(n_1181)
);

INVx4_ASAP7_75t_L g1182 ( 
.A(n_1122),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1097),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1094),
.B(n_1065),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1085),
.B(n_1086),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1087),
.B(n_1015),
.C(n_770),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1075),
.B(n_845),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1084),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1117),
.B(n_758),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1144),
.B(n_772),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1125),
.B(n_1127),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1128),
.Y(n_1192)
);

AND2x6_ASAP7_75t_L g1193 ( 
.A(n_1152),
.B(n_1004),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1115),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1115),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1160),
.B(n_1011),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_1109),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1153),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1146),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1140),
.B(n_773),
.Y(n_1200)
);

INVx4_ASAP7_75t_SL g1201 ( 
.A(n_1103),
.Y(n_1201)
);

NAND2x1p5_ASAP7_75t_L g1202 ( 
.A(n_1146),
.B(n_1020),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1129),
.A2(n_778),
.B1(n_779),
.B2(n_776),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1112),
.B(n_872),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1149),
.B(n_781),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1109),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1107),
.B(n_784),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1120),
.B(n_785),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1131),
.A2(n_1151),
.B1(n_1133),
.B2(n_1148),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1147),
.A2(n_787),
.B1(n_788),
.B2(n_786),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1158),
.Y(n_1211)
);

BUFx4f_ASAP7_75t_L g1212 ( 
.A(n_1108),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1112),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1124),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1073),
.B(n_790),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1124),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1159),
.Y(n_1217)
);

AND2x6_ASAP7_75t_L g1218 ( 
.A(n_1123),
.B(n_150),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1090),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1091),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_1141),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1154),
.A2(n_794),
.B1(n_796),
.B2(n_791),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1132),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1143),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1132),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1079),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1157),
.B(n_798),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1072),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1142),
.B(n_1155),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1093),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1113),
.B(n_800),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1156),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1119),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1078),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1156),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1145),
.B(n_802),
.Y(n_1236)
);

INVxp67_ASAP7_75t_SL g1237 ( 
.A(n_1111),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1116),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1077),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1081),
.Y(n_1240)
);

INVx5_ASAP7_75t_L g1241 ( 
.A(n_1141),
.Y(n_1241)
);

AND2x2_ASAP7_75t_SL g1242 ( 
.A(n_1150),
.B(n_1083),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1089),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1092),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1118),
.B(n_856),
.Y(n_1245)
);

BUFx10_ASAP7_75t_L g1246 ( 
.A(n_1096),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1121),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1072),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1114),
.B(n_874),
.C(n_864),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1099),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1100),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1101),
.Y(n_1252)
);

BUFx4f_ASAP7_75t_L g1253 ( 
.A(n_1074),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1105),
.B(n_807),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1110),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1130),
.B(n_809),
.Y(n_1256)
);

OR2x6_ASAP7_75t_L g1257 ( 
.A(n_1126),
.B(n_3),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1134),
.B(n_881),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1074),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1135),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1137),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1088),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1088),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1106),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1191),
.B(n_811),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1212),
.B(n_812),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1248),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1219),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1170),
.B(n_813),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1175),
.B(n_815),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1188),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1166),
.B(n_1139),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1184),
.B(n_816),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1194),
.B(n_819),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1230),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1195),
.B(n_821),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1198),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1178),
.B(n_1185),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1174),
.B(n_823),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1211),
.Y(n_1280)
);

OR2x6_ASAP7_75t_L g1281 ( 
.A(n_1179),
.B(n_3),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1192),
.B(n_826),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1190),
.B(n_827),
.Y(n_1283)
);

BUFx8_ASAP7_75t_L g1284 ( 
.A(n_1168),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1183),
.B(n_829),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1217),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1207),
.B(n_831),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1229),
.B(n_835),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1224),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1208),
.B(n_838),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1220),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1234),
.B(n_842),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1233),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1244),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1176),
.B(n_846),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1205),
.B(n_848),
.Y(n_1296)
);

O2A1O1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1181),
.A2(n_855),
.B(n_875),
.C(n_851),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1180),
.B(n_880),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1240),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1209),
.B(n_4),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1242),
.B(n_4),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1250),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1189),
.B(n_5),
.Y(n_1303)
);

NAND2xp33_ASAP7_75t_L g1304 ( 
.A(n_1218),
.B(n_151),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1171),
.B(n_5),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1252),
.Y(n_1306)
);

AOI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1226),
.A2(n_153),
.B1(n_154),
.B2(n_152),
.Y(n_1307)
);

INVx8_ASAP7_75t_L g1308 ( 
.A(n_1221),
.Y(n_1308)
);

OR2x6_ASAP7_75t_L g1309 ( 
.A(n_1179),
.B(n_7),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1251),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1215),
.B(n_7),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1200),
.B(n_8),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1255),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1172),
.Y(n_1314)
);

INVx8_ASAP7_75t_L g1315 ( 
.A(n_1221),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_SL g1316 ( 
.A(n_1177),
.B(n_155),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1236),
.B(n_8),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1260),
.Y(n_1318)
);

NOR2xp67_ASAP7_75t_L g1319 ( 
.A(n_1167),
.B(n_156),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1261),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1227),
.B(n_9),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1237),
.B(n_9),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1239),
.B(n_10),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1232),
.B(n_10),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1235),
.B(n_11),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1231),
.B(n_11),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1243),
.B(n_12),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1199),
.B(n_12),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1262),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_SL g1330 ( 
.A(n_1203),
.B(n_1249),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1222),
.B(n_13),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1169),
.B(n_158),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1254),
.B(n_160),
.Y(n_1333)
);

AO221x1_ASAP7_75t_L g1334 ( 
.A1(n_1228),
.A2(n_16),
.B1(n_13),
.B2(n_15),
.C(n_17),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1256),
.B(n_161),
.Y(n_1335)
);

INVxp67_ASAP7_75t_SL g1336 ( 
.A(n_1248),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1253),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1201),
.B(n_162),
.Y(n_1338)
);

AND2x2_ASAP7_75t_SL g1339 ( 
.A(n_1182),
.B(n_15),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1173),
.B(n_16),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1238),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1214),
.Y(n_1342)
);

AO22x2_ASAP7_75t_L g1343 ( 
.A1(n_1186),
.A2(n_25),
.B1(n_33),
.B2(n_17),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1278),
.B(n_1196),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1284),
.Y(n_1345)
);

BUFx12f_ASAP7_75t_SL g1346 ( 
.A(n_1337),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1265),
.B(n_1210),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1273),
.A2(n_1258),
.B1(n_1187),
.B2(n_1204),
.Y(n_1348)
);

NAND2x1p5_ASAP7_75t_L g1349 ( 
.A(n_1267),
.B(n_1225),
.Y(n_1349)
);

INVxp67_ASAP7_75t_L g1350 ( 
.A(n_1289),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1271),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1268),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1308),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1288),
.B(n_1218),
.Y(n_1354)
);

NAND2xp33_ASAP7_75t_L g1355 ( 
.A(n_1311),
.B(n_1218),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1294),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1276),
.B(n_1201),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1272),
.B(n_1246),
.Y(n_1358)
);

INVxp67_ASAP7_75t_SL g1359 ( 
.A(n_1314),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1287),
.B(n_1213),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1337),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1292),
.A2(n_1245),
.B1(n_1193),
.B2(n_1223),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1302),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1290),
.B(n_1216),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1308),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1275),
.Y(n_1366)
);

INVx4_ASAP7_75t_L g1367 ( 
.A(n_1315),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1315),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1331),
.A2(n_1257),
.B1(n_1247),
.B2(n_1193),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1277),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1330),
.A2(n_1193),
.B1(n_1257),
.B2(n_1259),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1305),
.A2(n_1264),
.B1(n_1263),
.B2(n_1206),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1310),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1341),
.B(n_1197),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1301),
.A2(n_1264),
.B1(n_1202),
.B2(n_1241),
.Y(n_1375)
);

AND2x6_ASAP7_75t_L g1376 ( 
.A(n_1338),
.B(n_1241),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1285),
.B(n_1282),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1267),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1283),
.B(n_18),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1291),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1317),
.B(n_163),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1270),
.B(n_18),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1328),
.B(n_19),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1342),
.B(n_1336),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1313),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1339),
.B(n_19),
.Y(n_1386)
);

BUFx12f_ASAP7_75t_L g1387 ( 
.A(n_1281),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1320),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1296),
.B(n_20),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1293),
.B(n_21),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1318),
.B(n_165),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1312),
.B(n_21),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1329),
.B(n_166),
.Y(n_1393)
);

BUFx2_ASAP7_75t_SL g1394 ( 
.A(n_1319),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1327),
.B(n_22),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1280),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1286),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1321),
.B(n_22),
.Y(n_1398)
);

INVx5_ASAP7_75t_L g1399 ( 
.A(n_1281),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1306),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1300),
.B(n_23),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1324),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1309),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1299),
.Y(n_1404)
);

OR2x2_ASAP7_75t_SL g1405 ( 
.A(n_1279),
.B(n_24),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1303),
.B(n_24),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1274),
.B(n_167),
.Y(n_1407)
);

NOR3xp33_ASAP7_75t_SL g1408 ( 
.A(n_1340),
.B(n_25),
.C(n_26),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1309),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1322),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1326),
.B(n_26),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1323),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1332),
.B(n_169),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1325),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1266),
.B(n_170),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1298),
.B(n_28),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1269),
.B(n_29),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1295),
.B(n_30),
.Y(n_1418)
);

AND3x2_ASAP7_75t_SL g1419 ( 
.A(n_1343),
.B(n_30),
.C(n_31),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1334),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1377),
.B(n_1316),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1356),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1344),
.B(n_1343),
.Y(n_1423)
);

AND2x4_ASAP7_75t_SL g1424 ( 
.A(n_1367),
.B(n_1307),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1363),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1373),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1410),
.B(n_1333),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1378),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1385),
.Y(n_1429)
);

INVx4_ASAP7_75t_L g1430 ( 
.A(n_1378),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1386),
.B(n_1335),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_SL g1432 ( 
.A(n_1399),
.B(n_1297),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1350),
.B(n_1304),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1388),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1414),
.B(n_31),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1351),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1349),
.Y(n_1437)
);

NOR2xp67_ASAP7_75t_L g1438 ( 
.A(n_1362),
.B(n_171),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1383),
.B(n_32),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1399),
.B(n_1402),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1382),
.B(n_33),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1370),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1353),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1380),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1395),
.B(n_34),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1397),
.Y(n_1446)
);

NAND2x1p5_ASAP7_75t_L g1447 ( 
.A(n_1365),
.B(n_176),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1402),
.B(n_34),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1396),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_R g1450 ( 
.A(n_1346),
.B(n_172),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1368),
.Y(n_1451)
);

AND2x2_ASAP7_75t_SL g1452 ( 
.A(n_1415),
.B(n_35),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1361),
.B(n_173),
.Y(n_1453)
);

NAND2xp33_ASAP7_75t_SL g1454 ( 
.A(n_1357),
.B(n_36),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1420),
.B(n_37),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1400),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1374),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1360),
.B(n_38),
.Y(n_1458)
);

INVx3_ASAP7_75t_SL g1459 ( 
.A(n_1403),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_SL g1460 ( 
.A(n_1348),
.B(n_38),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1347),
.B(n_39),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1384),
.B(n_174),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1359),
.B(n_175),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1364),
.B(n_39),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1379),
.B(n_40),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1352),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1366),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1404),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1390),
.Y(n_1469)
);

AO22x1_ASAP7_75t_L g1470 ( 
.A1(n_1376),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1389),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1471)
);

INVx5_ASAP7_75t_L g1472 ( 
.A(n_1376),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1401),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1392),
.B(n_43),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1398),
.B(n_44),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1406),
.B(n_44),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1345),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1393),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1411),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1409),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1417),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1418),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1358),
.B(n_45),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1416),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1391),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1376),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1394),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1412),
.Y(n_1488)
);

AND2x2_ASAP7_75t_SL g1489 ( 
.A(n_1419),
.B(n_46),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1387),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1413),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1405),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1407),
.Y(n_1493)
);

NAND2xp33_ASAP7_75t_L g1494 ( 
.A(n_1354),
.B(n_177),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1381),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1371),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1372),
.Y(n_1497)
);

AND2x2_ASAP7_75t_SL g1498 ( 
.A(n_1355),
.B(n_47),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1408),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1375),
.B(n_178),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1369),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1356),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1430),
.B(n_179),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_48),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1480),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1452),
.B(n_49),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1495),
.A2(n_1485),
.B(n_1432),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1494),
.A2(n_1421),
.B(n_1460),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1488),
.A2(n_181),
.B(n_180),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1479),
.B(n_49),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1496),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1428),
.Y(n_1512)
);

O2A1O1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1441),
.A2(n_53),
.B(n_50),
.C(n_51),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1422),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_SL g1515 ( 
.A(n_1433),
.B(n_53),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1455),
.A2(n_183),
.B(n_182),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1427),
.B(n_54),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1469),
.B(n_189),
.Y(n_1518)
);

AO31x2_ASAP7_75t_L g1519 ( 
.A1(n_1423),
.A2(n_191),
.A3(n_192),
.B(n_190),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1451),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1457),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1449),
.A2(n_194),
.B(n_193),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1434),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1438),
.A2(n_701),
.B(n_700),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1456),
.A2(n_196),
.B(n_195),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1425),
.A2(n_198),
.B(n_197),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1501),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1431),
.A2(n_690),
.B(n_689),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1436),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1493),
.A2(n_201),
.B(n_199),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1426),
.A2(n_203),
.B(n_202),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1477),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1481),
.B(n_56),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1429),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1484),
.B(n_57),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1482),
.B(n_57),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1500),
.B(n_58),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1461),
.A2(n_699),
.B(n_697),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1465),
.A2(n_206),
.B(n_205),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1492),
.B(n_207),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1499),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.C(n_61),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1454),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1542)
);

OAI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1458),
.A2(n_62),
.B(n_63),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1498),
.A2(n_691),
.B(n_688),
.Y(n_1544)
);

NAND2x1p5_ASAP7_75t_L g1545 ( 
.A(n_1472),
.B(n_208),
.Y(n_1545)
);

A2O1A1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1474),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_1546)
);

NAND2x1_ASAP7_75t_L g1547 ( 
.A(n_1493),
.B(n_209),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1464),
.A2(n_696),
.B(n_695),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1502),
.A2(n_211),
.B(n_210),
.Y(n_1549)
);

NOR2x1_ASAP7_75t_L g1550 ( 
.A(n_1487),
.B(n_213),
.Y(n_1550)
);

NOR2xp67_ASAP7_75t_L g1551 ( 
.A(n_1472),
.B(n_214),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1466),
.A2(n_216),
.B(n_215),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1467),
.A2(n_1468),
.B(n_1475),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1442),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1435),
.B(n_65),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1476),
.B(n_66),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1497),
.A2(n_1478),
.B1(n_1489),
.B2(n_1424),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1444),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1445),
.B(n_67),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1446),
.A2(n_1447),
.B(n_1440),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1462),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1448),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1483),
.A2(n_218),
.B(n_217),
.Y(n_1563)
);

NAND2x1_ASAP7_75t_L g1564 ( 
.A(n_1486),
.B(n_219),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1439),
.B(n_67),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1463),
.B(n_68),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1472),
.A2(n_1491),
.B1(n_1437),
.B2(n_1471),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1453),
.B(n_68),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1459),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1569)
);

NAND3xp33_ASAP7_75t_SL g1570 ( 
.A(n_1450),
.B(n_69),
.C(n_70),
.Y(n_1570)
);

AO22x2_ASAP7_75t_L g1571 ( 
.A1(n_1470),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1451),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1443),
.B(n_73),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1490),
.A2(n_74),
.B(n_75),
.Y(n_1574)
);

OA22x2_ASAP7_75t_L g1575 ( 
.A1(n_1499),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1494),
.A2(n_708),
.B(n_222),
.Y(n_1576)
);

NOR2xp67_ASAP7_75t_L g1577 ( 
.A(n_1472),
.B(n_220),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1421),
.A2(n_76),
.B(n_77),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1430),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1473),
.B(n_78),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1496),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_1581)
);

OAI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1421),
.A2(n_79),
.B(n_80),
.Y(n_1582)
);

OAI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1421),
.A2(n_81),
.B(n_82),
.Y(n_1583)
);

AOI21x1_ASAP7_75t_SL g1584 ( 
.A1(n_1441),
.A2(n_82),
.B(n_83),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1421),
.A2(n_83),
.B(n_84),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1422),
.Y(n_1586)
);

OA22x2_ASAP7_75t_L g1587 ( 
.A1(n_1499),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1473),
.B(n_85),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1494),
.A2(n_706),
.B(n_705),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1421),
.A2(n_87),
.B(n_88),
.Y(n_1590)
);

OAI21x1_ASAP7_75t_L g1591 ( 
.A1(n_1495),
.A2(n_224),
.B(n_223),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1495),
.A2(n_227),
.B(n_225),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1473),
.B(n_87),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1473),
.B(n_89),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1495),
.A2(n_229),
.B(n_228),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1422),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1473),
.B(n_90),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1494),
.A2(n_685),
.B(n_684),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1422),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1495),
.A2(n_231),
.B(n_230),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1473),
.B(n_90),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1421),
.B(n_91),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1480),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1473),
.B(n_91),
.Y(n_1604)
);

AO21x1_ASAP7_75t_L g1605 ( 
.A1(n_1441),
.A2(n_92),
.B(n_93),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1473),
.B(n_92),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1473),
.B(n_94),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1430),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1452),
.B(n_95),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1473),
.B(n_95),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1495),
.A2(n_233),
.B(n_232),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1422),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_SL g1613 ( 
.A1(n_1455),
.A2(n_96),
.B(n_97),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1494),
.A2(n_707),
.B(n_235),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1494),
.A2(n_704),
.B(n_236),
.Y(n_1615)
);

NAND2x1p5_ASAP7_75t_L g1616 ( 
.A(n_1472),
.B(n_234),
.Y(n_1616)
);

INVx4_ASAP7_75t_L g1617 ( 
.A(n_1472),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1421),
.A2(n_97),
.B(n_98),
.Y(n_1618)
);

AO31x2_ASAP7_75t_L g1619 ( 
.A1(n_1488),
.A2(n_239),
.A3(n_240),
.B(n_237),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1494),
.A2(n_242),
.B(n_241),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1523),
.B(n_98),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_SL g1622 ( 
.A(n_1608),
.B(n_243),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1534),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1603),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1562),
.B(n_99),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1602),
.B(n_99),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1572),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1517),
.B(n_100),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1514),
.B(n_100),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1529),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1515),
.B(n_101),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1506),
.B(n_244),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1609),
.B(n_246),
.Y(n_1633)
);

BUFx12f_ASAP7_75t_L g1634 ( 
.A(n_1532),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1558),
.B(n_247),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1554),
.B(n_102),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1561),
.B(n_248),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_R g1638 ( 
.A(n_1520),
.B(n_694),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1586),
.B(n_1596),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1557),
.B(n_250),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1599),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1512),
.B(n_253),
.Y(n_1642)
);

NAND2xp33_ASAP7_75t_L g1643 ( 
.A(n_1578),
.B(n_102),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1521),
.Y(n_1644)
);

INVx5_ASAP7_75t_L g1645 ( 
.A(n_1572),
.Y(n_1645)
);

NAND3xp33_ASAP7_75t_L g1646 ( 
.A(n_1543),
.B(n_103),
.C(n_104),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1509),
.A2(n_255),
.B(n_254),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1570),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1648)
);

BUFx12f_ASAP7_75t_L g1649 ( 
.A(n_1579),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1612),
.B(n_105),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1559),
.B(n_256),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1518),
.B(n_1555),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1537),
.B(n_1504),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1553),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1505),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1566),
.B(n_259),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1510),
.B(n_106),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1508),
.B(n_260),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1568),
.B(n_261),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1579),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1580),
.B(n_106),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1507),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1573),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1588),
.B(n_107),
.Y(n_1664)
);

BUFx3_ASAP7_75t_L g1665 ( 
.A(n_1503),
.Y(n_1665)
);

INVx4_ASAP7_75t_L g1666 ( 
.A(n_1617),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1560),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1533),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1551),
.B(n_262),
.Y(n_1669)
);

INVx3_ASAP7_75t_SL g1670 ( 
.A(n_1575),
.Y(n_1670)
);

NAND2x1p5_ASAP7_75t_L g1671 ( 
.A(n_1547),
.B(n_264),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1567),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1535),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1576),
.A2(n_266),
.B(n_265),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_SL g1675 ( 
.A(n_1540),
.B(n_267),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1577),
.B(n_268),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1536),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1565),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1589),
.A2(n_270),
.B(n_269),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1556),
.B(n_271),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1587),
.B(n_272),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1550),
.B(n_273),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1542),
.A2(n_111),
.B1(n_108),
.B2(n_109),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1593),
.Y(n_1685)
);

O2A1O1Ixp33_ASAP7_75t_L g1686 ( 
.A1(n_1585),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1564),
.Y(n_1687)
);

OR2x6_ASAP7_75t_SL g1688 ( 
.A(n_1569),
.B(n_1594),
.Y(n_1688)
);

OR2x6_ASAP7_75t_L g1689 ( 
.A(n_1530),
.B(n_274),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1597),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1598),
.A2(n_276),
.B(n_275),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1614),
.A2(n_1620),
.B(n_1615),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1601),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1604),
.B(n_112),
.Y(n_1694)
);

O2A1O1Ixp5_ASAP7_75t_L g1695 ( 
.A1(n_1590),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1618),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1606),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1545),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1607),
.B(n_1610),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1591),
.Y(n_1700)
);

NAND2x1p5_ASAP7_75t_L g1701 ( 
.A(n_1516),
.B(n_277),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1616),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1592),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1571),
.B(n_278),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1519),
.Y(n_1705)
);

INVx3_ASAP7_75t_SL g1706 ( 
.A(n_1539),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1538),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1595),
.B(n_279),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1581),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1519),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1563),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1541),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1544),
.B(n_280),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1600),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1605),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1546),
.B(n_120),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1513),
.B(n_120),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1619),
.Y(n_1718)
);

A2O1A1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1574),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1511),
.B(n_281),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1524),
.A2(n_283),
.B(n_282),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1611),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1528),
.A2(n_124),
.B(n_121),
.C(n_123),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1644),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1649),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1668),
.B(n_1571),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1623),
.B(n_1619),
.Y(n_1727)
);

O2A1O1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1643),
.A2(n_1527),
.B(n_1613),
.C(n_1548),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1673),
.B(n_1522),
.Y(n_1729)
);

INVxp67_ASAP7_75t_L g1730 ( 
.A(n_1655),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1624),
.B(n_1525),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1670),
.A2(n_1584),
.B1(n_1531),
.B2(n_1549),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1639),
.B(n_1526),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1697),
.B(n_1630),
.Y(n_1734)
);

OR2x6_ASAP7_75t_SL g1735 ( 
.A(n_1685),
.B(n_1552),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1641),
.B(n_124),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1677),
.B(n_125),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1632),
.B(n_125),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1633),
.B(n_126),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1645),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1654),
.Y(n_1741)
);

OA21x2_ASAP7_75t_L g1742 ( 
.A1(n_1718),
.A2(n_126),
.B(n_127),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1705),
.Y(n_1743)
);

O2A1O1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1719),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_1744)
);

NOR2x2_ASAP7_75t_L g1745 ( 
.A(n_1689),
.B(n_129),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1690),
.B(n_130),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1662),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1710),
.Y(n_1748)
);

A2O1A1Ixp33_ASAP7_75t_L g1749 ( 
.A1(n_1686),
.A2(n_133),
.B(n_131),
.C(n_132),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1696),
.A2(n_1682),
.B(n_1723),
.C(n_1717),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1667),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1693),
.B(n_131),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1715),
.Y(n_1753)
);

BUFx2_ASAP7_75t_L g1754 ( 
.A(n_1665),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1699),
.B(n_132),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1663),
.B(n_133),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1653),
.B(n_134),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1652),
.B(n_134),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1704),
.B(n_135),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1711),
.Y(n_1760)
);

NOR2xp67_ASAP7_75t_L g1761 ( 
.A(n_1666),
.B(n_135),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_SL g1762 ( 
.A(n_1675),
.B(n_284),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1712),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1763)
);

O2A1O1Ixp5_ASAP7_75t_L g1764 ( 
.A1(n_1695),
.A2(n_139),
.B(n_136),
.C(n_137),
.Y(n_1764)
);

A2O1A1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1646),
.A2(n_141),
.B(n_139),
.C(n_140),
.Y(n_1765)
);

O2A1O1Ixp5_ASAP7_75t_L g1766 ( 
.A1(n_1684),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_1766)
);

NOR2xp67_ASAP7_75t_L g1767 ( 
.A(n_1625),
.B(n_142),
.Y(n_1767)
);

OAI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1692),
.A2(n_286),
.B(n_285),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1678),
.B(n_143),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1658),
.A2(n_289),
.B(n_288),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1650),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1651),
.B(n_144),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1648),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1636),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1628),
.B(n_145),
.Y(n_1775)
);

AOI21x1_ASAP7_75t_SL g1776 ( 
.A1(n_1716),
.A2(n_146),
.B(n_147),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1634),
.B(n_290),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_SL g1778 ( 
.A(n_1622),
.B(n_291),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1700),
.Y(n_1779)
);

A2O1A1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1672),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1621),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1629),
.B(n_148),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1703),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1688),
.A2(n_149),
.B1(n_293),
.B2(n_292),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1645),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1722),
.Y(n_1786)
);

A2O1A1Ixp33_ASAP7_75t_L g1787 ( 
.A1(n_1720),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1680),
.B(n_693),
.Y(n_1788)
);

O2A1O1Ixp33_ASAP7_75t_L g1789 ( 
.A1(n_1709),
.A2(n_301),
.B(n_298),
.C(n_299),
.Y(n_1789)
);

AND2x2_ASAP7_75t_SL g1790 ( 
.A(n_1698),
.B(n_302),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1657),
.B(n_303),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1702),
.B(n_692),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1674),
.A2(n_305),
.B(n_307),
.Y(n_1793)
);

BUFx12f_ASAP7_75t_L g1794 ( 
.A(n_1660),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1661),
.B(n_308),
.Y(n_1795)
);

A2O1A1Ixp33_ASAP7_75t_L g1796 ( 
.A1(n_1679),
.A2(n_1691),
.B(n_1640),
.C(n_1721),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1714),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1681),
.B(n_686),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1659),
.B(n_1706),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1714),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1707),
.A2(n_317),
.B(n_318),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1664),
.B(n_319),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1694),
.B(n_320),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1627),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1642),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1626),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1635),
.B(n_322),
.Y(n_1807)
);

O2A1O1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1631),
.A2(n_325),
.B(n_323),
.C(n_324),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1689),
.A2(n_326),
.B(n_327),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1656),
.B(n_328),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_L g1811 ( 
.A(n_1687),
.B(n_329),
.Y(n_1811)
);

O2A1O1Ixp5_ASAP7_75t_L g1812 ( 
.A1(n_1713),
.A2(n_333),
.B(n_330),
.C(n_331),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1683),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.C(n_337),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1637),
.B(n_683),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1701),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1647),
.B(n_338),
.Y(n_1816)
);

NAND2x1p5_ASAP7_75t_L g1817 ( 
.A(n_1669),
.B(n_339),
.Y(n_1817)
);

BUFx8_ASAP7_75t_SL g1818 ( 
.A(n_1676),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1638),
.B(n_340),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1708),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1671),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_SL g1822 ( 
.A1(n_1670),
.A2(n_348),
.B1(n_344),
.B2(n_345),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1639),
.Y(n_1823)
);

CKINVDCx6p67_ASAP7_75t_R g1824 ( 
.A(n_1634),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1655),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1644),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1639),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1643),
.A2(n_354),
.B(n_349),
.C(n_351),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1668),
.B(n_356),
.Y(n_1829)
);

O2A1O1Ixp33_ASAP7_75t_L g1830 ( 
.A1(n_1643),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_1830)
);

NAND2x1p5_ASAP7_75t_L g1831 ( 
.A(n_1698),
.B(n_360),
.Y(n_1831)
);

A2O1A1Ixp33_ASAP7_75t_SL g1832 ( 
.A1(n_1715),
.A2(n_364),
.B(n_362),
.C(n_363),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1668),
.B(n_365),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1623),
.B(n_366),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1668),
.B(n_367),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1623),
.B(n_682),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1623),
.B(n_370),
.Y(n_1837)
);

O2A1O1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1643),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1623),
.B(n_375),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_SL g1840 ( 
.A1(n_1686),
.A2(n_376),
.B(n_377),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1623),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1623),
.B(n_681),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1655),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1668),
.B(n_378),
.Y(n_1844)
);

NOR2xp67_ASAP7_75t_L g1845 ( 
.A(n_1666),
.B(n_382),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1670),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1652),
.B(n_386),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1623),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1623),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1623),
.B(n_387),
.Y(n_1850)
);

OA21x2_ASAP7_75t_L g1851 ( 
.A1(n_1718),
.A2(n_389),
.B(n_392),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1623),
.B(n_679),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1623),
.B(n_394),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1623),
.B(n_678),
.Y(n_1854)
);

NOR3xp33_ASAP7_75t_L g1855 ( 
.A(n_1682),
.B(n_395),
.C(n_399),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1634),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1692),
.A2(n_400),
.B(n_401),
.Y(n_1857)
);

A2O1A1Ixp33_ASAP7_75t_L g1858 ( 
.A1(n_1643),
.A2(n_406),
.B(n_403),
.C(n_405),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1639),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1682),
.A2(n_407),
.B(n_408),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_SL g1861 ( 
.A1(n_1670),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_1861)
);

CKINVDCx20_ASAP7_75t_R g1862 ( 
.A(n_1644),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1623),
.B(n_412),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1623),
.Y(n_1864)
);

O2A1O1Ixp5_ASAP7_75t_SL g1865 ( 
.A1(n_1682),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_1865)
);

AOI21x1_ASAP7_75t_SL g1866 ( 
.A1(n_1717),
.A2(n_418),
.B(n_419),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1740),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1825),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1841),
.Y(n_1869)
);

BUFx3_ASAP7_75t_L g1870 ( 
.A(n_1794),
.Y(n_1870)
);

OAI21x1_ASAP7_75t_L g1871 ( 
.A1(n_1866),
.A2(n_1753),
.B(n_1857),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1848),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1843),
.B(n_421),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1730),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1785),
.Y(n_1875)
);

BUFx2_ASAP7_75t_L g1876 ( 
.A(n_1760),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1823),
.B(n_423),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1849),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1773),
.A2(n_427),
.B1(n_424),
.B2(n_425),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1864),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1734),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1799),
.B(n_428),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1822),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1743),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1748),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1741),
.Y(n_1886)
);

AO21x2_ASAP7_75t_L g1887 ( 
.A1(n_1729),
.A2(n_432),
.B(n_433),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1827),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1751),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1859),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1786),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_1725),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1727),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1783),
.Y(n_1894)
);

INVx3_ASAP7_75t_L g1895 ( 
.A(n_1754),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1779),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1781),
.B(n_434),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1747),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1797),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1726),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1742),
.Y(n_1901)
);

AOI21x1_ASAP7_75t_L g1902 ( 
.A1(n_1742),
.A2(n_435),
.B(n_439),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1800),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1806),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1771),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1774),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1731),
.B(n_440),
.Y(n_1907)
);

INVx1_ASAP7_75t_SL g1908 ( 
.A(n_1724),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1733),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1736),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1834),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1805),
.Y(n_1912)
);

OAI21x1_ASAP7_75t_L g1913 ( 
.A1(n_1768),
.A2(n_441),
.B(n_442),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1737),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1756),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1815),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1851),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1861),
.A2(n_1763),
.B1(n_1855),
.B2(n_1784),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1826),
.B(n_443),
.Y(n_1919)
);

AO21x1_ASAP7_75t_SL g1920 ( 
.A1(n_1820),
.A2(n_444),
.B(n_445),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1746),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1824),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1752),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1851),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1755),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1804),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1759),
.B(n_446),
.Y(n_1927)
);

BUFx4f_ASAP7_75t_SL g1928 ( 
.A(n_1862),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1850),
.Y(n_1929)
);

BUFx2_ASAP7_75t_L g1930 ( 
.A(n_1735),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1782),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1775),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1732),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1850),
.B(n_447),
.Y(n_1934)
);

NAND2x1p5_ASAP7_75t_L g1935 ( 
.A(n_1854),
.B(n_450),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1758),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1854),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1757),
.B(n_451),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1836),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1837),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1839),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1842),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1852),
.Y(n_1943)
);

BUFx6f_ASAP7_75t_L g1944 ( 
.A(n_1818),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1856),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1792),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1853),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1738),
.B(n_453),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1863),
.B(n_454),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1796),
.A2(n_456),
.B(n_457),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1750),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1745),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1795),
.B(n_1829),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1764),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1816),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1833),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1835),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1881),
.B(n_1769),
.Y(n_1958)
);

INVxp67_ASAP7_75t_SL g1959 ( 
.A(n_1876),
.Y(n_1959)
);

BUFx2_ASAP7_75t_L g1960 ( 
.A(n_1955),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1868),
.B(n_1739),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1895),
.B(n_1772),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1900),
.B(n_1790),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1944),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1874),
.B(n_1798),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1933),
.A2(n_1813),
.B1(n_1860),
.B2(n_1847),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1876),
.B(n_1767),
.Y(n_1967)
);

AOI22xp33_ASAP7_75t_L g1968 ( 
.A1(n_1918),
.A2(n_1762),
.B1(n_1846),
.B2(n_1793),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1889),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1928),
.B(n_1791),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1869),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1955),
.B(n_1816),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1944),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1872),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1904),
.B(n_1749),
.Y(n_1975)
);

OA21x2_ASAP7_75t_L g1976 ( 
.A1(n_1901),
.A2(n_1766),
.B(n_1765),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1878),
.Y(n_1977)
);

NOR2x1_ASAP7_75t_L g1978 ( 
.A(n_1930),
.B(n_1840),
.Y(n_1978)
);

HB1xp67_ASAP7_75t_L g1979 ( 
.A(n_1891),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1880),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1884),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1889),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1875),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1875),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1930),
.B(n_1819),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1951),
.A2(n_1778),
.B1(n_1801),
.B2(n_1809),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1885),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1899),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1936),
.B(n_1802),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1903),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1886),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1909),
.B(n_1788),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1893),
.B(n_1803),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1905),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1906),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1894),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1896),
.Y(n_1997)
);

BUFx2_ASAP7_75t_L g1998 ( 
.A(n_1867),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1890),
.B(n_1761),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1925),
.B(n_1844),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1916),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1888),
.Y(n_2002)
);

AO22x1_ASAP7_75t_L g2003 ( 
.A1(n_1952),
.A2(n_1792),
.B1(n_1810),
.B2(n_1830),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1917),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1926),
.B(n_1807),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1898),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1915),
.B(n_1831),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1892),
.B(n_1814),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1911),
.Y(n_2009)
);

INVx2_ASAP7_75t_SL g2010 ( 
.A(n_1912),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1924),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1910),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1914),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1940),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1912),
.B(n_1811),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1921),
.B(n_1780),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1941),
.Y(n_2017)
);

BUFx2_ASAP7_75t_L g2018 ( 
.A(n_1929),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1879),
.A2(n_1883),
.B1(n_1744),
.B2(n_1858),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1923),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1932),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1931),
.B(n_1817),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1956),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1957),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1942),
.Y(n_2025)
);

BUFx4f_ASAP7_75t_L g2026 ( 
.A(n_1945),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1954),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1939),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1902),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1937),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1953),
.B(n_1728),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1870),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1902),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1943),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1947),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1922),
.B(n_1845),
.Y(n_2036)
);

BUFx12f_ASAP7_75t_L g2037 ( 
.A(n_1948),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1871),
.Y(n_2038)
);

OAI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1950),
.A2(n_1828),
.B1(n_1787),
.B2(n_1838),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1908),
.B(n_1777),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1873),
.Y(n_2041)
);

AOI22xp5_ASAP7_75t_L g2042 ( 
.A1(n_1907),
.A2(n_1946),
.B1(n_1882),
.B2(n_1934),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2027),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1971),
.Y(n_2044)
);

INVx4_ASAP7_75t_L g2045 ( 
.A(n_1973),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1974),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_2032),
.B(n_1938),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1977),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1960),
.Y(n_2049)
);

INVxp67_ASAP7_75t_SL g2050 ( 
.A(n_2004),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1998),
.B(n_1919),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1972),
.B(n_1897),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1972),
.B(n_1927),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1979),
.B(n_1887),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1980),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2041),
.B(n_1877),
.Y(n_2056)
);

INVxp67_ASAP7_75t_SL g2057 ( 
.A(n_2031),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1969),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2023),
.B(n_1913),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1961),
.B(n_1920),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1981),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1987),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_2009),
.B(n_1935),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1991),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_1993),
.B(n_1982),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2018),
.B(n_1920),
.Y(n_2066)
);

INVx3_ASAP7_75t_L g2067 ( 
.A(n_2032),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2011),
.Y(n_2068)
);

OR2x2_ASAP7_75t_L g2069 ( 
.A(n_2014),
.B(n_1949),
.Y(n_2069)
);

OAI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1966),
.A2(n_1821),
.B1(n_1789),
.B2(n_1808),
.Y(n_2070)
);

HB1xp67_ASAP7_75t_L g2071 ( 
.A(n_1959),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1996),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1994),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_2039),
.A2(n_1770),
.B1(n_1776),
.B2(n_1812),
.Y(n_2074)
);

BUFx2_ASAP7_75t_L g2075 ( 
.A(n_1978),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1997),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1958),
.B(n_1865),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1985),
.B(n_458),
.Y(n_2078)
);

INVx1_ASAP7_75t_SL g2079 ( 
.A(n_1967),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2006),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2017),
.B(n_1832),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2024),
.Y(n_2082)
);

NOR2xp67_ASAP7_75t_L g2083 ( 
.A(n_2038),
.B(n_459),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_1962),
.B(n_460),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1965),
.B(n_461),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1973),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2025),
.B(n_462),
.Y(n_2087)
);

INVx2_ASAP7_75t_SL g2088 ( 
.A(n_2026),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_1992),
.B(n_463),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1995),
.Y(n_2090)
);

BUFx3_ASAP7_75t_L g2091 ( 
.A(n_1964),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_2038),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2005),
.B(n_464),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_1999),
.B(n_465),
.Y(n_2094)
);

HB1xp67_ASAP7_75t_L g2095 ( 
.A(n_2001),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_2057),
.B(n_2012),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_2075),
.B(n_2013),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2079),
.B(n_2030),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2060),
.B(n_2008),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2043),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2066),
.B(n_2010),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2077),
.B(n_1989),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2076),
.Y(n_2103)
);

INVxp67_ASAP7_75t_L g2104 ( 
.A(n_2075),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2049),
.B(n_1963),
.Y(n_2105)
);

AND2x2_ASAP7_75t_L g2106 ( 
.A(n_2052),
.B(n_2007),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2080),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2052),
.B(n_2036),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_2071),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2053),
.B(n_1984),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2090),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2082),
.B(n_2021),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_2092),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2092),
.Y(n_2114)
);

AND2x4_ASAP7_75t_SL g2115 ( 
.A(n_2045),
.B(n_1973),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_2067),
.B(n_2020),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2070),
.A2(n_2019),
.B1(n_1968),
.B2(n_1976),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2065),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2081),
.B(n_2050),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2059),
.B(n_2054),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2044),
.Y(n_2121)
);

INVx2_ASAP7_75t_SL g2122 ( 
.A(n_2086),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2046),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2051),
.B(n_2022),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_2088),
.B(n_2032),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2056),
.B(n_1983),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2073),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2058),
.B(n_2034),
.Y(n_2128)
);

AND2x4_ASAP7_75t_L g2129 ( 
.A(n_2048),
.B(n_2035),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2068),
.Y(n_2130)
);

BUFx2_ASAP7_75t_L g2131 ( 
.A(n_2091),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2055),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2061),
.Y(n_2133)
);

NAND2x1p5_ASAP7_75t_L g2134 ( 
.A(n_2083),
.B(n_2040),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_2063),
.Y(n_2135)
);

INVxp67_ASAP7_75t_SL g2136 ( 
.A(n_2095),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2062),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_2064),
.B(n_2016),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2069),
.B(n_2035),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2072),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2087),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_2109),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2123),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2117),
.B(n_2000),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_2115),
.Y(n_2145)
);

AOI21xp33_ASAP7_75t_L g2146 ( 
.A1(n_2102),
.A2(n_2074),
.B(n_1976),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2131),
.Y(n_2147)
);

AO21x2_ASAP7_75t_L g2148 ( 
.A1(n_2104),
.A2(n_2033),
.B(n_2029),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2108),
.B(n_2086),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2126),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2099),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2106),
.B(n_2047),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2141),
.B(n_1975),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2101),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2134),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2122),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2124),
.Y(n_2157)
);

HB1xp67_ASAP7_75t_L g2158 ( 
.A(n_2138),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2116),
.Y(n_2159)
);

INVx2_ASAP7_75t_SL g2160 ( 
.A(n_2125),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2116),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2141),
.A2(n_1986),
.B1(n_2003),
.B2(n_2094),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2123),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2132),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2119),
.B(n_2028),
.Y(n_2165)
);

INVxp67_ASAP7_75t_L g2166 ( 
.A(n_2136),
.Y(n_2166)
);

OAI33xp33_ASAP7_75t_L g2167 ( 
.A1(n_2132),
.A2(n_2033),
.A3(n_2029),
.B1(n_1990),
.B2(n_1988),
.B3(n_2002),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2140),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_2118),
.B(n_2085),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2097),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2140),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2139),
.B(n_2094),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2147),
.B(n_2135),
.Y(n_2173)
);

OR2x2_ASAP7_75t_L g2174 ( 
.A(n_2153),
.B(n_2096),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2145),
.B(n_2105),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_2145),
.B(n_2113),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2142),
.B(n_2166),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2149),
.B(n_2110),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2152),
.B(n_2098),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2143),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2143),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2150),
.Y(n_2182)
);

BUFx2_ASAP7_75t_SL g2183 ( 
.A(n_2156),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2160),
.Y(n_2184)
);

NAND2x1p5_ASAP7_75t_L g2185 ( 
.A(n_2155),
.B(n_2078),
.Y(n_2185)
);

NOR2x1p5_ASAP7_75t_L g2186 ( 
.A(n_2154),
.B(n_2037),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2151),
.B(n_2157),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2159),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2161),
.B(n_2170),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_2144),
.B(n_2112),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2158),
.B(n_2127),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2165),
.B(n_2130),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_2172),
.B(n_2100),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2146),
.B(n_2162),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2182),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_2178),
.B(n_2164),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2180),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2183),
.B(n_2171),
.Y(n_2198)
);

OR2x2_ASAP7_75t_L g2199 ( 
.A(n_2177),
.B(n_2169),
.Y(n_2199)
);

INVx4_ASAP7_75t_L g2200 ( 
.A(n_2176),
.Y(n_2200)
);

AND2x4_ASAP7_75t_L g2201 ( 
.A(n_2186),
.B(n_2097),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2181),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_2184),
.B(n_2167),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2175),
.B(n_2137),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2183),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2191),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_2173),
.B(n_2103),
.Y(n_2207)
);

HB1xp67_ASAP7_75t_L g2208 ( 
.A(n_2176),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2174),
.B(n_2120),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2192),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2189),
.B(n_2190),
.Y(n_2211)
);

NOR3xp33_ASAP7_75t_L g2212 ( 
.A(n_2195),
.B(n_2194),
.C(n_2188),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2208),
.B(n_2193),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2200),
.B(n_2179),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2205),
.B(n_2187),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2206),
.B(n_2163),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2210),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2196),
.B(n_2163),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2197),
.Y(n_2219)
);

INVx1_ASAP7_75t_SL g2220 ( 
.A(n_2201),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2196),
.B(n_2168),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_2211),
.B(n_2185),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_SL g2223 ( 
.A1(n_2203),
.A2(n_2168),
.B1(n_2003),
.B2(n_2114),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2204),
.B(n_2107),
.Y(n_2224)
);

AND2x2_ASAP7_75t_L g2225 ( 
.A(n_2199),
.B(n_2209),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2207),
.B(n_2111),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2214),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2225),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2220),
.B(n_2212),
.Y(n_2229)
);

INVxp67_ASAP7_75t_L g2230 ( 
.A(n_2215),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2218),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2213),
.B(n_2198),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2222),
.B(n_2202),
.Y(n_2233)
);

INVx1_ASAP7_75t_SL g2234 ( 
.A(n_2223),
.Y(n_2234)
);

INVxp67_ASAP7_75t_SL g2235 ( 
.A(n_2221),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2217),
.Y(n_2236)
);

NAND2x1p5_ASAP7_75t_L g2237 ( 
.A(n_2219),
.B(n_2093),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2226),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2224),
.B(n_2148),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_2216),
.B(n_2133),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2228),
.Y(n_2241)
);

NAND2x1_ASAP7_75t_L g2242 ( 
.A(n_2227),
.B(n_2121),
.Y(n_2242)
);

INVxp67_ASAP7_75t_L g2243 ( 
.A(n_2229),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2238),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2235),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2236),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2234),
.B(n_2129),
.Y(n_2247)
);

AOI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2232),
.A2(n_2015),
.B1(n_1970),
.B2(n_2129),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2231),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2233),
.B(n_2128),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2230),
.B(n_2084),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2231),
.Y(n_2252)
);

OAI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2237),
.A2(n_2042),
.B1(n_2089),
.B2(n_469),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2247),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2250),
.B(n_2240),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2241),
.B(n_2239),
.Y(n_2256)
);

NOR2xp67_ASAP7_75t_L g2257 ( 
.A(n_2243),
.B(n_466),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_2245),
.B(n_467),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2244),
.B(n_470),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2251),
.B(n_471),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2246),
.B(n_473),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_2242),
.B(n_474),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2249),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2252),
.B(n_475),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2248),
.B(n_476),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2253),
.B(n_478),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_2250),
.B(n_480),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2250),
.B(n_481),
.Y(n_2268)
);

INVx2_ASAP7_75t_L g2269 ( 
.A(n_2260),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2255),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2254),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2256),
.Y(n_2272)
);

XOR2x2_ASAP7_75t_L g2273 ( 
.A(n_2257),
.B(n_482),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2258),
.B(n_483),
.Y(n_2274)
);

CKINVDCx5p33_ASAP7_75t_R g2275 ( 
.A(n_2267),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2266),
.B(n_484),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2262),
.B(n_485),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2268),
.B(n_486),
.Y(n_2278)
);

NOR2xp33_ASAP7_75t_R g2279 ( 
.A(n_2263),
.B(n_677),
.Y(n_2279)
);

AO22x2_ASAP7_75t_L g2280 ( 
.A1(n_2270),
.A2(n_2264),
.B1(n_2259),
.B2(n_2261),
.Y(n_2280)
);

AOI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2269),
.A2(n_2265),
.B1(n_489),
.B2(n_487),
.Y(n_2281)
);

NAND2xp33_ASAP7_75t_L g2282 ( 
.A(n_2279),
.B(n_488),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2276),
.B(n_493),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_2271),
.B(n_494),
.Y(n_2284)
);

BUFx2_ASAP7_75t_L g2285 ( 
.A(n_2273),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2275),
.B(n_495),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2272),
.B(n_496),
.Y(n_2287)
);

OAI211xp5_ASAP7_75t_L g2288 ( 
.A1(n_2278),
.A2(n_500),
.B(n_497),
.C(n_499),
.Y(n_2288)
);

AOI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_2282),
.A2(n_2277),
.B(n_2274),
.Y(n_2289)
);

NOR2xp33_ASAP7_75t_L g2290 ( 
.A(n_2285),
.B(n_501),
.Y(n_2290)
);

NAND4xp25_ASAP7_75t_L g2291 ( 
.A(n_2281),
.B(n_509),
.C(n_506),
.D(n_508),
.Y(n_2291)
);

AOI221xp5_ASAP7_75t_L g2292 ( 
.A1(n_2280),
.A2(n_510),
.B1(n_512),
.B2(n_513),
.C(n_514),
.Y(n_2292)
);

NOR3xp33_ASAP7_75t_L g2293 ( 
.A(n_2286),
.B(n_2283),
.C(n_2287),
.Y(n_2293)
);

OA22x2_ASAP7_75t_SL g2294 ( 
.A1(n_2280),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_2288),
.B(n_519),
.Y(n_2295)
);

NAND3xp33_ASAP7_75t_L g2296 ( 
.A(n_2284),
.B(n_520),
.C(n_521),
.Y(n_2296)
);

NOR2x1_ASAP7_75t_L g2297 ( 
.A(n_2282),
.B(n_523),
.Y(n_2297)
);

AOI221xp5_ASAP7_75t_L g2298 ( 
.A1(n_2285),
.A2(n_524),
.B1(n_525),
.B2(n_526),
.C(n_527),
.Y(n_2298)
);

A2O1A1Ixp33_ASAP7_75t_L g2299 ( 
.A1(n_2281),
.A2(n_530),
.B(n_528),
.C(n_529),
.Y(n_2299)
);

NOR4xp25_ASAP7_75t_L g2300 ( 
.A(n_2282),
.B(n_533),
.C(n_531),
.D(n_532),
.Y(n_2300)
);

NOR3xp33_ASAP7_75t_L g2301 ( 
.A(n_2285),
.B(n_534),
.C(n_535),
.Y(n_2301)
);

NAND3x1_ASAP7_75t_SL g2302 ( 
.A(n_2297),
.B(n_537),
.C(n_538),
.Y(n_2302)
);

AOI32xp33_ASAP7_75t_L g2303 ( 
.A1(n_2290),
.A2(n_540),
.A3(n_541),
.B1(n_542),
.B2(n_543),
.Y(n_2303)
);

INVxp67_ASAP7_75t_L g2304 ( 
.A(n_2295),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2293),
.Y(n_2305)
);

OAI21xp5_ASAP7_75t_SL g2306 ( 
.A1(n_2289),
.A2(n_545),
.B(n_546),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2296),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2300),
.B(n_548),
.Y(n_2308)
);

OAI21xp33_ASAP7_75t_SL g2309 ( 
.A1(n_2292),
.A2(n_549),
.B(n_550),
.Y(n_2309)
);

AOI221xp5_ASAP7_75t_L g2310 ( 
.A1(n_2301),
.A2(n_551),
.B1(n_552),
.B2(n_553),
.C(n_554),
.Y(n_2310)
);

NOR2x1_ASAP7_75t_L g2311 ( 
.A(n_2291),
.B(n_558),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_2299),
.B(n_676),
.Y(n_2312)
);

NOR2x1_ASAP7_75t_L g2313 ( 
.A(n_2294),
.B(n_559),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2298),
.Y(n_2314)
);

AOI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2290),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_2297),
.Y(n_2316)
);

NOR2x1_ASAP7_75t_L g2317 ( 
.A(n_2313),
.B(n_564),
.Y(n_2317)
);

NAND3xp33_ASAP7_75t_L g2318 ( 
.A(n_2316),
.B(n_565),
.C(n_566),
.Y(n_2318)
);

NOR2x1_ASAP7_75t_L g2319 ( 
.A(n_2306),
.B(n_674),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2312),
.B(n_567),
.Y(n_2320)
);

NOR2x1_ASAP7_75t_L g2321 ( 
.A(n_2308),
.B(n_671),
.Y(n_2321)
);

NOR3x2_ASAP7_75t_L g2322 ( 
.A(n_2302),
.B(n_568),
.C(n_569),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_2304),
.B(n_570),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2311),
.B(n_571),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2309),
.B(n_572),
.Y(n_2325)
);

OAI21xp33_ASAP7_75t_L g2326 ( 
.A1(n_2305),
.A2(n_573),
.B(n_574),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2314),
.B(n_576),
.Y(n_2327)
);

NAND2xp33_ASAP7_75t_SL g2328 ( 
.A(n_2307),
.B(n_577),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2310),
.B(n_578),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2315),
.Y(n_2330)
);

NAND3xp33_ASAP7_75t_SL g2331 ( 
.A(n_2303),
.B(n_579),
.C(n_580),
.Y(n_2331)
);

NOR3x1_ASAP7_75t_L g2332 ( 
.A(n_2306),
.B(n_582),
.C(n_583),
.Y(n_2332)
);

NOR3x2_ASAP7_75t_L g2333 ( 
.A(n_2302),
.B(n_584),
.C(n_585),
.Y(n_2333)
);

NOR3xp33_ASAP7_75t_L g2334 ( 
.A(n_2305),
.B(n_587),
.C(n_589),
.Y(n_2334)
);

NOR2xp67_ASAP7_75t_L g2335 ( 
.A(n_2316),
.B(n_590),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2313),
.B(n_591),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2335),
.B(n_592),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2322),
.Y(n_2338)
);

NAND3x1_ASAP7_75t_L g2339 ( 
.A(n_2317),
.B(n_594),
.C(n_595),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2336),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2333),
.Y(n_2341)
);

INVx1_ASAP7_75t_SL g2342 ( 
.A(n_2328),
.Y(n_2342)
);

INVxp67_ASAP7_75t_L g2343 ( 
.A(n_2325),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2324),
.B(n_596),
.Y(n_2344)
);

NAND2x1p5_ASAP7_75t_L g2345 ( 
.A(n_2321),
.B(n_597),
.Y(n_2345)
);

NOR3xp33_ASAP7_75t_L g2346 ( 
.A(n_2323),
.B(n_598),
.C(n_599),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2320),
.Y(n_2347)
);

AND4x1_ASAP7_75t_L g2348 ( 
.A(n_2332),
.B(n_600),
.C(n_601),
.D(n_603),
.Y(n_2348)
);

INVxp33_ASAP7_75t_SL g2349 ( 
.A(n_2327),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2338),
.B(n_2319),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2342),
.A2(n_2331),
.B1(n_2330),
.B2(n_2329),
.Y(n_2351)
);

NAND2x1_ASAP7_75t_L g2352 ( 
.A(n_2341),
.B(n_2318),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2344),
.B(n_2348),
.Y(n_2353)
);

NAND4xp75_ASAP7_75t_L g2354 ( 
.A(n_2340),
.B(n_2334),
.C(n_2326),
.D(n_606),
.Y(n_2354)
);

OR3x2_ASAP7_75t_L g2355 ( 
.A(n_2347),
.B(n_604),
.C(n_605),
.Y(n_2355)
);

NOR2xp33_ASAP7_75t_L g2356 ( 
.A(n_2343),
.B(n_607),
.Y(n_2356)
);

AOI22xp5_ASAP7_75t_L g2357 ( 
.A1(n_2349),
.A2(n_608),
.B1(n_609),
.B2(n_610),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2345),
.Y(n_2358)
);

AND2x2_ASAP7_75t_SL g2359 ( 
.A(n_2350),
.B(n_2337),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2353),
.Y(n_2360)
);

O2A1O1Ixp33_ASAP7_75t_L g2361 ( 
.A1(n_2352),
.A2(n_2346),
.B(n_2339),
.C(n_613),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2356),
.B(n_2358),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2361),
.Y(n_2363)
);

AOI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2360),
.A2(n_2355),
.B1(n_2351),
.B2(n_2354),
.Y(n_2364)
);

A2O1A1Ixp33_ASAP7_75t_L g2365 ( 
.A1(n_2362),
.A2(n_2357),
.B(n_612),
.C(n_614),
.Y(n_2365)
);

AOI22xp33_ASAP7_75t_L g2366 ( 
.A1(n_2363),
.A2(n_2359),
.B1(n_615),
.B2(n_616),
.Y(n_2366)
);

XNOR2xp5_ASAP7_75t_L g2367 ( 
.A(n_2364),
.B(n_611),
.Y(n_2367)
);

OAI22xp5_ASAP7_75t_L g2368 ( 
.A1(n_2366),
.A2(n_2367),
.B1(n_2365),
.B2(n_619),
.Y(n_2368)
);

OAI21xp33_ASAP7_75t_L g2369 ( 
.A1(n_2367),
.A2(n_617),
.B(n_618),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2368),
.Y(n_2370)
);

NOR4xp25_ASAP7_75t_L g2371 ( 
.A(n_2369),
.B(n_620),
.C(n_621),
.D(n_622),
.Y(n_2371)
);

AOI22xp33_ASAP7_75t_R g2372 ( 
.A1(n_2370),
.A2(n_623),
.B1(n_624),
.B2(n_625),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2371),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2373),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2372),
.Y(n_2375)
);

NAND3xp33_ASAP7_75t_L g2376 ( 
.A(n_2374),
.B(n_626),
.C(n_628),
.Y(n_2376)
);

AOI21xp33_ASAP7_75t_L g2377 ( 
.A1(n_2375),
.A2(n_631),
.B(n_632),
.Y(n_2377)
);

AOI21xp33_ASAP7_75t_L g2378 ( 
.A1(n_2374),
.A2(n_633),
.B(n_634),
.Y(n_2378)
);

OA21x2_ASAP7_75t_L g2379 ( 
.A1(n_2374),
.A2(n_635),
.B(n_636),
.Y(n_2379)
);

INVxp67_ASAP7_75t_L g2380 ( 
.A(n_2379),
.Y(n_2380)
);

BUFx2_ASAP7_75t_SL g2381 ( 
.A(n_2377),
.Y(n_2381)
);

INVxp67_ASAP7_75t_SL g2382 ( 
.A(n_2376),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_2378),
.Y(n_2383)
);

OA21x2_ASAP7_75t_L g2384 ( 
.A1(n_2380),
.A2(n_637),
.B(n_638),
.Y(n_2384)
);

OR2x6_ASAP7_75t_L g2385 ( 
.A(n_2381),
.B(n_639),
.Y(n_2385)
);

OR2x6_ASAP7_75t_L g2386 ( 
.A(n_2383),
.B(n_640),
.Y(n_2386)
);

AOI21xp5_ASAP7_75t_L g2387 ( 
.A1(n_2385),
.A2(n_2382),
.B(n_641),
.Y(n_2387)
);

AOI211xp5_ASAP7_75t_L g2388 ( 
.A1(n_2387),
.A2(n_2384),
.B(n_2386),
.C(n_643),
.Y(n_2388)
);


endmodule