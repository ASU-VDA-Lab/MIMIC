module fake_jpeg_12620_n_268 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_268);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_268;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_20),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_20),
.CON(n_65),
.SN(n_65)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_21),
.B1(n_34),
.B2(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_53),
.B1(n_56),
.B2(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_52),
.Y(n_78)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_18),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_17),
.B1(n_24),
.B2(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_28),
.B1(n_24),
.B2(n_23),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_70),
.B1(n_41),
.B2(n_44),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_55),
.A2(n_60),
.B1(n_67),
.B2(n_42),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_30),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_27),
.B1(n_26),
.B2(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_20),
.B1(n_33),
.B2(n_19),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_42),
.B1(n_37),
.B2(n_3),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_65),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_45),
.B1(n_44),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_35),
.B1(n_32),
.B2(n_20),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_74),
.Y(n_131)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_46),
.C(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_81),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_36),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_86),
.Y(n_114)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_49),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_32),
.B(n_35),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_42),
.B(n_37),
.C(n_73),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_33),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_88),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_92),
.B1(n_102),
.B2(n_64),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_32),
.B1(n_29),
.B2(n_22),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_22),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_19),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_61),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_50),
.B(n_1),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_4),
.Y(n_130)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_65),
.A2(n_41),
.B1(n_42),
.B2(n_37),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_104),
.B1(n_68),
.B2(n_61),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_56),
.A2(n_42),
.B1(n_37),
.B2(n_3),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_71),
.B1(n_51),
.B2(n_68),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_105),
.A2(n_75),
.B1(n_79),
.B2(n_101),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_109),
.A2(n_112),
.B1(n_90),
.B2(n_5),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_128),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_93),
.A2(n_84),
.B1(n_103),
.B2(n_80),
.Y(n_112)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_96),
.Y(n_136)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_118),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_2),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_87),
.Y(n_132)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_126),
.B1(n_93),
.B2(n_74),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_68),
.B1(n_61),
.B2(n_37),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_78),
.B(n_4),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_130),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_120),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_134),
.A2(n_144),
.B1(n_154),
.B2(n_125),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_81),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_135),
.B(n_147),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_136),
.A2(n_158),
.B(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_83),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_143),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_76),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_97),
.B1(n_82),
.B2(n_74),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_99),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_113),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_101),
.C(n_75),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_115),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_75),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_155),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_77),
.B1(n_79),
.B2(n_91),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_85),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_156),
.A2(n_113),
.B1(n_118),
.B2(n_125),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_4),
.B(n_5),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_6),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_6),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_165),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_119),
.B(n_111),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_168),
.B(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_108),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_129),
.B(n_106),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_144),
.B1(n_146),
.B2(n_138),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_108),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_152),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_180),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_143),
.C(n_137),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_134),
.A2(n_127),
.B1(n_107),
.B2(n_8),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_127),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_9),
.B(n_10),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_135),
.B(n_133),
.Y(n_193)
);

OA21x2_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_156),
.B(n_142),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_200),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_151),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_204),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_189),
.A2(n_193),
.B1(n_185),
.B2(n_180),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_162),
.C(n_178),
.Y(n_223)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_152),
.B(n_132),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_201),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_191),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_SL g204 ( 
.A(n_163),
.B(n_133),
.C(n_159),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_145),
.C(n_140),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_206),
.C(n_164),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_139),
.C(n_148),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_211),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_181),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_193),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_175),
.B1(n_174),
.B2(n_183),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_212),
.A2(n_222),
.B1(n_197),
.B2(n_202),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_218),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_182),
.B1(n_169),
.B2(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_164),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_175),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_223),
.C(n_206),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_171),
.B(n_168),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_197),
.B1(n_202),
.B2(n_194),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_186),
.A2(n_181),
.B1(n_173),
.B2(n_169),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_219),
.C(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_215),
.Y(n_238)
);

NAND4xp25_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_233),
.C(n_226),
.D(n_236),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_192),
.A3(n_204),
.B1(n_201),
.B2(n_190),
.C1(n_200),
.C2(n_195),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_232),
.Y(n_240)
);

AO221x1_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_187),
.B1(n_201),
.B2(n_157),
.C(n_146),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_189),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_157),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_222),
.B1(n_207),
.B2(n_220),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_218),
.B1(n_211),
.B2(n_213),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_241),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_187),
.C(n_208),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_166),
.C(n_10),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_246),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_234),
.B(n_232),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_249),
.B(n_242),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_234),
.B(n_233),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_228),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_248),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_254),
.A2(n_256),
.B(n_257),
.Y(n_261)
);

OAI211xp5_ASAP7_75t_L g255 ( 
.A1(n_253),
.A2(n_245),
.B(n_244),
.C(n_243),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_255),
.A2(n_258),
.B(n_250),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_247),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

NOR4xp25_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_9),
.C(n_11),
.D(n_12),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_257),
.A2(n_237),
.B(n_235),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_260),
.B(n_262),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_257),
.A2(n_231),
.B(n_11),
.Y(n_262)
);

NOR4xp25_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_261),
.C(n_13),
.D(n_14),
.Y(n_265)
);

OAI21xp33_ASAP7_75t_L g266 ( 
.A1(n_265),
.A2(n_12),
.B(n_13),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g267 ( 
.A(n_266),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_264),
.Y(n_268)
);


endmodule