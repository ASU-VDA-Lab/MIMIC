module real_aes_8025_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_792;
wire n_673;
wire n_386;
wire n_503;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_852;
wire n_857;
wire n_461;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_397;
wire n_275;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_691;
wire n_765;
wire n_498;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_0), .A2(n_240), .B1(n_440), .B2(n_540), .Y(n_539) );
AOI22xp33_ASAP7_75t_SL g541 ( .A1(n_1), .A2(n_111), .B1(n_432), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_2), .A2(n_252), .B1(n_451), .B2(n_454), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_3), .A2(n_251), .B1(n_300), .B2(n_479), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_4), .A2(n_41), .B1(n_284), .B2(n_300), .C(n_305), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_5), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_6), .B(n_344), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_7), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_8), .A2(n_259), .B1(n_339), .B2(n_673), .Y(n_863) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_9), .A2(n_99), .B1(n_482), .B2(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_10), .A2(n_162), .B1(n_405), .B2(n_476), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_11), .B(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_12), .A2(n_73), .B1(n_479), .B2(n_481), .Y(n_478) );
XOR2x2_ASAP7_75t_L g591 ( .A(n_13), .B(n_592), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_14), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_15), .A2(n_175), .B1(n_308), .B2(n_482), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_16), .Y(n_821) );
AOI22xp33_ASAP7_75t_SL g632 ( .A1(n_17), .A2(n_119), .B1(n_476), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_18), .A2(n_214), .B1(n_408), .B2(n_547), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_19), .A2(n_215), .B1(n_339), .B2(n_343), .C(n_345), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_20), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_21), .A2(n_134), .B1(n_628), .B2(n_635), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_22), .A2(n_157), .B1(n_860), .B2(n_861), .Y(n_859) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_23), .A2(n_183), .B1(n_628), .B2(n_629), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_24), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_25), .A2(n_33), .B1(n_396), .B2(n_454), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_26), .A2(n_470), .B1(n_512), .B2(n_513), .Y(n_469) );
INVx1_ASAP7_75t_L g513 ( .A(n_26), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_27), .A2(n_260), .B1(n_454), .B2(n_531), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_28), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_29), .A2(n_38), .B1(n_438), .B2(n_786), .Y(n_836) );
AO22x2_ASAP7_75t_L g297 ( .A1(n_30), .A2(n_84), .B1(n_289), .B2(n_294), .Y(n_297) );
INVx1_ASAP7_75t_L g810 ( .A(n_30), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_31), .A2(n_46), .B1(n_571), .B2(n_573), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_32), .A2(n_39), .B1(n_396), .B2(n_620), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_34), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_35), .B(n_673), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_36), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_37), .A2(n_49), .B1(n_431), .B2(n_835), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_40), .A2(n_77), .B1(n_489), .B2(n_491), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_42), .A2(n_163), .B1(n_370), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_43), .A2(n_59), .B1(n_776), .B2(n_777), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_44), .A2(n_262), .B1(n_452), .B2(n_500), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_45), .A2(n_237), .B1(n_324), .B2(n_832), .Y(n_831) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_47), .A2(n_86), .B1(n_289), .B2(n_290), .Y(n_299) );
INVx1_ASAP7_75t_L g811 ( .A(n_47), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_48), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_50), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_51), .A2(n_185), .B1(n_551), .B2(n_737), .Y(n_736) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_52), .A2(n_100), .B1(n_491), .B2(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_53), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_54), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_55), .A2(n_269), .B1(n_324), .B2(n_552), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_56), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_57), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_58), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_60), .A2(n_246), .B1(n_531), .B2(n_776), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_61), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_62), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_63), .A2(n_194), .B1(n_440), .B2(n_442), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_64), .A2(n_241), .B1(n_284), .B2(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_65), .A2(n_187), .B1(n_441), .B2(n_629), .Y(n_760) );
AOI222xp33_ASAP7_75t_L g359 ( .A1(n_66), .A2(n_90), .B1(n_146), .B2(n_360), .C1(n_363), .C2(n_369), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_67), .A2(n_144), .B1(n_395), .B2(n_451), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_68), .B(n_340), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_69), .Y(n_398) );
INVx1_ASAP7_75t_L g608 ( .A(n_70), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_71), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_72), .A2(n_122), .B1(n_319), .B2(n_324), .C(n_328), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_74), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_75), .A2(n_155), .B1(n_302), .B2(n_635), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_76), .A2(n_255), .B1(n_371), .B2(n_526), .Y(n_609) );
AOI22xp33_ASAP7_75t_SL g654 ( .A1(n_78), .A2(n_239), .B1(n_489), .B2(n_655), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g346 ( .A(n_79), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_80), .A2(n_141), .B1(n_430), .B2(n_432), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_81), .A2(n_203), .B1(n_455), .B2(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g575 ( .A1(n_82), .A2(n_139), .B1(n_413), .B2(n_576), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_83), .A2(n_123), .B1(n_324), .B2(n_438), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_85), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_87), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g732 ( .A1(n_88), .A2(n_174), .B1(n_479), .B2(n_569), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_89), .Y(n_849) );
INVx1_ASAP7_75t_L g278 ( .A(n_91), .Y(n_278) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_92), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g684 ( .A1(n_93), .A2(n_153), .B1(n_573), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_94), .A2(n_192), .B1(n_395), .B2(n_396), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_95), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_96), .A2(n_182), .B1(n_302), .B2(n_635), .Y(n_749) );
INVx1_ASAP7_75t_L g274 ( .A(n_97), .Y(n_274) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_98), .A2(n_222), .B1(n_451), .B2(n_526), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_101), .A2(n_235), .B1(n_598), .B2(n_691), .Y(n_869) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_102), .A2(n_231), .B1(n_413), .B2(n_416), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_103), .A2(n_113), .B1(n_416), .B2(n_438), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_104), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_105), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_106), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_107), .A2(n_229), .B1(n_482), .B2(n_573), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_108), .A2(n_206), .B1(n_308), .B2(n_319), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_109), .A2(n_814), .B1(n_837), .B2(n_838), .Y(n_813) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_109), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_110), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_112), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_114), .A2(n_129), .B1(n_452), .B2(n_526), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_115), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_116), .A2(n_208), .B1(n_435), .B2(n_571), .Y(n_784) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_117), .A2(n_230), .B1(n_284), .B2(n_302), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g865 ( .A1(n_118), .A2(n_210), .B1(n_324), .B2(n_866), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_120), .B(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_121), .A2(n_213), .B1(n_310), .B2(n_544), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_124), .A2(n_258), .B1(n_371), .B2(n_620), .Y(n_822) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_125), .A2(n_158), .B1(n_405), .B2(n_408), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_126), .A2(n_199), .B1(n_365), .B2(n_530), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_127), .Y(n_351) );
XOR2x2_ASAP7_75t_L g714 ( .A(n_128), .B(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_130), .A2(n_211), .B1(n_549), .B2(n_551), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_131), .Y(n_534) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_132), .A2(n_154), .B1(n_691), .B2(n_692), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_133), .A2(n_169), .B1(n_435), .B2(n_437), .Y(n_434) );
AND2x2_ASAP7_75t_L g277 ( .A(n_135), .B(n_278), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_136), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_137), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_138), .A2(n_145), .B1(n_416), .B2(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_140), .A2(n_228), .B1(n_540), .B2(n_598), .Y(n_659) );
INVx1_ASAP7_75t_L g636 ( .A(n_142), .Y(n_636) );
OA22x2_ASAP7_75t_L g667 ( .A1(n_143), .A2(n_668), .B1(n_669), .B2(n_694), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_143), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_147), .B(n_344), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_148), .B(n_602), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_149), .A2(n_263), .B1(n_734), .B2(n_786), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g867 ( .A1(n_150), .A2(n_166), .B1(n_432), .B2(n_542), .Y(n_867) );
AND2x6_ASAP7_75t_L g273 ( .A(n_151), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_151), .Y(n_804) );
AO22x2_ASAP7_75t_L g288 ( .A1(n_152), .A2(n_221), .B1(n_289), .B2(n_290), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_156), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_159), .A2(n_253), .B1(n_454), .B2(n_531), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_160), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_161), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_164), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_165), .A2(n_207), .B1(n_366), .B2(n_452), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_167), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_168), .B(n_562), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_170), .Y(n_646) );
XNOR2x1_ASAP7_75t_L g553 ( .A(n_171), .B(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_172), .A2(n_268), .B1(n_343), .B2(n_602), .Y(n_601) );
AO22x2_ASAP7_75t_L g293 ( .A1(n_173), .A2(n_242), .B1(n_289), .B2(n_294), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_176), .A2(n_265), .B1(n_413), .B2(n_441), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_177), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_178), .A2(n_423), .B1(n_465), .B2(n_466), .Y(n_422) );
INVx1_ASAP7_75t_L g465 ( .A(n_178), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_179), .A2(n_218), .B1(n_441), .B2(n_547), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_180), .A2(n_254), .B1(n_416), .B2(n_431), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_181), .Y(n_817) );
AOI22xp5_ASAP7_75t_SL g379 ( .A1(n_184), .A2(n_380), .B1(n_417), .B2(n_418), .Y(n_379) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_184), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_186), .A2(n_209), .B1(n_687), .B2(n_688), .Y(n_686) );
XNOR2x1_ASAP7_75t_L g637 ( .A(n_188), .B(n_638), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_189), .Y(n_505) );
AO22x1_ASAP7_75t_L g281 ( .A1(n_190), .A2(n_282), .B1(n_373), .B2(n_374), .Y(n_281) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_190), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_191), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_193), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_195), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_196), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_197), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_198), .A2(n_264), .B1(n_476), .B2(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_200), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_201), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_202), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_204), .B(n_344), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_205), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_212), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_216), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_217), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_219), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_220), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_221), .B(n_809), .Y(n_808) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_223), .A2(n_271), .B(n_279), .C(n_812), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_224), .Y(n_329) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_225), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_226), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_227), .Y(n_428) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_232), .A2(n_236), .B1(n_628), .B2(n_658), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_233), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g759 ( .A1(n_234), .A2(n_266), .B1(n_321), .B2(n_406), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_238), .Y(n_497) );
INVx1_ASAP7_75t_L g807 ( .A(n_242), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_243), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_244), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_245), .B(n_365), .Y(n_725) );
OA22x2_ASAP7_75t_L g763 ( .A1(n_247), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_763) );
CKINVDCx16_ASAP7_75t_R g764 ( .A(n_247), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_248), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g870 ( .A1(n_249), .A2(n_267), .B1(n_405), .B2(n_871), .Y(n_870) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_250), .Y(n_521) );
INVx1_ASAP7_75t_L g289 ( .A(n_256), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_256), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_257), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_261), .Y(n_824) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_274), .Y(n_803) );
OAI21xp5_ASAP7_75t_L g847 ( .A1(n_275), .A2(n_802), .B(n_848), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_585), .B1(n_797), .B2(n_798), .C(n_799), .Y(n_279) );
INVx1_ASAP7_75t_L g798 ( .A(n_280), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_375), .B1(n_583), .B2(n_584), .Y(n_280) );
INVx1_ASAP7_75t_L g583 ( .A(n_281), .Y(n_583) );
INVx1_ASAP7_75t_L g374 ( .A(n_282), .Y(n_374) );
AND4x1_ASAP7_75t_L g282 ( .A(n_283), .B(n_318), .C(n_338), .D(n_359), .Y(n_282) );
BUFx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_285), .Y(n_441) );
INVx2_ASAP7_75t_L g572 ( .A(n_285), .Y(n_572) );
BUFx2_ASAP7_75t_SL g687 ( .A(n_285), .Y(n_687) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_295), .Y(n_285) );
AND2x4_ASAP7_75t_L g310 ( .A(n_286), .B(n_311), .Y(n_310) );
AND2x6_ASAP7_75t_L g321 ( .A(n_286), .B(n_322), .Y(n_321) );
AND2x6_ASAP7_75t_L g362 ( .A(n_286), .B(n_356), .Y(n_362) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_292), .Y(n_286) );
AND2x2_ASAP7_75t_L g304 ( .A(n_287), .B(n_293), .Y(n_304) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_288), .B(n_293), .Y(n_327) );
AND2x2_ASAP7_75t_L g349 ( .A(n_288), .B(n_297), .Y(n_349) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g294 ( .A(n_291), .Y(n_294) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g317 ( .A(n_293), .Y(n_317) );
INVx1_ASAP7_75t_L g368 ( .A(n_293), .Y(n_368) );
AND2x4_ASAP7_75t_L g303 ( .A(n_295), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_295), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g325 ( .A(n_295), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g407 ( .A(n_295), .B(n_316), .Y(n_407) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_296), .B(n_299), .Y(n_311) );
OR2x2_ASAP7_75t_L g323 ( .A(n_296), .B(n_299), .Y(n_323) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g356 ( .A(n_297), .B(n_299), .Y(n_356) );
INVx1_ASAP7_75t_L g350 ( .A(n_298), .Y(n_350) );
AND2x2_ASAP7_75t_L g367 ( .A(n_298), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g337 ( .A(n_299), .Y(n_337) );
INVx4_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx4_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx3_ASAP7_75t_L g438 ( .A(n_303), .Y(n_438) );
INVx2_ASAP7_75t_L g484 ( .A(n_303), .Y(n_484) );
BUFx3_ASAP7_75t_L g552 ( .A(n_303), .Y(n_552) );
BUFx3_ASAP7_75t_L g578 ( .A(n_303), .Y(n_578) );
AND2x4_ASAP7_75t_L g342 ( .A(n_304), .B(n_322), .Y(n_342) );
AND2x6_ASAP7_75t_L g344 ( .A(n_304), .B(n_311), .Y(n_344) );
INVx1_ASAP7_75t_L g386 ( .A(n_304), .Y(n_386) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_304), .B(n_311), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B1(n_312), .B2(n_313), .Y(n_305) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_307), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_787) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx3_ASAP7_75t_L g576 ( .A(n_309), .Y(n_576) );
INVx2_ASAP7_75t_L g691 ( .A(n_309), .Y(n_691) );
INVx2_ASAP7_75t_L g835 ( .A(n_309), .Y(n_835) );
INVx6_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g442 ( .A(n_310), .Y(n_442) );
BUFx3_ASAP7_75t_L g476 ( .A(n_310), .Y(n_476) );
BUFx3_ASAP7_75t_L g540 ( .A(n_310), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_311), .B(n_316), .Y(n_331) );
AND2x2_ASAP7_75t_L g415 ( .A(n_311), .B(n_316), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g425 ( .A1(n_313), .A2(n_426), .B1(n_427), .B2(n_428), .C(n_429), .Y(n_425) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g790 ( .A(n_314), .Y(n_790) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g358 ( .A(n_317), .Y(n_358) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx4_ASAP7_75t_L g598 ( .A(n_320), .Y(n_598) );
INVx2_ASAP7_75t_SL g737 ( .A(n_320), .Y(n_737) );
INVx11_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx11_ASAP7_75t_L g436 ( .A(n_321), .Y(n_436) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g385 ( .A(n_323), .B(n_386), .Y(n_385) );
BUFx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_SL g408 ( .A(n_325), .Y(n_408) );
INVx1_ASAP7_75t_L g486 ( .A(n_325), .Y(n_486) );
BUFx2_ASAP7_75t_SL g569 ( .A(n_325), .Y(n_569) );
BUFx3_ASAP7_75t_L g629 ( .A(n_325), .Y(n_629) );
BUFx2_ASAP7_75t_L g688 ( .A(n_325), .Y(n_688) );
AND2x2_ASAP7_75t_L g635 ( .A(n_326), .B(n_350), .Y(n_635) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x6_ASAP7_75t_L g336 ( .A(n_327), .B(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_330), .B1(n_332), .B2(n_333), .Y(n_328) );
BUFx2_ASAP7_75t_R g330 ( .A(n_331), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_334), .Y(n_333) );
BUFx4f_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g416 ( .A(n_335), .Y(n_416) );
BUFx2_ASAP7_75t_L g786 ( .A(n_335), .Y(n_786) );
INVx6_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g432 ( .A(n_336), .Y(n_432) );
INVx1_ASAP7_75t_L g491 ( .A(n_336), .Y(n_491) );
INVx1_ASAP7_75t_SL g655 ( .A(n_336), .Y(n_655) );
INVx1_ASAP7_75t_L g453 ( .A(n_337), .Y(n_453) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx5_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g562 ( .A(n_341), .Y(n_562) );
INVx2_ASAP7_75t_L g602 ( .A(n_341), .Y(n_602) );
INVx2_ASAP7_75t_L g676 ( .A(n_341), .Y(n_676) );
INVx4_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx4f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g564 ( .A(n_344), .Y(n_564) );
INVx1_ASAP7_75t_SL g674 ( .A(n_344), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_351), .B2(n_352), .Y(n_345) );
OAI22xp5_ASAP7_75t_SL g533 ( .A1(n_347), .A2(n_534), .B1(n_535), .B2(n_536), .Y(n_533) );
BUFx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx4_ASAP7_75t_L g400 ( .A(n_348), .Y(n_400) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_348), .Y(n_728) );
OAI22xp33_ASAP7_75t_SL g779 ( .A1(n_348), .A2(n_535), .B1(n_780), .B2(n_781), .Y(n_779) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x4_ASAP7_75t_L g366 ( .A(n_349), .B(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g371 ( .A(n_349), .B(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g452 ( .A(n_349), .B(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_352), .A2(n_399), .B1(n_649), .B2(n_650), .Y(n_648) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g535 ( .A(n_353), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g353 ( .A(n_354), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_398), .B1(n_399), .B2(n_401), .Y(n_397) );
BUFx2_ASAP7_75t_L g511 ( .A(n_354), .Y(n_511) );
OR2x6_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g455 ( .A(n_356), .B(n_358), .Y(n_455) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx4_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI21xp5_ASAP7_75t_SL g556 ( .A1(n_361), .A2(n_557), .B(n_558), .Y(n_556) );
BUFx2_ASAP7_75t_L g679 ( .A(n_361), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_361), .A2(n_703), .B(n_704), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g751 ( .A1(n_361), .A2(n_752), .B(n_753), .Y(n_751) );
INVx4_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g392 ( .A(n_362), .Y(n_392) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_362), .Y(n_460) );
INVx2_ASAP7_75t_L g502 ( .A(n_362), .Y(n_502) );
BUFx3_ASAP7_75t_L g607 ( .A(n_362), .Y(n_607) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx4_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g776 ( .A(n_365), .Y(n_776) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
BUFx4f_ASAP7_75t_SL g500 ( .A(n_366), .Y(n_500) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_366), .Y(n_526) );
BUFx2_ASAP7_75t_L g826 ( .A(n_366), .Y(n_826) );
INVx1_ASAP7_75t_L g372 ( .A(n_368), .Y(n_372) );
INVx2_ASAP7_75t_L g723 ( .A(n_369), .Y(n_723) );
BUFx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g463 ( .A(n_370), .Y(n_463) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx12f_ASAP7_75t_L g396 ( .A(n_371), .Y(n_396) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_371), .Y(n_531) );
INVx1_ASAP7_75t_L g584 ( .A(n_375), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_419), .B2(n_582), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g417 ( .A(n_380), .Y(n_417) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_402), .Y(n_380) );
NOR3xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_391), .C(n_397), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B1(n_387), .B2(n_388), .Y(n_382) );
OAI221xp5_ASAP7_75t_SL g444 ( .A1(n_384), .A2(n_445), .B1(n_446), .B2(n_449), .C(n_450), .Y(n_444) );
OAI22xp5_ASAP7_75t_SL g520 ( .A1(n_384), .A2(n_448), .B1(n_521), .B2(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g770 ( .A(n_384), .Y(n_770) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g496 ( .A(n_385), .Y(n_496) );
BUFx3_ASAP7_75t_L g642 ( .A(n_385), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_385), .A2(n_817), .B1(n_818), .B2(n_819), .Y(n_816) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g819 ( .A(n_389), .Y(n_819) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g448 ( .A(n_390), .Y(n_448) );
OAI21xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_393), .B(n_394), .Y(n_391) );
OAI222xp33_ASAP7_75t_L g523 ( .A1(n_392), .A2(n_524), .B1(n_527), .B2(n_528), .C1(n_529), .C2(n_532), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_395), .Y(n_457) );
BUFx4f_ASAP7_75t_SL g509 ( .A(n_396), .Y(n_509) );
INVx2_ASAP7_75t_L g778 ( .A(n_396), .Y(n_778) );
INVx3_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g504 ( .A(n_400), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_410), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_409), .Y(n_403) );
BUFx4f_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g550 ( .A(n_406), .Y(n_550) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx3_ASAP7_75t_L g482 ( .A(n_407), .Y(n_482) );
BUFx3_ASAP7_75t_L g628 ( .A(n_407), .Y(n_628) );
BUFx3_ASAP7_75t_L g685 ( .A(n_407), .Y(n_685) );
INVx1_ASAP7_75t_L g427 ( .A(n_408), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g431 ( .A(n_414), .Y(n_431) );
BUFx3_ASAP7_75t_L g490 ( .A(n_414), .Y(n_490) );
INVx4_ASAP7_75t_L g544 ( .A(n_414), .Y(n_544) );
INVx5_ASAP7_75t_L g633 ( .A(n_414), .Y(n_633) );
INVx1_ASAP7_75t_L g692 ( .A(n_414), .Y(n_692) );
INVx8_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g582 ( .A(n_419), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_467), .B2(n_581), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
AND2x2_ASAP7_75t_SL g423 ( .A(n_424), .B(n_443), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_433), .Y(n_424) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_439), .Y(n_433) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_436), .Y(n_473) );
INVx5_ASAP7_75t_SL g547 ( .A(n_436), .Y(n_547) );
INVx4_ASAP7_75t_L g573 ( .A(n_436), .Y(n_573) );
INVx2_ASAP7_75t_SL g711 ( .A(n_436), .Y(n_711) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g480 ( .A(n_441), .Y(n_480) );
BUFx6f_ASAP7_75t_L g871 ( .A(n_441), .Y(n_871) );
NOR2xp33_ASAP7_75t_SL g443 ( .A(n_444), .B(n_456), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_446), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_717) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_448), .A2(n_494), .B1(n_495), .B2(n_497), .Y(n_493) );
BUFx3_ASAP7_75t_L g644 ( .A(n_448), .Y(n_644) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx3_ASAP7_75t_L g604 ( .A(n_452), .Y(n_604) );
BUFx2_ASAP7_75t_L g860 ( .A(n_452), .Y(n_860) );
INVx1_ASAP7_75t_SL g862 ( .A(n_454), .Y(n_862) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_SL g559 ( .A(n_455), .Y(n_559) );
BUFx3_ASAP7_75t_L g620 ( .A(n_455), .Y(n_620) );
OAI222xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_459), .B2(n_461), .C1(n_462), .C2(n_464), .Y(n_456) );
INVx2_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g855 ( .A(n_460), .Y(n_855) );
INVxp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g581 ( .A(n_467), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_514), .B2(n_515), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g512 ( .A(n_470), .Y(n_512) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_471), .B(n_492), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_472), .B(n_483), .Y(n_471) );
OAI221xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_474), .B1(n_475), .B2(n_477), .C(n_478), .Y(n_472) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI221xp5_ASAP7_75t_SL g483 ( .A1(n_484), .A2(n_485), .B1(n_486), .B2(n_487), .C(n_488), .Y(n_483) );
INVx2_ASAP7_75t_L g866 ( .A(n_484), .Y(n_866) );
INVx1_ASAP7_75t_L g658 ( .A(n_486), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_486), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_791) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_498), .C(n_506), .Y(n_492) );
INVx1_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g719 ( .A(n_496), .Y(n_719) );
OAI222xp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_501), .B1(n_502), .B2(n_503), .C1(n_504), .C2(n_505), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_502), .A2(n_618), .B(n_619), .Y(n_617) );
OAI21xp33_ASAP7_75t_SL g645 ( .A1(n_502), .A2(n_646), .B(n_647), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_502), .A2(n_722), .B1(n_723), .B2(n_724), .C(n_725), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_504), .A2(n_824), .B1(n_825), .B2(n_827), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B1(n_510), .B2(n_511), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_553), .B1(n_579), .B2(n_580), .Y(n_515) );
INVx2_ASAP7_75t_L g579 ( .A(n_516), .Y(n_579) );
XNOR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_537), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_523), .C(n_533), .Y(n_519) );
INVx2_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx4f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_535), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_545), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g734 ( .A(n_544), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g580 ( .A(n_553), .Y(n_580) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_566), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_560), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .C(n_565), .Y(n_560) );
NOR2x1_ASAP7_75t_L g566 ( .A(n_567), .B(n_574), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx3_ASAP7_75t_L g832 ( .A(n_572), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx1_ASAP7_75t_L g793 ( .A(n_578), .Y(n_793) );
INVx1_ASAP7_75t_L g797 ( .A(n_585), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_660), .B2(n_796), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AO22x1_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_610), .B2(n_611), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
NOR4xp75_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .C(n_600), .D(n_605), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_597), .B(n_599), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_601), .B(n_603), .Y(n_600) );
OAI21xp5_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_608), .B(n_609), .Y(n_605) );
OAI21xp33_ASAP7_75t_SL g773 ( .A1(n_606), .A2(n_774), .B(n_775), .Y(n_773) );
OAI21xp33_ASAP7_75t_L g820 ( .A1(n_606), .A2(n_821), .B(n_822), .Y(n_820) );
INVx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
XNOR2x1_ASAP7_75t_SL g611 ( .A(n_612), .B(n_637), .Y(n_611) );
INVx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
XOR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_636), .Y(n_614) );
NAND2x1p5_ASAP7_75t_L g615 ( .A(n_616), .B(n_625), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_621), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .C(n_624), .Y(n_621) );
NOR2x1_ASAP7_75t_L g625 ( .A(n_626), .B(n_631), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_630), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
AND2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_651), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_645), .C(n_648), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B1(n_643), .B2(n_644), .Y(n_640) );
OAI22xp5_ASAP7_75t_SL g768 ( .A1(n_644), .A2(n_769), .B1(n_771), .B2(n_772), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_656), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g796 ( .A(n_660), .Y(n_796) );
XOR2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_740), .Y(n_660) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_714), .B2(n_739), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_667), .B1(n_695), .B2(n_696), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_SL g694 ( .A(n_669), .Y(n_694) );
NAND2x1p5_ASAP7_75t_L g669 ( .A(n_670), .B(n_682), .Y(n_669) );
NOR2xp67_ASAP7_75t_SL g670 ( .A(n_671), .B(n_678), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .C(n_677), .Y(n_671) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_680), .B(n_681), .Y(n_678) );
NOR2x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_689), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_695), .A2(n_741), .B1(n_742), .B2(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_695), .Y(n_741) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
XOR2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_713), .Y(n_696) );
NAND3x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .C(n_709), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
NOR2x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .C(n_708), .Y(n_705) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx2_ASAP7_75t_L g739 ( .A(n_714), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_730), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_721), .C(n_726), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_735), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_762), .B1(n_763), .B2(n_795), .Y(n_744) );
INVx3_ASAP7_75t_L g795 ( .A(n_745), .Y(n_795) );
XOR2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_761), .Y(n_745) );
NAND3x1_ASAP7_75t_SL g746 ( .A(n_747), .B(n_750), .C(n_758), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
NOR2x1_ASAP7_75t_L g750 ( .A(n_751), .B(n_754), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .C(n_757), .Y(n_754) );
AND2x2_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_782), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_773), .C(n_779), .Y(n_767) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx3_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_787), .C(n_791), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
INVx1_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
NOR2x1_ASAP7_75t_L g800 ( .A(n_801), .B(n_805), .Y(n_800) );
OR2x2_ASAP7_75t_SL g874 ( .A(n_801), .B(n_806), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_804), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_802), .Y(n_841) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_803), .B(n_845), .Y(n_848) );
CKINVDCx16_ASAP7_75t_R g845 ( .A(n_804), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
OAI322xp33_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_839), .A3(n_842), .B1(n_846), .B2(n_849), .C1(n_850), .C2(n_872), .Y(n_812) );
INVx1_ASAP7_75t_L g838 ( .A(n_814), .Y(n_838) );
AND2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_828), .Y(n_814) );
NOR3xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_820), .C(n_823), .Y(n_815) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_833), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_836), .Y(n_833) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
BUFx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
CKINVDCx16_ASAP7_75t_R g846 ( .A(n_847), .Y(n_846) );
XNOR2xp5_ASAP7_75t_L g851 ( .A(n_849), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_864), .C(n_868), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_858), .Y(n_853) );
OAI21xp5_ASAP7_75t_SL g854 ( .A1(n_855), .A2(n_856), .B(n_857), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_863), .Y(n_858) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
AND2x2_ASAP7_75t_L g864 ( .A(n_865), .B(n_867), .Y(n_864) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_873), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
endmodule