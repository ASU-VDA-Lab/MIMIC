module real_aes_7273_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_316;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g483 ( .A1(n_0), .A2(n_187), .B(n_484), .C(n_487), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_1), .B(n_478), .Y(n_489) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g121 ( .A(n_2), .Y(n_121) );
INVx1_ASAP7_75t_L g236 ( .A(n_3), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_4), .B(n_175), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_5), .A2(n_462), .B(n_532), .Y(n_531) );
OAI22xp5_ASAP7_75t_SL g759 ( .A1(n_6), .A2(n_9), .B1(n_445), .B2(n_760), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_6), .Y(n_760) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_7), .A2(n_192), .B(n_541), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_8), .A2(n_39), .B1(n_148), .B2(n_160), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_9), .A2(n_132), .B1(n_133), .B2(n_445), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_9), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_10), .B(n_192), .Y(n_225) );
AND2x6_ASAP7_75t_L g163 ( .A(n_11), .B(n_164), .Y(n_163) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_12), .A2(n_163), .B(n_465), .C(n_554), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_13), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_14), .B(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_14), .B(n_40), .Y(n_122) );
INVx1_ASAP7_75t_L g144 ( .A(n_15), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_16), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g230 ( .A(n_17), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_18), .B(n_175), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_19), .B(n_190), .Y(n_208) );
AO32x2_ASAP7_75t_L g184 ( .A1(n_20), .A2(n_185), .A3(n_189), .B1(n_191), .B2(n_192), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_21), .A2(n_100), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_21), .Y(n_127) );
AND2x2_ASAP7_75t_L g526 ( .A(n_22), .B(n_140), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_23), .B(n_148), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_24), .B(n_190), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_25), .A2(n_55), .B1(n_148), .B2(n_160), .Y(n_188) );
AOI22xp33_ASAP7_75t_SL g201 ( .A1(n_26), .A2(n_82), .B1(n_148), .B2(n_152), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_27), .B(n_148), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_28), .A2(n_191), .B(n_465), .C(n_467), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_29), .A2(n_191), .B(n_465), .C(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_30), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_31), .B(n_140), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_32), .A2(n_462), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_33), .B(n_140), .Y(n_182) );
INVx2_ASAP7_75t_L g150 ( .A(n_34), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_35), .A2(n_496), .B(n_497), .C(n_501), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_36), .B(n_148), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_37), .B(n_140), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_38), .B(n_155), .Y(n_545) );
INVx1_ASAP7_75t_L g108 ( .A(n_40), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_41), .B(n_461), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_42), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_43), .B(n_175), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_44), .B(n_462), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_45), .A2(n_496), .B(n_501), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_46), .B(n_148), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_47), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g485 ( .A(n_48), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_49), .A2(n_91), .B1(n_160), .B2(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g524 ( .A(n_50), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_51), .B(n_148), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_52), .B(n_148), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_53), .B(n_462), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_54), .B(n_223), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g212 ( .A1(n_56), .A2(n_60), .B1(n_148), .B2(n_152), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_57), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_58), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_59), .B(n_148), .Y(n_249) );
INVx1_ASAP7_75t_L g164 ( .A(n_61), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_62), .B(n_462), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_63), .B(n_478), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_64), .A2(n_223), .B(n_233), .C(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_65), .B(n_148), .Y(n_237) );
INVx1_ASAP7_75t_L g143 ( .A(n_66), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_67), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_68), .B(n_175), .Y(n_499) );
AO32x2_ASAP7_75t_L g197 ( .A1(n_69), .A2(n_191), .A3(n_192), .B1(n_198), .B2(n_202), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_70), .B(n_176), .Y(n_555) );
INVx1_ASAP7_75t_L g248 ( .A(n_71), .Y(n_248) );
INVx1_ASAP7_75t_L g173 ( .A(n_72), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_73), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_74), .A2(n_103), .B1(n_114), .B2(n_765), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_75), .B(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_76), .A2(n_465), .B(n_501), .C(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_77), .B(n_757), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_77), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_78), .B(n_152), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_79), .Y(n_533) );
INVx1_ASAP7_75t_L g113 ( .A(n_80), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_81), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_83), .B(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_84), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_85), .B(n_152), .Y(n_179) );
INVx2_ASAP7_75t_L g141 ( .A(n_86), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_87), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_88), .B(n_162), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_89), .B(n_152), .Y(n_219) );
INVx2_ASAP7_75t_L g110 ( .A(n_90), .Y(n_110) );
OR2x2_ASAP7_75t_L g118 ( .A(n_90), .B(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g448 ( .A(n_90), .B(n_120), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_92), .A2(n_101), .B1(n_152), .B2(n_153), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_93), .B(n_462), .Y(n_494) );
INVx1_ASAP7_75t_L g498 ( .A(n_94), .Y(n_498) );
INVxp67_ASAP7_75t_L g536 ( .A(n_95), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_96), .B(n_152), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_97), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g511 ( .A(n_98), .Y(n_511) );
INVx1_ASAP7_75t_L g551 ( .A(n_99), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_100), .Y(n_126) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx12_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g766 ( .A(n_106), .Y(n_766) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
OR2x2_ASAP7_75t_L g742 ( .A(n_110), .B(n_120), .Y(n_742) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_110), .B(n_119), .Y(n_750) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_123), .Y(n_115) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g764 ( .A(n_118), .Y(n_764) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
OAI32xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_747), .A3(n_751), .B1(n_752), .B2(n_755), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_128), .B1(n_743), .B2(n_744), .Y(n_124) );
INVx1_ASAP7_75t_L g743 ( .A(n_125), .Y(n_743) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22x1_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_446), .B1(n_449), .B2(n_740), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_131), .A2(n_450), .B1(n_740), .B2(n_746), .Y(n_745) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_132), .A2(n_133), .B1(n_758), .B2(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_367), .Y(n_133) );
NAND5xp2_ASAP7_75t_L g134 ( .A(n_135), .B(n_286), .C(n_301), .D(n_327), .E(n_349), .Y(n_134) );
NOR2xp33_ASAP7_75t_SL g135 ( .A(n_136), .B(n_266), .Y(n_135) );
OAI221xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_203), .B1(n_239), .B2(n_255), .C(n_256), .Y(n_136) );
NOR2xp33_ASAP7_75t_SL g137 ( .A(n_138), .B(n_193), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_138), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g443 ( .A(n_138), .Y(n_443) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_166), .Y(n_138) );
INVx1_ASAP7_75t_L g283 ( .A(n_139), .Y(n_283) );
AND2x2_ASAP7_75t_L g285 ( .A(n_139), .B(n_184), .Y(n_285) );
AND2x2_ASAP7_75t_L g295 ( .A(n_139), .B(n_183), .Y(n_295) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_139), .Y(n_313) );
INVx1_ASAP7_75t_L g323 ( .A(n_139), .Y(n_323) );
OR2x2_ASAP7_75t_L g361 ( .A(n_139), .B(n_260), .Y(n_361) );
INVx2_ASAP7_75t_L g411 ( .A(n_139), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_139), .B(n_259), .Y(n_428) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_145), .B(n_165), .Y(n_139) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_140), .A2(n_170), .B(n_182), .Y(n_169) );
INVx2_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
INVx1_ASAP7_75t_L g475 ( .A(n_140), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_140), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_140), .A2(n_521), .B(n_522), .Y(n_520) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_L g190 ( .A(n_141), .B(n_142), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_157), .B(n_163), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_151), .B(n_154), .Y(n_146) );
INVx3_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_148), .Y(n_513) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
BUFx3_ASAP7_75t_L g200 ( .A(n_149), .Y(n_200) );
AND2x6_ASAP7_75t_L g465 ( .A(n_149), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g153 ( .A(n_150), .Y(n_153) );
INVx1_ASAP7_75t_L g224 ( .A(n_150), .Y(n_224) );
INVx2_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_156), .Y(n_162) );
INVx3_ASAP7_75t_L g176 ( .A(n_156), .Y(n_176) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
AND2x2_ASAP7_75t_L g463 ( .A(n_156), .B(n_224), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_156), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_161), .Y(n_157) );
O2A1O1Ixp5_ASAP7_75t_L g247 ( .A1(n_161), .A2(n_235), .B(n_248), .C(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_162), .A2(n_186), .B1(n_187), .B2(n_188), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g198 ( .A1(n_162), .A2(n_176), .B1(n_199), .B2(n_201), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_162), .A2(n_187), .B1(n_211), .B2(n_212), .Y(n_210) );
INVx4_ASAP7_75t_L g486 ( .A(n_162), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_163), .A2(n_171), .B(n_177), .Y(n_170) );
BUFx3_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_163), .A2(n_217), .B(n_220), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_163), .A2(n_229), .B(n_234), .Y(n_228) );
AND2x4_ASAP7_75t_L g462 ( .A(n_163), .B(n_463), .Y(n_462) );
INVx4_ASAP7_75t_SL g488 ( .A(n_163), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g552 ( .A(n_163), .B(n_463), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g166 ( .A(n_167), .B(n_183), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_168), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_168), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_SL g343 ( .A(n_168), .B(n_283), .Y(n_343) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_169), .Y(n_195) );
INVx2_ASAP7_75t_L g260 ( .A(n_169), .Y(n_260) );
OR2x2_ASAP7_75t_L g322 ( .A(n_169), .B(n_323), .Y(n_322) );
O2A1O1Ixp5_ASAP7_75t_SL g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_175), .Y(n_171) );
INVx2_ASAP7_75t_L g187 ( .A(n_175), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_175), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_175), .A2(n_245), .B(n_246), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_175), .B(n_536), .Y(n_535) );
INVx5_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_180), .Y(n_177) );
INVx1_ASAP7_75t_L g233 ( .A(n_180), .Y(n_233) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g469 ( .A(n_181), .Y(n_469) );
AND2x2_ASAP7_75t_L g261 ( .A(n_183), .B(n_197), .Y(n_261) );
AND2x2_ASAP7_75t_L g278 ( .A(n_183), .B(n_258), .Y(n_278) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g196 ( .A(n_184), .B(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g281 ( .A(n_184), .Y(n_281) );
AND2x2_ASAP7_75t_L g410 ( .A(n_184), .B(n_411), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_187), .A2(n_221), .B(n_222), .Y(n_220) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_187), .A2(n_235), .B(n_236), .C(n_237), .Y(n_234) );
INVx2_ASAP7_75t_L g227 ( .A(n_189), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_189), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_190), .Y(n_192) );
NAND3xp33_ASAP7_75t_L g209 ( .A(n_191), .B(n_210), .C(n_213), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_191), .A2(n_244), .B(n_247), .Y(n_243) );
INVx4_ASAP7_75t_L g213 ( .A(n_192), .Y(n_213) );
OA21x2_ASAP7_75t_L g215 ( .A1(n_192), .A2(n_216), .B(n_225), .Y(n_215) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_192), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_192), .A2(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g255 ( .A(n_193), .Y(n_255) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_196), .Y(n_193) );
AND2x2_ASAP7_75t_L g373 ( .A(n_194), .B(n_261), .Y(n_373) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g374 ( .A(n_195), .B(n_285), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_196), .A2(n_342), .B(n_344), .C(n_346), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_196), .B(n_342), .Y(n_351) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_196), .A2(n_272), .B1(n_415), .B2(n_416), .C(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g258 ( .A(n_197), .Y(n_258) );
INVx1_ASAP7_75t_L g294 ( .A(n_197), .Y(n_294) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_197), .Y(n_303) );
INVx2_ASAP7_75t_L g487 ( .A(n_200), .Y(n_487) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_200), .Y(n_500) );
INVx1_ASAP7_75t_L g472 ( .A(n_202), .Y(n_472) );
INVx1_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_214), .Y(n_204) );
AND2x2_ASAP7_75t_L g320 ( .A(n_205), .B(n_265), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_205), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_206), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g412 ( .A(n_206), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g444 ( .A(n_206), .Y(n_444) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g274 ( .A(n_207), .Y(n_274) );
AND2x2_ASAP7_75t_L g300 ( .A(n_207), .B(n_254), .Y(n_300) );
NOR2x1_ASAP7_75t_L g309 ( .A(n_207), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g316 ( .A(n_207), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
INVx1_ASAP7_75t_L g252 ( .A(n_208), .Y(n_252) );
AO21x1_ASAP7_75t_L g251 ( .A1(n_210), .A2(n_213), .B(n_252), .Y(n_251) );
INVx3_ASAP7_75t_L g478 ( .A(n_213), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_213), .B(n_503), .Y(n_502) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_213), .A2(n_508), .B(n_515), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_213), .B(n_516), .Y(n_515) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_213), .A2(n_550), .B(n_557), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_214), .B(n_356), .Y(n_391) );
INVx1_ASAP7_75t_SL g395 ( .A(n_214), .Y(n_395) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_226), .Y(n_214) );
INVx3_ASAP7_75t_L g254 ( .A(n_215), .Y(n_254) );
AND2x2_ASAP7_75t_L g265 ( .A(n_215), .B(n_242), .Y(n_265) );
AND2x2_ASAP7_75t_L g287 ( .A(n_215), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g332 ( .A(n_215), .B(n_326), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_215), .B(n_264), .Y(n_413) );
INVx2_ASAP7_75t_L g235 ( .A(n_223), .Y(n_235) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g253 ( .A(n_226), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g264 ( .A(n_226), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_226), .B(n_242), .Y(n_289) );
AND2x2_ASAP7_75t_L g325 ( .A(n_226), .B(n_326), .Y(n_325) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_238), .Y(n_226) );
OA21x2_ASAP7_75t_L g242 ( .A1(n_227), .A2(n_243), .B(n_250), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .C(n_233), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_231), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_231), .A2(n_555), .B(n_556), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_L g510 ( .A1(n_233), .A2(n_511), .B(n_512), .C(n_513), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_235), .A2(n_468), .B(n_470), .Y(n_467) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_253), .Y(n_240) );
INVx1_ASAP7_75t_L g305 ( .A(n_241), .Y(n_305) );
AND2x2_ASAP7_75t_L g347 ( .A(n_241), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_241), .B(n_268), .Y(n_353) );
AOI21xp5_ASAP7_75t_SL g427 ( .A1(n_241), .A2(n_259), .B(n_282), .Y(n_427) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_251), .Y(n_241) );
OR2x2_ASAP7_75t_L g270 ( .A(n_242), .B(n_251), .Y(n_270) );
AND2x2_ASAP7_75t_L g317 ( .A(n_242), .B(n_254), .Y(n_317) );
INVx2_ASAP7_75t_L g326 ( .A(n_242), .Y(n_326) );
INVx1_ASAP7_75t_L g432 ( .A(n_242), .Y(n_432) );
AND2x2_ASAP7_75t_L g356 ( .A(n_251), .B(n_326), .Y(n_356) );
INVx1_ASAP7_75t_L g381 ( .A(n_251), .Y(n_381) );
AND2x2_ASAP7_75t_L g290 ( .A(n_253), .B(n_274), .Y(n_290) );
AND2x2_ASAP7_75t_L g302 ( .A(n_253), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_SL g420 ( .A(n_253), .Y(n_420) );
INVx2_ASAP7_75t_L g310 ( .A(n_254), .Y(n_310) );
AND2x2_ASAP7_75t_L g348 ( .A(n_254), .B(n_264), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_254), .B(n_432), .Y(n_431) );
OAI21xp33_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_261), .B(n_262), .Y(n_256) );
AND2x2_ASAP7_75t_L g363 ( .A(n_257), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g417 ( .A(n_257), .Y(n_417) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g337 ( .A(n_258), .Y(n_337) );
BUFx2_ASAP7_75t_L g436 ( .A(n_258), .Y(n_436) );
BUFx2_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
AND2x2_ASAP7_75t_L g409 ( .A(n_259), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g392 ( .A(n_260), .Y(n_392) );
AND2x4_ASAP7_75t_L g319 ( .A(n_261), .B(n_282), .Y(n_319) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_261), .B(n_343), .Y(n_355) );
AOI32xp33_ASAP7_75t_L g279 ( .A1(n_262), .A2(n_280), .A3(n_282), .B1(n_284), .B2(n_285), .Y(n_279) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
INVx3_ASAP7_75t_L g268 ( .A(n_263), .Y(n_268) );
OR2x2_ASAP7_75t_L g404 ( .A(n_263), .B(n_360), .Y(n_404) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g273 ( .A(n_264), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g380 ( .A(n_264), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g272 ( .A(n_265), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g284 ( .A(n_265), .B(n_274), .Y(n_284) );
INVx1_ASAP7_75t_L g405 ( .A(n_265), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_265), .B(n_380), .Y(n_438) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_271), .B(n_275), .C(n_279), .Y(n_266) );
OAI322xp33_ASAP7_75t_L g375 ( .A1(n_267), .A2(n_312), .A3(n_376), .B1(n_378), .B2(n_382), .C1(n_383), .C2(n_387), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVxp67_ASAP7_75t_L g340 ( .A(n_268), .Y(n_340) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g394 ( .A(n_270), .B(n_395), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_270), .B(n_310), .Y(n_441) );
INVxp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g333 ( .A(n_273), .Y(n_333) );
OR2x2_ASAP7_75t_L g419 ( .A(n_274), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_277), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g328 ( .A(n_278), .B(n_307), .Y(n_328) );
AND2x2_ASAP7_75t_L g399 ( .A(n_278), .B(n_312), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_278), .B(n_386), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_280), .A2(n_287), .B1(n_290), .B2(n_291), .C(n_296), .Y(n_286) );
OR2x2_ASAP7_75t_L g297 ( .A(n_280), .B(n_293), .Y(n_297) );
AND2x2_ASAP7_75t_L g385 ( .A(n_280), .B(n_386), .Y(n_385) );
AOI32xp33_ASAP7_75t_L g424 ( .A1(n_280), .A2(n_310), .A3(n_425), .B1(n_426), .B2(n_429), .Y(n_424) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND3xp33_ASAP7_75t_L g358 ( .A(n_281), .B(n_317), .C(n_340), .Y(n_358) );
AND2x2_ASAP7_75t_L g384 ( .A(n_281), .B(n_377), .Y(n_384) );
INVxp67_ASAP7_75t_L g364 ( .A(n_282), .Y(n_364) );
BUFx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_285), .B(n_337), .Y(n_393) );
INVx2_ASAP7_75t_L g403 ( .A(n_285), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_285), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g372 ( .A(n_288), .Y(n_372) );
OR2x2_ASAP7_75t_L g298 ( .A(n_289), .B(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_291), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_295), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_294), .Y(n_377) );
AND2x2_ASAP7_75t_L g336 ( .A(n_295), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g382 ( .A(n_295), .Y(n_382) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_295), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AOI21xp33_ASAP7_75t_SL g321 ( .A1(n_297), .A2(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g415 ( .A(n_300), .B(n_325), .Y(n_415) );
AOI211xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_304), .B(n_314), .C(n_321), .Y(n_301) );
AND2x2_ASAP7_75t_L g345 ( .A(n_303), .B(n_313), .Y(n_345) );
INVx2_ASAP7_75t_L g360 ( .A(n_303), .Y(n_360) );
OR2x2_ASAP7_75t_L g398 ( .A(n_303), .B(n_361), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_303), .B(n_441), .Y(n_440) );
AOI211xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_306), .B(n_308), .C(n_311), .Y(n_304) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_307), .B(n_345), .Y(n_344) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_308), .A2(n_403), .B(n_427), .C(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g324 ( .A(n_309), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g366 ( .A(n_310), .B(n_356), .Y(n_366) );
INVx1_ASAP7_75t_L g371 ( .A(n_310), .Y(n_371) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_315), .B(n_318), .Y(n_314) );
INVxp33_ASAP7_75t_L g422 ( .A(n_316), .Y(n_422) );
AND2x2_ASAP7_75t_L g401 ( .A(n_317), .B(n_380), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_322), .A2(n_384), .B(n_385), .Y(n_383) );
OAI322xp33_ASAP7_75t_L g402 ( .A1(n_324), .A2(n_403), .A3(n_404), .B1(n_405), .B2(n_406), .C1(n_408), .C2(n_412), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_329), .B1(n_334), .B2(n_338), .C(n_341), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g379 ( .A(n_332), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g423 ( .A(n_336), .Y(n_423) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_339), .B(n_359), .Y(n_425) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g388 ( .A(n_348), .B(n_356), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_352), .B1(n_354), .B2(n_356), .C(n_357), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_352), .A2(n_369), .B1(n_373), .B2(n_374), .C(n_375), .Y(n_368) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_356), .B(n_371), .Y(n_370) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_362), .B2(n_365), .Y(n_357) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx2_ASAP7_75t_SL g386 ( .A(n_361), .Y(n_386) );
INVxp67_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND5xp2_ASAP7_75t_L g367 ( .A(n_368), .B(n_389), .C(n_414), .D(n_424), .E(n_434), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_372), .Y(n_369) );
NOR4xp25_ASAP7_75t_L g442 ( .A(n_371), .B(n_377), .C(n_443), .D(n_444), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g434 ( .A1(n_374), .A2(n_435), .B1(n_437), .B2(n_439), .C(n_442), .Y(n_434) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g433 ( .A(n_380), .Y(n_433) );
OAI322xp33_ASAP7_75t_L g390 ( .A1(n_384), .A2(n_391), .A3(n_392), .B1(n_393), .B2(n_394), .C1(n_396), .C2(n_400), .Y(n_390) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_402), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g435 ( .A(n_410), .B(n_436), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g746 ( .A(n_447), .Y(n_746) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_SL g450 ( .A(n_451), .B(n_695), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_630), .Y(n_451) );
NAND4xp25_ASAP7_75t_SL g452 ( .A(n_453), .B(n_575), .C(n_599), .D(n_622), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_517), .B1(n_547), .B2(n_559), .C(n_562), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_490), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_456), .A2(n_476), .B1(n_518), .B2(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_456), .B(n_491), .Y(n_633) );
AND2x2_ASAP7_75t_L g652 ( .A(n_456), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_456), .B(n_636), .Y(n_722) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_476), .Y(n_456) );
AND2x2_ASAP7_75t_L g590 ( .A(n_457), .B(n_491), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_457), .B(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g613 ( .A(n_457), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g618 ( .A(n_457), .B(n_477), .Y(n_618) );
INVx2_ASAP7_75t_L g650 ( .A(n_457), .Y(n_650) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_457), .Y(n_694) );
AND2x2_ASAP7_75t_L g711 ( .A(n_457), .B(n_588), .Y(n_711) );
INVx5_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g629 ( .A(n_458), .B(n_588), .Y(n_629) );
AND2x4_ASAP7_75t_L g643 ( .A(n_458), .B(n_476), .Y(n_643) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_458), .Y(n_647) );
AND2x2_ASAP7_75t_L g667 ( .A(n_458), .B(n_582), .Y(n_667) );
AND2x2_ASAP7_75t_L g717 ( .A(n_458), .B(n_492), .Y(n_717) );
AND2x2_ASAP7_75t_L g727 ( .A(n_458), .B(n_477), .Y(n_727) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_473), .Y(n_458) );
AOI21xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_464), .B(n_472), .Y(n_459) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx5_ASAP7_75t_L g482 ( .A(n_465), .Y(n_482) );
INVx2_ASAP7_75t_L g471 ( .A(n_469), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_471), .A2(n_498), .B(n_499), .C(n_500), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_471), .A2(n_500), .B(n_524), .C(n_525), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
AND2x2_ASAP7_75t_L g583 ( .A(n_476), .B(n_491), .Y(n_583) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_476), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_476), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g673 ( .A(n_476), .Y(n_673) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g561 ( .A(n_477), .B(n_506), .Y(n_561) );
AND2x2_ASAP7_75t_L g588 ( .A(n_477), .B(n_507), .Y(n_588) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_489), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_482), .B(n_483), .C(n_488), .Y(n_480) );
INVx2_ASAP7_75t_L g496 ( .A(n_482), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_482), .A2(n_488), .B(n_533), .C(n_534), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g501 ( .A(n_488), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_490), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_504), .Y(n_490) );
OR2x2_ASAP7_75t_L g614 ( .A(n_491), .B(n_505), .Y(n_614) );
AND2x2_ASAP7_75t_L g651 ( .A(n_491), .B(n_561), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_491), .B(n_582), .Y(n_662) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_491), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_491), .B(n_618), .Y(n_735) );
INVx5_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g560 ( .A(n_492), .Y(n_560) );
AND2x2_ASAP7_75t_L g569 ( .A(n_492), .B(n_505), .Y(n_569) );
AND2x2_ASAP7_75t_L g685 ( .A(n_492), .B(n_580), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_492), .B(n_618), .Y(n_707) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_502), .Y(n_492) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_505), .Y(n_653) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_506), .Y(n_605) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g582 ( .A(n_507), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_527), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_518), .B(n_595), .Y(n_714) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_519), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g566 ( .A(n_519), .B(n_567), .Y(n_566) );
INVx5_ASAP7_75t_SL g574 ( .A(n_519), .Y(n_574) );
OR2x2_ASAP7_75t_L g597 ( .A(n_519), .B(n_567), .Y(n_597) );
OR2x2_ASAP7_75t_L g607 ( .A(n_519), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g670 ( .A(n_519), .B(n_529), .Y(n_670) );
AND2x2_ASAP7_75t_SL g708 ( .A(n_519), .B(n_528), .Y(n_708) );
NOR4xp25_ASAP7_75t_L g729 ( .A(n_519), .B(n_650), .C(n_730), .D(n_731), .Y(n_729) );
AND2x2_ASAP7_75t_L g739 ( .A(n_519), .B(n_571), .Y(n_739) );
OR2x6_ASAP7_75t_L g519 ( .A(n_520), .B(n_526), .Y(n_519) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g564 ( .A(n_528), .B(n_560), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_528), .B(n_566), .Y(n_733) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
OR2x2_ASAP7_75t_L g573 ( .A(n_529), .B(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g580 ( .A(n_529), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_529), .B(n_549), .Y(n_592) );
INVxp67_ASAP7_75t_L g595 ( .A(n_529), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_529), .B(n_567), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_529), .B(n_539), .Y(n_661) );
AND2x2_ASAP7_75t_L g676 ( .A(n_529), .B(n_571), .Y(n_676) );
OR2x2_ASAP7_75t_L g705 ( .A(n_529), .B(n_539), .Y(n_705) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_537), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_538), .B(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_538), .B(n_574), .Y(n_713) );
OR2x2_ASAP7_75t_L g734 ( .A(n_538), .B(n_611), .Y(n_734) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g548 ( .A(n_539), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g571 ( .A(n_539), .B(n_567), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_539), .B(n_549), .Y(n_586) );
AND2x2_ASAP7_75t_L g656 ( .A(n_539), .B(n_580), .Y(n_656) );
AND2x2_ASAP7_75t_L g690 ( .A(n_539), .B(n_574), .Y(n_690) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_540), .B(n_574), .Y(n_593) );
AND2x2_ASAP7_75t_L g621 ( .A(n_540), .B(n_549), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_547), .B(n_629), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_548), .A2(n_636), .B1(n_672), .B2(n_689), .C(n_691), .Y(n_688) );
INVx5_ASAP7_75t_SL g567 ( .A(n_549), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .B(n_553), .Y(n_550) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
OAI33xp33_ASAP7_75t_L g587 ( .A1(n_560), .A2(n_588), .A3(n_589), .B1(n_591), .B2(n_594), .B3(n_598), .Y(n_587) );
OR2x2_ASAP7_75t_L g603 ( .A(n_560), .B(n_604), .Y(n_603) );
AOI322xp5_ASAP7_75t_L g712 ( .A1(n_560), .A2(n_629), .A3(n_636), .B1(n_713), .B2(n_714), .C1(n_715), .C2(n_718), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_560), .B(n_588), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_SL g736 ( .A1(n_560), .A2(n_588), .B(n_737), .C(n_739), .Y(n_736) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_561), .A2(n_576), .B1(n_581), .B2(n_584), .C(n_587), .Y(n_575) );
INVx1_ASAP7_75t_L g668 ( .A(n_561), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_561), .B(n_717), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .B1(n_568), .B2(n_570), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g645 ( .A(n_566), .B(n_580), .Y(n_645) );
AND2x2_ASAP7_75t_L g703 ( .A(n_566), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g611 ( .A(n_567), .B(n_574), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_567), .B(n_580), .Y(n_639) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_569), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_569), .B(n_647), .Y(n_701) );
OAI321xp33_ASAP7_75t_L g720 ( .A1(n_569), .A2(n_642), .A3(n_721), .B1(n_722), .B2(n_723), .C(n_724), .Y(n_720) );
INVx1_ASAP7_75t_L g687 ( .A(n_570), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_571), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g626 ( .A(n_571), .B(n_574), .Y(n_626) );
AOI321xp33_ASAP7_75t_L g684 ( .A1(n_571), .A2(n_588), .A3(n_685), .B1(n_686), .B2(n_687), .C(n_688), .Y(n_684) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g601 ( .A(n_573), .B(n_586), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_574), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_574), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_574), .B(n_660), .Y(n_697) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g620 ( .A(n_578), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g585 ( .A(n_579), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g693 ( .A(n_580), .Y(n_693) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_583), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g616 ( .A(n_588), .Y(n_616) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_590), .B(n_625), .Y(n_674) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
OR2x2_ASAP7_75t_L g638 ( .A(n_593), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g683 ( .A(n_593), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_594), .A2(n_641), .B1(n_644), .B2(n_646), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g738 ( .A(n_597), .B(n_661), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_602), .B1(n_606), .B2(n_612), .C(n_615), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx2_ASAP7_75t_L g636 ( .A(n_605), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_SL g682 ( .A(n_608), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_610), .B(n_660), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_610), .A2(n_678), .B(n_680), .Y(n_677) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g723 ( .A(n_611), .B(n_705), .Y(n_723) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_SL g625 ( .A(n_614), .Y(n_625) );
AOI21xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B(n_619), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g669 ( .A(n_621), .B(n_670), .Y(n_669) );
INVxp67_ASAP7_75t_L g731 ( .A(n_621), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B(n_627), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_625), .B(n_643), .Y(n_679) );
INVxp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g700 ( .A(n_629), .Y(n_700) );
NAND5xp2_ASAP7_75t_L g630 ( .A(n_631), .B(n_648), .C(n_657), .D(n_677), .E(n_684), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B(n_637), .C(n_640), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g672 ( .A(n_636), .Y(n_672) );
CKINVDCx16_ASAP7_75t_R g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_644), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g686 ( .A(n_646), .Y(n_686) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_652), .B(n_654), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_649), .A2(n_703), .B1(n_706), .B2(n_708), .C(n_709), .Y(n_702) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
AOI321xp33_ASAP7_75t_L g657 ( .A1(n_650), .A2(n_658), .A3(n_662), .B1(n_663), .B2(n_669), .C(n_671), .Y(n_657) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g728 ( .A(n_662), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_664), .B(n_668), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g680 ( .A(n_665), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NOR2xp67_ASAP7_75t_SL g692 ( .A(n_666), .B(n_673), .Y(n_692) );
AOI321xp33_ASAP7_75t_SL g724 ( .A1(n_669), .A2(n_725), .A3(n_726), .B1(n_727), .B2(n_728), .C(n_729), .Y(n_724) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_674), .C(n_675), .Y(n_671) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_682), .B(n_690), .Y(n_719) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .C(n_694), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_720), .C(n_732), .Y(n_695) );
OAI211xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_698), .B(n_702), .C(n_712), .Y(n_696) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_700), .B(n_701), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g732 ( .A1(n_701), .A2(n_733), .B1(n_734), .B2(n_735), .C(n_736), .Y(n_732) );
INVx1_ASAP7_75t_L g721 ( .A(n_703), .Y(n_721) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g725 ( .A(n_723), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
CKINVDCx14_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx3_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
BUFx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NOR3xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_761), .C(n_764), .Y(n_755) );
INVx1_ASAP7_75t_L g763 ( .A(n_757), .Y(n_763) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
endmodule