module fake_jpeg_18306_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_5),
.B(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_6),
.B(n_11),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_5),
.B(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_28),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_26),
.B(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_33),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_14),
.B1(n_32),
.B2(n_27),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_54),
.B1(n_37),
.B2(n_47),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_27),
.B1(n_36),
.B2(n_35),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_19),
.B1(n_35),
.B2(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_62),
.B1(n_64),
.B2(n_37),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_46),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_18),
.B1(n_22),
.B2(n_13),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_13),
.B1(n_22),
.B2(n_16),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_24),
.B(n_17),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_16),
.B1(n_17),
.B2(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_26),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_72),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_39),
.C(n_50),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_23),
.B(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_76),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_49),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_78),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_23),
.B(n_2),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_17),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_80),
.B1(n_44),
.B2(n_61),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_54),
.B1(n_57),
.B2(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_84),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_17),
.B(n_57),
.C(n_23),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_88),
.B(n_93),
.Y(n_103)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_23),
.B(n_15),
.C(n_53),
.D(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_90),
.B(n_56),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_78),
.C(n_69),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_53),
.C(n_42),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_83),
.A2(n_70),
.B1(n_74),
.B2(n_80),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_71),
.B1(n_67),
.B2(n_44),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_89),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_98),
.B(n_100),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_101),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_56),
.B(n_3),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_81),
.C(n_89),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_112),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_88),
.C(n_84),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_100),
.B1(n_95),
.B2(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_101),
.C(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_118),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_96),
.C(n_104),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_92),
.A3(n_82),
.B1(n_102),
.B2(n_85),
.C1(n_9),
.C2(n_11),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_120),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_111),
.C(n_9),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_106),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_119),
.C(n_3),
.Y(n_126)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_123),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_129),
.B(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_1),
.Y(n_129)
);

AOI31xp67_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_122),
.A3(n_4),
.B(n_7),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_1),
.C(n_4),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);


endmodule