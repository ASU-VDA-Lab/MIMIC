module fake_aes_9992_n_43 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_43);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx3_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_8), .B(n_13), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_4), .B(n_2), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_10), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_6), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_0), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_5), .Y(n_21) );
OAI22xp5_ASAP7_75t_L g22 ( .A1(n_12), .A2(n_9), .B1(n_3), .B2(n_7), .Y(n_22) );
NAND2xp5_ASAP7_75t_SL g23 ( .A(n_15), .B(n_0), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_20), .B(n_1), .Y(n_25) );
OAI21x1_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_21), .B(n_19), .Y(n_26) );
A2O1A1Ixp33_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_16), .B(n_18), .C(n_17), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_27), .B(n_25), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
INVx1_ASAP7_75t_SL g33 ( .A(n_30), .Y(n_33) );
NAND2xp33_ASAP7_75t_L g34 ( .A(n_32), .B(n_22), .Y(n_34) );
BUFx2_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
NOR3xp33_ASAP7_75t_L g37 ( .A(n_34), .B(n_23), .C(n_16), .Y(n_37) );
INVxp67_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
INVx1_ASAP7_75t_SL g39 ( .A(n_35), .Y(n_39) );
BUFx2_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
OAI22xp5_ASAP7_75t_SL g41 ( .A1(n_38), .A2(n_34), .B1(n_2), .B2(n_3), .Y(n_41) );
AOI22xp33_ASAP7_75t_L g42 ( .A1(n_41), .A2(n_37), .B1(n_26), .B2(n_1), .Y(n_42) );
OAI21xp5_ASAP7_75t_L g43 ( .A1(n_42), .A2(n_40), .B(n_14), .Y(n_43) );
endmodule