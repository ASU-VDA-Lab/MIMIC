module real_jpeg_32979_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_215;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_0),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_0),
.Y(n_245)
);

AOI22x1_ASAP7_75t_L g46 ( 
.A1(n_1),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_96),
.B1(n_103),
.B2(n_107),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_2),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_2),
.A2(n_107),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_3),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_4),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g16 ( 
.A1(n_5),
.A2(n_17),
.A3(n_21),
.B1(n_24),
.B2(n_35),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_5),
.A2(n_36),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g248 ( 
.A1(n_5),
.A2(n_168),
.B(n_180),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_62),
.B1(n_66),
.B2(n_67),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_6),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_6),
.A2(n_66),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

OAI22x1_ASAP7_75t_SL g154 ( 
.A1(n_6),
.A2(n_66),
.B1(n_155),
.B2(n_159),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_7),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_8),
.A2(n_92),
.B1(n_96),
.B2(n_100),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_8),
.A2(n_100),
.B1(n_226),
.B2(n_229),
.Y(n_225)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_9),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_186),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_183),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_145),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_145),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_71),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_42),
.Y(n_15)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_20),
.Y(n_119)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_23),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_23),
.Y(n_130)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_23),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_34),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_R g165 ( 
.A(n_36),
.B(n_111),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_36),
.B(n_211),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_36),
.A2(n_210),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_36),
.B(n_149),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_36),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_40),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_41),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_55),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_45),
.Y(n_182)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_49),
.Y(n_194)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx2_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_54),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_55),
.A2(n_225),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_56),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_56),
.A2(n_224),
.B1(n_233),
.B2(n_236),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_60),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_60),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_60),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_61),
.B(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22x1_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_80),
.B1(n_86),
.B2(n_88),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_108),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_91),
.B1(n_101),
.B2(n_102),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_73),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_85),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_80),
.B2(n_83),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_82),
.Y(n_209)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp67_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_86),
.Y(n_207)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_131),
.B(n_135),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_111)
);

INVx5_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.Y(n_120)
);

BUFx4f_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_164),
.C(n_166),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_147),
.A2(n_148),
.B1(n_164),
.B2(n_165),
.Y(n_218)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.B(n_153),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_154),
.Y(n_213)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_215),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_218),
.Y(n_217)
);

OAI21x1_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B(n_180),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_219),
.Y(n_186)
);

INVxp67_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_217),
.Y(n_188)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_212),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_212),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_195),
.B(n_206),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx4f_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B(n_210),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_217),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_260),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_238),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_237),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_237),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx2_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

OAI21x1_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_247),
.B(n_259),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_242),
.B(n_246),
.Y(n_259)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx4f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);


endmodule