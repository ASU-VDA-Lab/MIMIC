module real_aes_15695_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_860, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_860;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g120 ( .A(n_0), .B(n_121), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_1), .A2(n_33), .B1(n_156), .B2(n_192), .Y(n_191) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_2), .A2(n_9), .B1(n_146), .B2(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g121 ( .A(n_3), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_4), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_5), .A2(n_10), .B1(n_205), .B2(n_208), .Y(n_204) );
OR2x2_ASAP7_75t_L g111 ( .A(n_6), .B(n_29), .Y(n_111) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_7), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_8), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_11), .B(n_147), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_12), .A2(n_101), .B1(n_146), .B2(n_149), .Y(n_145) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_13), .A2(n_30), .B1(n_181), .B2(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_14), .B(n_147), .Y(n_178) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_15), .A2(n_44), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_16), .B(n_548), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_17), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_18), .A2(n_89), .B1(n_812), .B2(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_18), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_19), .A2(n_37), .B1(n_194), .B2(n_195), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g485 ( .A(n_20), .Y(n_485) );
XOR2x2_ASAP7_75t_L g124 ( .A(n_21), .B(n_125), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_22), .A2(n_42), .B1(n_146), .B2(n_195), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_23), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_24), .B(n_181), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_25), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_26), .B(n_206), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_27), .B(n_187), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_28), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_31), .A2(n_83), .B1(n_156), .B2(n_233), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_32), .A2(n_36), .B1(n_156), .B2(n_177), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_34), .A2(n_47), .B1(n_146), .B2(n_155), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_35), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_38), .B(n_147), .Y(n_533) );
INVx2_ASAP7_75t_L g119 ( .A(n_39), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_40), .B(n_152), .Y(n_543) );
BUFx3_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
INVx1_ASAP7_75t_L g823 ( .A(n_41), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_43), .B(n_493), .Y(n_550) );
AND2x2_ASAP7_75t_L g492 ( .A(n_45), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_46), .B(n_221), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_48), .B(n_206), .Y(n_515) );
XOR2xp5_ASAP7_75t_L g123 ( .A(n_49), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_50), .B(n_194), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_51), .A2(n_90), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_51), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_52), .A2(n_71), .B1(n_155), .B2(n_194), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_53), .A2(n_74), .B1(n_156), .B2(n_177), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_54), .B(n_519), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_55), .A2(n_236), .B(n_484), .C(n_486), .Y(n_483) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_56), .A2(n_98), .B1(n_146), .B2(n_208), .Y(n_254) );
AND2x4_ASAP7_75t_L g142 ( .A(n_57), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g165 ( .A(n_58), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_59), .A2(n_60), .B1(n_195), .B2(n_224), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_61), .B(n_187), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_62), .B(n_493), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_63), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_64), .B(n_195), .Y(n_536) );
INVx1_ASAP7_75t_L g143 ( .A(n_65), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_66), .A2(n_830), .B1(n_853), .B2(n_855), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_67), .A2(n_227), .B1(n_830), .B2(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g831 ( .A(n_67), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_68), .A2(n_828), .B1(n_829), .B2(n_832), .Y(n_827) );
CKINVDCx14_ASAP7_75t_R g828 ( .A(n_68), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_69), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_70), .B(n_187), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_72), .B(n_156), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_73), .B(n_152), .C(n_192), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_75), .B(n_156), .Y(n_499) );
INVx2_ASAP7_75t_L g153 ( .A(n_76), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_77), .B(n_147), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_78), .B(n_211), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_79), .B(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_80), .A2(n_97), .B1(n_195), .B2(n_236), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_81), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_82), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_84), .A2(n_92), .B1(n_206), .B2(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_85), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_86), .B(n_147), .Y(n_569) );
NAND2xp33_ASAP7_75t_SL g598 ( .A(n_87), .B(n_182), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_88), .B(n_150), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_89), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g812 ( .A(n_89), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_90), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_91), .B(n_187), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_93), .Y(n_215) );
INVx1_ASAP7_75t_L g115 ( .A(n_94), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_94), .B(n_843), .Y(n_842) );
NAND2xp33_ASAP7_75t_L g183 ( .A(n_95), .B(n_147), .Y(n_183) );
NAND2xp33_ASAP7_75t_L g500 ( .A(n_96), .B(n_182), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_99), .B(n_493), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_100), .B(n_182), .C(n_211), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_102), .B(n_156), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_103), .B(n_206), .Y(n_517) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_122), .B(n_816), .Y(n_104) );
BUFx4f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx3_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_112), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g113 ( .A(n_109), .B(n_114), .Y(n_113) );
NOR2x1_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g825 ( .A(n_111), .Y(n_825) );
OR2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
AND2x2_ASAP7_75t_L g853 ( .A(n_113), .B(n_854), .Y(n_853) );
BUFx8_ASAP7_75t_SL g469 ( .A(n_114), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_114), .Y(n_815) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g824 ( .A(n_115), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_116), .B(n_839), .Y(n_854) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_117), .B(n_120), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g849 ( .A(n_118), .B(n_850), .Y(n_849) );
INVx3_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_119), .B(n_858), .Y(n_857) );
INVx2_ASAP7_75t_SL g851 ( .A(n_120), .Y(n_851) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_128), .Y(n_122) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_470), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_469), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_372), .Y(n_130) );
NAND4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_296), .C(n_327), .D(n_356), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_263), .Y(n_132) );
OAI322xp33_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_199), .A3(n_228), .B1(n_241), .B2(n_249), .C1(n_258), .C2(n_260), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_135), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_169), .Y(n_135) );
AND2x2_ASAP7_75t_L g293 ( .A(n_136), .B(n_294), .Y(n_293) );
INVx4_ASAP7_75t_L g329 ( .A(n_136), .Y(n_329) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g304 ( .A(n_137), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g307 ( .A(n_137), .B(n_201), .Y(n_307) );
AND2x2_ASAP7_75t_L g324 ( .A(n_137), .B(n_217), .Y(n_324) );
AND2x2_ASAP7_75t_L g422 ( .A(n_137), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g245 ( .A(n_138), .Y(n_245) );
AND2x4_ASAP7_75t_L g428 ( .A(n_138), .B(n_423), .Y(n_428) );
AO31x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_144), .A3(n_160), .B(n_166), .Y(n_138) );
AO31x2_ASAP7_75t_L g252 ( .A1(n_139), .A2(n_212), .A3(n_253), .B(n_256), .Y(n_252) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp67_ASAP7_75t_SL g481 ( .A(n_140), .B(n_161), .Y(n_481) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AO31x2_ASAP7_75t_L g189 ( .A1(n_141), .A2(n_190), .A3(n_196), .B(n_197), .Y(n_189) );
AO31x2_ASAP7_75t_L g202 ( .A1(n_141), .A2(n_203), .A3(n_212), .B(n_214), .Y(n_202) );
AO31x2_ASAP7_75t_L g217 ( .A1(n_141), .A2(n_218), .A3(n_225), .B(n_226), .Y(n_217) );
AO31x2_ASAP7_75t_L g552 ( .A1(n_141), .A2(n_162), .A3(n_553), .B(n_557), .Y(n_552) );
BUFx10_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
BUFx10_ASAP7_75t_L g508 ( .A(n_142), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_151), .B1(n_154), .B2(n_157), .Y(n_144) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g548 ( .A(n_147), .Y(n_548) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_147), .A2(n_594), .B(n_595), .Y(n_593) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g150 ( .A(n_148), .Y(n_150) );
INVx3_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_148), .Y(n_182) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_148), .Y(n_192) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_148), .Y(n_195) );
INVx1_ASAP7_75t_L g207 ( .A(n_148), .Y(n_207) );
INVx1_ASAP7_75t_L g221 ( .A(n_148), .Y(n_221) );
INVx1_ASAP7_75t_L g224 ( .A(n_148), .Y(n_224) );
INVx2_ASAP7_75t_L g234 ( .A(n_148), .Y(n_234) );
INVx1_ASAP7_75t_L g236 ( .A(n_148), .Y(n_236) );
O2A1O1Ixp5_ASAP7_75t_L g567 ( .A1(n_149), .A2(n_152), .B(n_568), .C(n_569), .Y(n_567) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_151), .A2(n_180), .B(n_183), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_151), .A2(n_157), .B1(n_191), .B2(n_193), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_151), .A2(n_204), .B1(n_209), .B2(n_210), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_151), .A2(n_157), .B1(n_219), .B2(n_222), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_151), .A2(n_232), .B1(n_235), .B2(n_237), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_151), .A2(n_210), .B1(n_254), .B2(n_255), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g272 ( .A1(n_151), .A2(n_157), .B1(n_273), .B2(n_274), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_151), .A2(n_157), .B1(n_554), .B2(n_556), .Y(n_553) );
INVx6_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
O2A1O1Ixp5_ASAP7_75t_L g175 ( .A1(n_152), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_152), .A2(n_535), .B(n_536), .Y(n_534) );
BUFx8_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
INVx1_ASAP7_75t_L g211 ( .A(n_153), .Y(n_211) );
INVx1_ASAP7_75t_L g487 ( .A(n_153), .Y(n_487) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx4_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
INVx1_ASAP7_75t_L g208 ( .A(n_156), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_156), .A2(n_195), .B1(n_490), .B2(n_491), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_157), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g520 ( .A(n_158), .Y(n_520) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g504 ( .A(n_159), .Y(n_504) );
AO31x2_ASAP7_75t_L g271 ( .A1(n_160), .A2(n_238), .A3(n_272), .B(n_275), .Y(n_271) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_SL g214 ( .A(n_162), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_162), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g168 ( .A(n_163), .Y(n_168) );
INVx2_ASAP7_75t_L g213 ( .A(n_163), .Y(n_213) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_164), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_168), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g493 ( .A(n_168), .Y(n_493) );
INVx2_ASAP7_75t_L g511 ( .A(n_168), .Y(n_511) );
AND2x4_ASAP7_75t_L g433 ( .A(n_169), .B(n_334), .Y(n_433) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g262 ( .A(n_170), .Y(n_262) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_170), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_188), .Y(n_170) );
AND2x2_ASAP7_75t_L g250 ( .A(n_171), .B(n_189), .Y(n_250) );
INVx1_ASAP7_75t_L g291 ( .A(n_171), .Y(n_291) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_174), .B(n_186), .Y(n_171) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_172), .A2(n_174), .B(n_186), .Y(n_286) );
INVx2_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g187 ( .A(n_173), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_173), .B(n_198), .Y(n_197) );
BUFx3_ASAP7_75t_L g225 ( .A(n_173), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_173), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_173), .B(n_257), .Y(n_256) );
AND2x4_ASAP7_75t_SL g507 ( .A(n_173), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g529 ( .A(n_173), .Y(n_529) );
INVx1_ASAP7_75t_SL g591 ( .A(n_173), .Y(n_591) );
OAI21x1_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_179), .B(n_184), .Y(n_174) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g194 ( .A(n_182), .Y(n_194) );
INVx2_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_SL g238 ( .A(n_185), .Y(n_238) );
INVx2_ASAP7_75t_L g196 ( .A(n_187), .Y(n_196) );
INVx2_ASAP7_75t_L g282 ( .A(n_188), .Y(n_282) );
AND2x2_ASAP7_75t_L g346 ( .A(n_188), .B(n_285), .Y(n_346) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g300 ( .A(n_189), .Y(n_300) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_189), .Y(n_353) );
OR2x2_ASAP7_75t_L g424 ( .A(n_189), .B(n_230), .Y(n_424) );
INVx2_ASAP7_75t_L g519 ( .A(n_192), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_195), .A2(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g555 ( .A(n_195), .Y(n_555) );
NAND4xp25_ASAP7_75t_L g302 ( .A(n_199), .B(n_303), .C(n_306), .D(n_308), .Y(n_302) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_L g440 ( .A(n_200), .B(n_428), .Y(n_440) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_216), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_201), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g294 ( .A(n_201), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g314 ( .A(n_201), .Y(n_314) );
INVx1_ASAP7_75t_L g331 ( .A(n_201), .Y(n_331) );
INVx1_ASAP7_75t_L g339 ( .A(n_201), .Y(n_339) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_201), .Y(n_453) );
INVx4_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_202), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g371 ( .A(n_202), .B(n_271), .Y(n_371) );
AND2x2_ASAP7_75t_L g379 ( .A(n_202), .B(n_217), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_202), .B(n_402), .Y(n_401) );
BUFx2_ASAP7_75t_L g444 ( .A(n_202), .Y(n_444) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g237 ( .A(n_211), .Y(n_237) );
INVx1_ASAP7_75t_L g549 ( .A(n_211), .Y(n_549) );
BUFx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_213), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g248 ( .A(n_217), .Y(n_248) );
OR2x2_ASAP7_75t_L g309 ( .A(n_217), .B(n_271), .Y(n_309) );
INVx2_ASAP7_75t_L g316 ( .A(n_217), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_217), .B(n_269), .Y(n_340) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_217), .Y(n_427) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AO31x2_ASAP7_75t_L g230 ( .A1(n_225), .A2(n_231), .A3(n_238), .B(n_239), .Y(n_230) );
INVx1_ASAP7_75t_L g830 ( .A(n_227), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_228), .B(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g251 ( .A(n_230), .B(n_252), .Y(n_251) );
BUFx2_ASAP7_75t_L g261 ( .A(n_230), .Y(n_261) );
INVx2_ASAP7_75t_L g279 ( .A(n_230), .Y(n_279) );
AND2x4_ASAP7_75t_L g311 ( .A(n_230), .B(n_283), .Y(n_311) );
OR2x2_ASAP7_75t_L g391 ( .A(n_230), .B(n_291), .Y(n_391) );
INVx2_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_234), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g505 ( .A(n_236), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_246), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_243), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g308 ( .A(n_243), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_243), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_244), .B(n_314), .Y(n_322) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g267 ( .A(n_245), .Y(n_267) );
OR2x2_ASAP7_75t_L g360 ( .A(n_245), .B(n_270), .Y(n_360) );
INVx1_ASAP7_75t_L g287 ( .A(n_246), .Y(n_287) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g259 ( .A(n_247), .Y(n_259) );
INVx1_ASAP7_75t_L g295 ( .A(n_248), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
OAI322xp33_ASAP7_75t_L g263 ( .A1(n_250), .A2(n_264), .A3(n_277), .B1(n_280), .B2(n_287), .C1(n_288), .C2(n_292), .Y(n_263) );
AND2x4_ASAP7_75t_L g310 ( .A(n_250), .B(n_311), .Y(n_310) );
AOI211xp5_ASAP7_75t_SL g341 ( .A1(n_250), .A2(n_342), .B(n_343), .C(n_347), .Y(n_341) );
AND2x2_ASAP7_75t_L g361 ( .A(n_250), .B(n_251), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_250), .B(n_278), .Y(n_367) );
AND2x4_ASAP7_75t_SL g289 ( .A(n_251), .B(n_290), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g380 ( .A(n_251), .B(n_307), .C(n_335), .Y(n_380) );
AND2x2_ASAP7_75t_L g411 ( .A(n_251), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g278 ( .A(n_252), .B(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g283 ( .A(n_252), .Y(n_283) );
BUFx2_ASAP7_75t_L g351 ( .A(n_252), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_261), .B(n_285), .Y(n_284) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_261), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g344 ( .A(n_261), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_262), .B(n_278), .Y(n_409) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g352 ( .A(n_267), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_271), .Y(n_305) );
AND2x4_ASAP7_75t_L g315 ( .A(n_271), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g402 ( .A(n_271), .Y(n_402) );
INVx2_ASAP7_75t_L g423 ( .A(n_271), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_277), .A2(n_436), .B1(n_438), .B2(n_439), .Y(n_435) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g347 ( .A(n_278), .B(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g301 ( .A(n_279), .B(n_285), .Y(n_301) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x4_ASAP7_75t_L g290 ( .A(n_282), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g412 ( .A(n_282), .Y(n_412) );
INVx2_ASAP7_75t_L g298 ( .A(n_283), .Y(n_298) );
AND2x2_ASAP7_75t_L g326 ( .A(n_283), .B(n_285), .Y(n_326) );
INVx3_ASAP7_75t_L g334 ( .A(n_283), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_283), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g319 ( .A(n_284), .Y(n_319) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g335 ( .A(n_286), .Y(n_335) );
OAI222xp33_ASAP7_75t_L g458 ( .A1(n_288), .A2(n_448), .B1(n_459), .B2(n_462), .C1(n_464), .C2(n_466), .Y(n_458) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g399 ( .A(n_290), .Y(n_399) );
AND2x2_ASAP7_75t_L g463 ( .A(n_290), .B(n_333), .Y(n_463) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_293), .B(n_384), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_302), .B1(n_310), .B2(n_312), .C(n_317), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g385 ( .A(n_298), .Y(n_385) );
INVx2_ASAP7_75t_L g447 ( .A(n_299), .Y(n_447) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx2_ASAP7_75t_L g348 ( .A(n_300), .Y(n_348) );
AND2x2_ASAP7_75t_L g384 ( .A(n_300), .B(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g350 ( .A(n_301), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g376 ( .A(n_301), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g465 ( .A(n_301), .Y(n_465) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g414 ( .A(n_305), .Y(n_414) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g437 ( .A(n_307), .B(n_315), .Y(n_437) );
AND2x2_ASAP7_75t_L g460 ( .A(n_307), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g321 ( .A(n_309), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g456 ( .A(n_309), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_310), .A2(n_364), .B1(n_398), .B2(n_400), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g425 ( .A1(n_310), .A2(n_426), .B(n_429), .Y(n_425) );
INVxp67_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
INVx2_ASAP7_75t_SL g446 ( .A(n_311), .Y(n_446) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
OR2x2_ASAP7_75t_L g359 ( .A(n_313), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g457 ( .A(n_313), .B(n_456), .Y(n_457) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g330 ( .A(n_315), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_315), .B(n_339), .Y(n_355) );
INVx2_ASAP7_75t_L g382 ( .A(n_315), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B1(n_323), .B2(n_325), .Y(n_317) );
NOR2xp33_ASAP7_75t_SL g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_319), .A2(n_393), .B1(n_406), .B2(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g415 ( .A(n_324), .B(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_332), .B(n_336), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g396 ( .A(n_329), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_329), .B(n_379), .Y(n_407) );
INVx1_ASAP7_75t_L g365 ( .A(n_331), .Y(n_365) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_333), .B(n_346), .Y(n_438) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI21xp33_ASAP7_75t_L g451 ( .A1(n_334), .A2(n_452), .B(n_454), .Y(n_451) );
OAI21xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_341), .B(n_349), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_L g395 ( .A(n_340), .Y(n_395) );
INVx1_ASAP7_75t_L g461 ( .A(n_340), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_L g434 ( .A(n_344), .Y(n_434) );
OR2x2_ASAP7_75t_L g445 ( .A(n_345), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND3xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .C(n_354), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_350), .A2(n_411), .B1(n_413), .B2(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g377 ( .A(n_351), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_352), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_355), .B(n_359), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g417 ( .A1(n_355), .A2(n_418), .B1(n_421), .B2(n_424), .C(n_425), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_361), .B(n_362), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g366 ( .A(n_360), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_368), .B2(n_860), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AND2x4_ASAP7_75t_L g449 ( .A(n_371), .B(n_427), .Y(n_449) );
NAND4xp25_ASAP7_75t_L g372 ( .A(n_373), .B(n_403), .C(n_430), .D(n_450), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_386), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_380), .B2(n_381), .C(n_383), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_376), .A2(n_433), .B1(n_455), .B2(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g429 ( .A(n_378), .Y(n_429) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g413 ( .A(n_379), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_379), .B(n_422), .Y(n_421) );
NAND2x1_ASAP7_75t_L g466 ( .A(n_379), .B(n_467), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_381), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g388 ( .A(n_385), .B(n_389), .Y(n_388) );
OAI21xp33_ASAP7_75t_SL g386 ( .A1(n_387), .A2(n_392), .B(n_397), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g416 ( .A(n_402), .Y(n_416) );
AOI211xp5_ASAP7_75t_L g430 ( .A1(n_402), .A2(n_431), .B(n_435), .C(n_441), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_417), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_405), .B(n_410), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g464 ( .A(n_412), .B(n_465), .Y(n_464) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx3_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp33_ASAP7_75t_R g441 ( .A1(n_442), .A2(n_445), .B1(n_447), .B2(n_448), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g455 ( .A(n_444), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_458), .Y(n_450) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_471), .B(n_811), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_472), .A2(n_473), .B1(n_834), .B2(n_835), .Y(n_833) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_473), .A2(n_812), .B(n_813), .Y(n_811) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_699), .Y(n_473) );
NOR4xp75_ASAP7_75t_L g474 ( .A(n_475), .B(n_638), .C(n_662), .D(n_681), .Y(n_474) );
NAND3x1_ASAP7_75t_L g475 ( .A(n_476), .B(n_579), .C(n_629), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_522), .B1(n_559), .B2(n_575), .Y(n_476) );
AND2x2_ASAP7_75t_L g760 ( .A(n_477), .B(n_635), .Y(n_760) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_494), .Y(n_477) );
AND2x2_ASAP7_75t_L g710 ( .A(n_478), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_478), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g737 ( .A(n_478), .Y(n_737) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g583 ( .A(n_479), .Y(n_583) );
INVx2_ASAP7_75t_L g604 ( .A(n_479), .Y(n_604) );
AND2x2_ASAP7_75t_L g698 ( .A(n_479), .B(n_661), .Y(n_698) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g578 ( .A(n_480), .Y(n_578) );
AND2x2_ASAP7_75t_L g677 ( .A(n_480), .B(n_590), .Y(n_677) );
AOI21x1_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_482), .B(n_492), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_488), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_486), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_486), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_486), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_486), .A2(n_597), .B(n_598), .Y(n_596) );
BUFx4f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g630 ( .A(n_494), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g745 ( .A(n_494), .Y(n_745) );
AND2x2_ASAP7_75t_L g751 ( .A(n_494), .B(n_615), .Y(n_751) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_509), .Y(n_494) );
INVx1_ASAP7_75t_L g588 ( .A(n_495), .Y(n_588) );
INVx4_ASAP7_75t_L g608 ( .A(n_495), .Y(n_608) );
OR2x2_ASAP7_75t_L g657 ( .A(n_495), .B(n_637), .Y(n_657) );
BUFx2_ASAP7_75t_L g726 ( .A(n_495), .Y(n_726) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
OAI21x1_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_501), .B(n_507), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_503), .A2(n_571), .B(n_572), .Y(n_570) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_508), .A2(n_513), .B(n_516), .Y(n_512) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_508), .A2(n_531), .B(n_534), .Y(n_530) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_508), .A2(n_542), .B(n_545), .Y(n_541) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_508), .A2(n_567), .B(n_570), .Y(n_566) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_508), .A2(n_593), .B(n_596), .Y(n_592) );
AND2x2_ASAP7_75t_L g577 ( .A(n_509), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g679 ( .A(n_509), .Y(n_679) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g603 ( .A(n_510), .Y(n_603) );
OAI21x1_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_521), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_511), .A2(n_566), .B(n_573), .Y(n_565) );
OAI21xp33_ASAP7_75t_SL g617 ( .A1(n_511), .A2(n_512), .B(n_521), .Y(n_617) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_511), .A2(n_566), .B(n_573), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_520), .Y(n_516) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2x1_ASAP7_75t_L g748 ( .A(n_524), .B(n_688), .Y(n_748) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_538), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g633 ( .A(n_526), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g653 ( .A(n_526), .B(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_526), .Y(n_687) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g643 ( .A(n_527), .B(n_540), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g798 ( .A(n_527), .B(n_539), .Y(n_798) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g720 ( .A(n_528), .Y(n_720) );
OAI21x1_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_537), .Y(n_528) );
OAI21x1_ASAP7_75t_L g540 ( .A1(n_529), .A2(n_541), .B(n_550), .Y(n_540) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_529), .A2(n_530), .B(n_537), .Y(n_563) );
OA21x2_ASAP7_75t_L g574 ( .A1(n_529), .A2(n_541), .B(n_550), .Y(n_574) );
INVx2_ASAP7_75t_L g741 ( .A(n_538), .Y(n_741) );
AND2x4_ASAP7_75t_L g779 ( .A(n_538), .B(n_718), .Y(n_779) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_551), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g619 ( .A(n_540), .Y(n_619) );
AND2x2_ASAP7_75t_L g654 ( .A(n_540), .B(n_552), .Y(n_654) );
AND2x2_ASAP7_75t_L g777 ( .A(n_540), .B(n_627), .Y(n_777) );
AND2x2_ASAP7_75t_L g788 ( .A(n_540), .B(n_565), .Y(n_788) );
AOI21x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_549), .Y(n_545) );
AND2x2_ASAP7_75t_L g646 ( .A(n_551), .B(n_563), .Y(n_646) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g562 ( .A(n_552), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g620 ( .A(n_552), .B(n_563), .Y(n_620) );
OR2x2_ASAP7_75t_L g634 ( .A(n_552), .B(n_574), .Y(n_634) );
AND2x2_ASAP7_75t_L g719 ( .A(n_552), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_552), .B(n_574), .Y(n_730) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_552), .Y(n_772) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g668 ( .A(n_562), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g775 ( .A(n_562), .B(n_776), .C(n_778), .Y(n_775) );
INVx1_ASAP7_75t_L g612 ( .A(n_563), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_564), .B(n_620), .Y(n_742) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_574), .Y(n_564) );
INVx1_ASAP7_75t_L g586 ( .A(n_565), .Y(n_586) );
AND2x2_ASAP7_75t_L g791 ( .A(n_574), .B(n_627), .Y(n_791) );
INVx1_ASAP7_75t_L g794 ( .A(n_575), .Y(n_794) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g773 ( .A(n_576), .B(n_606), .Y(n_773) );
OR2x2_ASAP7_75t_L g784 ( .A(n_576), .B(n_657), .Y(n_784) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g660 ( .A(n_577), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g808 ( .A(n_577), .B(n_587), .Y(n_808) );
AND2x2_ASAP7_75t_L g616 ( .A(n_578), .B(n_617), .Y(n_616) );
A2O1A1O1Ixp25_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_584), .B(n_600), .C(n_609), .D(n_613), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g694 ( .A(n_582), .B(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g631 ( .A(n_583), .Y(n_631) );
INVx1_ASAP7_75t_L g666 ( .A(n_584), .Y(n_666) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
AND2x2_ASAP7_75t_L g645 ( .A(n_585), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g636 ( .A(n_586), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g665 ( .A(n_587), .Y(n_665) );
AND2x2_ASAP7_75t_L g736 ( .A(n_587), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g782 ( .A(n_587), .B(n_616), .Y(n_782) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g607 ( .A(n_589), .Y(n_607) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_589), .Y(n_615) );
INVx2_ASAP7_75t_L g661 ( .A(n_589), .Y(n_661) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g637 ( .A(n_590), .Y(n_637) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B(n_599), .Y(n_590) );
INVx1_ASAP7_75t_L g732 ( .A(n_600), .Y(n_732) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_605), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g656 ( .A1(n_601), .A2(n_606), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
AND2x2_ASAP7_75t_L g622 ( .A(n_602), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g727 ( .A(n_602), .B(n_677), .Y(n_727) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g659 ( .A(n_603), .B(n_637), .Y(n_659) );
AND2x2_ASAP7_75t_L g683 ( .A(n_604), .B(n_608), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g767 ( .A(n_604), .B(n_623), .Y(n_767) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g711 ( .A(n_606), .Y(n_711) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx2_ASAP7_75t_L g623 ( .A(n_608), .Y(n_623) );
NAND2x1_ASAP7_75t_L g678 ( .A(n_608), .B(n_679), .Y(n_678) );
OAI32xp33_ASAP7_75t_L g799 ( .A1(n_609), .A2(n_675), .A3(n_783), .B1(n_800), .B2(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g673 ( .A(n_611), .Y(n_673) );
AND2x2_ASAP7_75t_L g696 ( .A(n_611), .B(n_654), .Y(n_696) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g693 ( .A(n_612), .B(n_627), .Y(n_693) );
OAI22xp33_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_618), .B1(n_621), .B2(n_624), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g650 ( .A(n_616), .B(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g669 ( .A(n_617), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_L g783 ( .A(n_619), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_620), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g762 ( .A(n_620), .Y(n_762) );
AND2x2_ASAP7_75t_L g790 ( .A(n_620), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_L g697 ( .A(n_622), .B(n_698), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_L g746 ( .A1(n_622), .A2(n_677), .B(n_747), .C(n_749), .Y(n_746) );
INVx1_ASAP7_75t_L g651 ( .A(n_623), .Y(n_651) );
AND2x2_ASAP7_75t_L g695 ( .A(n_623), .B(n_661), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_625), .B(n_646), .Y(n_664) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVxp67_ASAP7_75t_SL g642 ( .A(n_627), .Y(n_642) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_627), .Y(n_689) );
INVx1_ASAP7_75t_L g718 ( .A(n_627), .Y(n_718) );
BUFx3_ASAP7_75t_L g731 ( .A(n_627), .Y(n_731) );
INVx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .C(n_635), .Y(n_629) );
INVx1_ASAP7_75t_L g753 ( .A(n_630), .Y(n_753) );
OR2x2_ASAP7_75t_L g680 ( .A(n_631), .B(n_665), .Y(n_680) );
OR2x2_ASAP7_75t_L g644 ( .A(n_632), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_633), .A2(n_671), .B1(n_675), .B2(n_680), .Y(n_670) );
INVx2_ASAP7_75t_L g674 ( .A(n_634), .Y(n_674) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_634), .Y(n_686) );
INVx1_ASAP7_75t_L g705 ( .A(n_634), .Y(n_705) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVxp67_ASAP7_75t_L g649 ( .A(n_637), .Y(n_649) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_637), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_647), .B1(n_652), .B2(n_655), .Y(n_638) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_644), .Y(n_639) );
BUFx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_646), .Y(n_724) );
NAND2x1p5_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g715 ( .A(n_648), .Y(n_715) );
BUFx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI221x1_ASAP7_75t_L g701 ( .A1(n_650), .A2(n_702), .B1(n_706), .B2(n_708), .C(n_712), .Y(n_701) );
BUFx2_ASAP7_75t_L g804 ( .A(n_651), .Y(n_804) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_654), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_654), .B(n_731), .Y(n_756) );
AND2x2_ASAP7_75t_L g810 ( .A(n_654), .B(n_689), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .B(n_660), .Y(n_655) );
AOI211xp5_ASAP7_75t_L g792 ( .A1(n_657), .A2(n_793), .B(n_799), .C(n_802), .Y(n_792) );
OAI222xp33_ASAP7_75t_L g780 ( .A1(n_658), .A2(n_781), .B1(n_783), .B2(n_784), .C1(n_785), .C2(n_789), .Y(n_780) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AO21x1_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_669), .B(n_670), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_666), .B2(n_667), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g806 ( .A(n_669), .Y(n_806) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x4_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
AND2x2_ASAP7_75t_L g707 ( .A(n_674), .B(n_693), .Y(n_707) );
INVx1_ASAP7_75t_L g733 ( .A(n_674), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_675), .A2(n_729), .B1(n_732), .B2(n_733), .Y(n_728) );
INVx1_ASAP7_75t_L g759 ( .A(n_675), .Y(n_759) );
OR2x6_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx1_ASAP7_75t_L g805 ( .A(n_676), .Y(n_805) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g766 ( .A(n_679), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_679), .B(n_695), .Y(n_800) );
OAI21xp33_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_684), .B(n_690), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR3x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .C(n_688), .Y(n_685) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_694), .B1(n_696), .B2(n_697), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_693), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g778 ( .A(n_693), .Y(n_778) );
INVx2_ASAP7_75t_L g752 ( .A(n_696), .Y(n_752) );
INVx3_ASAP7_75t_L g713 ( .A(n_697), .Y(n_713) );
NOR2x1_ASAP7_75t_L g699 ( .A(n_700), .B(n_757), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_721), .C(n_746), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g769 ( .A(n_718), .Y(n_769) );
BUFx2_ASAP7_75t_L g740 ( .A(n_720), .Y(n_740) );
AOI211xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_725), .B(n_728), .C(n_734), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AND2x4_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
OR2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_731), .B(n_798), .Y(n_797) );
OAI22xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_738), .B1(n_742), .B2(n_743), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
AND2x2_ASAP7_75t_L g786 ( .A(n_739), .B(n_777), .Y(n_786) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g787 ( .A(n_740), .B(n_788), .Y(n_787) );
OR2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_749) );
INVx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVxp67_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_763), .C(n_792), .Y(n_757) );
OAI21xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_780), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_768), .B1(n_773), .B2(n_774), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
NOR2xp67_ASAP7_75t_L g774 ( .A(n_775), .B(n_779), .Y(n_774) );
INVx2_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NOR2xp33_ASAP7_75t_SL g785 ( .A(n_786), .B(n_787), .Y(n_785) );
INVx2_ASAP7_75t_L g801 ( .A(n_787), .Y(n_801) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AOI21xp33_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_807), .B(n_809), .Y(n_802) );
NAND3x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .C(n_806), .Y(n_803) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
INVx4_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
BUFx12f_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI21xp33_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_845), .B(n_852), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_826), .B(n_837), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx3_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx4_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
AND3x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .C(n_825), .Y(n_821) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g843 ( .A(n_823), .Y(n_843) );
AND2x6_ASAP7_75t_SL g841 ( .A(n_825), .B(n_842), .Y(n_841) );
XOR2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_833), .Y(n_826) );
INVx1_ASAP7_75t_L g832 ( .A(n_829), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_844), .Y(n_837) );
INVx4_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
CKINVDCx8_ASAP7_75t_R g840 ( .A(n_841), .Y(n_840) );
INVx3_ASAP7_75t_L g858 ( .A(n_841), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_846), .Y(n_845) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_847), .Y(n_846) );
INVx4_ASAP7_75t_SL g847 ( .A(n_848), .Y(n_847) );
BUFx3_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
OR2x4_ASAP7_75t_L g856 ( .A(n_850), .B(n_857), .Y(n_856) );
BUFx2_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
BUFx3_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
endmodule