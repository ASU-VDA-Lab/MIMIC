module fake_jpeg_28599_n_113 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_18),
.B1(n_38),
.B2(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_17),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_1),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_60),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_47),
.C(n_57),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_1),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_44),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_45),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_49),
.C(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_2),
.Y(n_81)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_9),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_70),
.A2(n_48),
.B1(n_45),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_10),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_81),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_41),
.B1(n_43),
.B2(n_40),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_19),
.B1(n_33),
.B2(n_32),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_64),
.B(n_68),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_84),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_2),
.B(n_3),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_83),
.B(n_12),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_4),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_86),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_91),
.B1(n_96),
.B2(n_94),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_95),
.B(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_14),
.C(n_15),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g97 ( 
.A(n_79),
.B(n_24),
.C(n_25),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_100),
.B1(n_95),
.B2(n_85),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_30),
.Y(n_99)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_97),
.C(n_90),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_91),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_105),
.B(n_89),
.Y(n_108)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_101),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_108),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_93),
.C(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_99),
.Y(n_113)
);


endmodule