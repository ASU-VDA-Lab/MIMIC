module fake_jpeg_14297_n_648 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_63),
.B(n_66),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_64),
.B(n_76),
.Y(n_134)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_22),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_16),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_77),
.B(n_51),
.Y(n_197)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_82),
.Y(n_216)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_85),
.Y(n_166)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_87),
.Y(n_169)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_89),
.Y(n_205)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_92),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_20),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_105),
.Y(n_138)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_95),
.Y(n_201)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_96),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_98),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_100),
.Y(n_212)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_103),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_43),
.B(n_16),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_104),
.B(n_106),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_19),
.B(n_0),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_19),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_1),
.Y(n_160)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_36),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_122),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_38),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_46),
.Y(n_123)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_29),
.Y(n_126)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

NAND2x1_ASAP7_75t_SL g195 ( 
.A(n_127),
.B(n_59),
.Y(n_195)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_30),
.Y(n_129)
);

BUFx4f_ASAP7_75t_SL g207 ( 
.A(n_129),
.Y(n_207)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_85),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_141),
.B(n_146),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_87),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_77),
.B(n_49),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_147),
.B(n_152),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_62),
.A2(n_40),
.B1(n_50),
.B2(n_32),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_150),
.A2(n_100),
.B1(n_119),
.B2(n_125),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_87),
.Y(n_152)
);

BUFx16f_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

BUFx8_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_94),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_158),
.B(n_159),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_94),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_160),
.B(n_173),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_107),
.B(n_54),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_189),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_84),
.B(n_54),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_99),
.B(n_26),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_176),
.B(n_186),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_78),
.B(n_49),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_98),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_81),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_202),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_89),
.A2(n_40),
.B1(n_50),
.B2(n_37),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_191),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_195),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_26),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_68),
.A2(n_30),
.B1(n_32),
.B2(n_37),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_198),
.A2(n_129),
.B1(n_127),
.B2(n_124),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_130),
.B(n_24),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_83),
.B(n_24),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_116),
.B(n_53),
.Y(n_202)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_70),
.Y(n_203)
);

INVx5_ASAP7_75t_SL g282 ( 
.A(n_203),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_121),
.B(n_53),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_210),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_82),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_55),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_217),
.B(n_240),
.Y(n_317)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_220),
.Y(n_296)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_222),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_L g339 ( 
.A1(n_223),
.A2(n_228),
.B(n_237),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_86),
.B1(n_128),
.B2(n_101),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_225),
.A2(n_229),
.B1(n_182),
.B2(n_211),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_144),
.B(n_161),
.C(n_177),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_227),
.B(n_244),
.C(n_290),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_131),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_230),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_231),
.Y(n_323)
);

AOI21xp33_ASAP7_75t_L g232 ( 
.A1(n_175),
.A2(n_51),
.B(n_55),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_232),
.B(n_264),
.Y(n_348)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_137),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_154),
.Y(n_234)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_171),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_236),
.B(n_243),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_134),
.Y(n_237)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_164),
.B(n_184),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_241),
.Y(n_325)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_148),
.Y(n_242)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_242),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_138),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_214),
.C(n_201),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_245),
.Y(n_326)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_246),
.Y(n_341)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_247),
.Y(n_293)
);

CKINVDCx9p33_ASAP7_75t_R g248 ( 
.A(n_169),
.Y(n_248)
);

INVx4_ASAP7_75t_SL g331 ( 
.A(n_248),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_137),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVx3_ASAP7_75t_SL g252 ( 
.A(n_203),
.Y(n_252)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_253),
.A2(n_135),
.B1(n_132),
.B2(n_211),
.Y(n_304)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

INVx8_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_145),
.Y(n_256)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_136),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_287),
.Y(n_301)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_145),
.Y(n_259)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_259),
.Y(n_347)
);

CKINVDCx12_ASAP7_75t_R g261 ( 
.A(n_153),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_261),
.Y(n_309)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_151),
.Y(n_262)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_262),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_140),
.B(n_41),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_183),
.Y(n_265)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_194),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_266),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_133),
.B(n_41),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_267),
.B(n_271),
.Y(n_312)
);

CKINVDCx9p33_ASAP7_75t_R g268 ( 
.A(n_187),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_268),
.Y(n_302)
);

CKINVDCx12_ASAP7_75t_R g269 ( 
.A(n_207),
.Y(n_269)
);

NAND2x1_ASAP7_75t_SL g298 ( 
.A(n_269),
.B(n_289),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_187),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_276),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_180),
.B(n_57),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_206),
.Y(n_272)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_151),
.Y(n_273)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_273),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_L g274 ( 
.A1(n_198),
.A2(n_79),
.B1(n_118),
.B2(n_117),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_278),
.B1(n_281),
.B2(n_165),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_139),
.B(n_39),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_275),
.B(n_279),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_195),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_207),
.A2(n_39),
.B(n_61),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_285),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_156),
.A2(n_40),
.B1(n_50),
.B2(n_103),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_139),
.B(n_57),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_157),
.B(n_60),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_280),
.B(n_165),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_156),
.A2(n_123),
.B1(n_114),
.B2(n_92),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_143),
.Y(n_283)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_283),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_155),
.B(n_61),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_284),
.B(n_288),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_174),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_167),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_291),
.Y(n_334)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_170),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_170),
.B(n_60),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_157),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_172),
.B(n_30),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_172),
.B(n_45),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_218),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_295),
.B(n_243),
.Y(n_355)
);

OA22x2_ASAP7_75t_L g379 ( 
.A1(n_299),
.A2(n_338),
.B1(n_331),
.B2(n_311),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_304),
.A2(n_335),
.B1(n_268),
.B2(n_229),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_224),
.A2(n_45),
.B(n_38),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_307),
.A2(n_328),
.B(n_333),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_319),
.A2(n_332),
.B1(n_282),
.B2(n_254),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_224),
.A2(n_135),
.B1(n_132),
.B2(n_216),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_320),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_322),
.B(n_270),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_274),
.A2(n_192),
.B(n_216),
.Y(n_328)
);

AND2x2_ASAP7_75t_SL g329 ( 
.A(n_240),
.B(n_174),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_329),
.B(n_330),
.C(n_290),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_227),
.B(n_178),
.C(n_162),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_292),
.A2(n_75),
.B1(n_182),
.B2(n_212),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_221),
.A2(n_59),
.B(n_47),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_280),
.A2(n_178),
.B1(n_212),
.B2(n_162),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_221),
.B(n_196),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_344),
.Y(n_356)
);

O2A1O1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_248),
.A2(n_179),
.B(n_174),
.C(n_192),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_228),
.A2(n_179),
.B(n_193),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_342),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_263),
.B(n_196),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_249),
.B(n_213),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_302),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_260),
.B(n_237),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_349),
.B(n_272),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_353),
.A2(n_363),
.B1(n_368),
.B2(n_376),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_354),
.B(n_360),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_355),
.B(n_357),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_294),
.B(n_255),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_358),
.Y(n_405)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_359),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_322),
.B(n_317),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_362),
.B(n_370),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_299),
.A2(n_219),
.B1(n_226),
.B2(n_244),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_332),
.A2(n_252),
.B1(n_282),
.B2(n_239),
.Y(n_364)
);

OAI22x1_ASAP7_75t_L g419 ( 
.A1(n_364),
.A2(n_385),
.B1(n_311),
.B2(n_318),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_234),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_365),
.B(n_369),
.Y(n_436)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_296),
.Y(n_366)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_366),
.Y(n_425)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_367),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_337),
.A2(n_304),
.B1(n_328),
.B2(n_314),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_312),
.B(n_230),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_317),
.B(n_250),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_217),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_371),
.A2(n_338),
.B(n_301),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_298),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_373),
.B(n_380),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_315),
.B(n_223),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_321),
.C(n_305),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_375),
.A2(n_381),
.B1(n_399),
.B2(n_323),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_335),
.A2(n_220),
.B1(n_167),
.B2(n_213),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_296),
.Y(n_377)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_377),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_333),
.A2(n_188),
.B1(n_289),
.B2(n_242),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_378),
.A2(n_387),
.B1(n_343),
.B2(n_324),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_298),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_329),
.A2(n_223),
.B1(n_290),
.B2(n_228),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_222),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_354),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_389),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_301),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_392),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g385 ( 
.A1(n_300),
.A2(n_256),
.B1(n_259),
.B2(n_262),
.Y(n_385)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_331),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_386),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_310),
.A2(n_315),
.B1(n_330),
.B2(n_320),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_388),
.B(n_246),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_327),
.B(n_241),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_346),
.B(n_287),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_308),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_394),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_301),
.Y(n_394)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_297),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_396),
.Y(n_422)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_341),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_308),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_398),
.Y(n_431)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_306),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_334),
.B(n_257),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_361),
.A2(n_342),
.B(n_307),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_401),
.A2(n_435),
.B(n_377),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_368),
.A2(n_329),
.B1(n_339),
.B2(n_350),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_402),
.A2(n_380),
.B(n_372),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_361),
.A2(n_362),
.B1(n_356),
.B2(n_382),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_406),
.A2(n_423),
.B1(n_424),
.B2(n_427),
.Y(n_450)
);

OAI32xp33_ASAP7_75t_L g408 ( 
.A1(n_356),
.A2(n_321),
.A3(n_336),
.B1(n_305),
.B2(n_325),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_413),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_415),
.C(n_420),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_325),
.C(n_336),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_417),
.B(n_394),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_419),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_343),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_391),
.A2(n_188),
.B1(n_233),
.B2(n_345),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_426),
.A2(n_428),
.B1(n_393),
.B2(n_397),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_391),
.A2(n_273),
.B1(n_251),
.B2(n_283),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_363),
.A2(n_313),
.B1(n_347),
.B2(n_352),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_303),
.C(n_323),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_429),
.B(n_430),
.C(n_434),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_370),
.B(n_352),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_373),
.A2(n_326),
.B(n_318),
.Y(n_435)
);

OA22x2_ASAP7_75t_L g438 ( 
.A1(n_375),
.A2(n_347),
.B1(n_313),
.B2(n_293),
.Y(n_438)
);

OA22x2_ASAP7_75t_L g455 ( 
.A1(n_438),
.A2(n_353),
.B1(n_379),
.B2(n_384),
.Y(n_455)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_440),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_455),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_425),
.Y(n_442)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_432),
.Y(n_443)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_443),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g444 ( 
.A1(n_407),
.A2(n_378),
.B(n_379),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_444),
.B(n_438),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_431),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_460),
.Y(n_475)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_432),
.Y(n_446)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_446),
.Y(n_499)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_433),
.Y(n_447)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_448),
.A2(n_451),
.B1(n_468),
.B2(n_470),
.Y(n_498)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_433),
.Y(n_449)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_449),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_414),
.A2(n_372),
.B1(n_360),
.B2(n_381),
.Y(n_451)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_453),
.Y(n_506)
);

OAI21xp33_ASAP7_75t_L g491 ( 
.A1(n_456),
.A2(n_471),
.B(n_466),
.Y(n_491)
);

FAx1_ASAP7_75t_SL g457 ( 
.A(n_437),
.B(n_371),
.CI(n_366),
.CON(n_457),
.SN(n_457)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_467),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_459),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_396),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_408),
.B(n_390),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_464),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_411),
.B(n_371),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_462),
.B(n_463),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_412),
.B(n_436),
.Y(n_463)
);

OAI32xp33_ASAP7_75t_L g464 ( 
.A1(n_418),
.A2(n_379),
.A3(n_376),
.B1(n_293),
.B2(n_340),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_422),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_466),
.Y(n_484)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_412),
.B(n_359),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_414),
.A2(n_395),
.B1(n_398),
.B2(n_358),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_434),
.B(n_326),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_471),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_407),
.A2(n_297),
.B1(n_316),
.B2(n_286),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_403),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_405),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_421),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_426),
.A2(n_316),
.B1(n_265),
.B2(n_266),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_473),
.A2(n_427),
.B1(n_423),
.B2(n_438),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_400),
.B(n_340),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_421),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_420),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_477),
.B(n_489),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_430),
.C(n_429),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_478),
.B(n_497),
.C(n_448),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_461),
.A2(n_418),
.B1(n_402),
.B2(n_406),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_482),
.A2(n_492),
.B1(n_451),
.B2(n_502),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_460),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_486),
.B(n_488),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_459),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_409),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_491),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_439),
.A2(n_428),
.B1(n_401),
.B2(n_404),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_441),
.B(n_435),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_493),
.B(n_508),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_454),
.B(n_415),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_494),
.B(n_502),
.Y(n_531)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_495),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_496),
.B(n_504),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_413),
.C(n_417),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_439),
.B(n_416),
.Y(n_502)
);

NOR3xp33_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_367),
.C(n_419),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_457),
.B(n_416),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_505),
.B(n_473),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_507),
.A2(n_450),
.B1(n_452),
.B2(n_442),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_SL g509 ( 
.A(n_484),
.B(n_465),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_509),
.B(n_517),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_510),
.A2(n_538),
.B1(n_507),
.B2(n_500),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_475),
.B(n_445),
.Y(n_512)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_512),
.Y(n_547)
);

MAJx2_ASAP7_75t_L g554 ( 
.A(n_513),
.B(n_258),
.C(n_238),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_514),
.A2(n_521),
.B1(n_534),
.B2(n_483),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_450),
.C(n_468),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_515),
.B(n_519),
.C(n_525),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_484),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_501),
.A2(n_493),
.B(n_483),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_518),
.A2(n_536),
.B(n_524),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_477),
.B(n_444),
.C(n_449),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_495),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_520),
.B(n_523),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_480),
.A2(n_444),
.B1(n_464),
.B2(n_455),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_475),
.Y(n_522)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_522),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_482),
.B(n_440),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_478),
.B(n_447),
.C(n_455),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_453),
.Y(n_526)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_526),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_489),
.B(n_455),
.C(n_472),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_527),
.B(n_529),
.C(n_537),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_446),
.C(n_443),
.Y(n_529)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_530),
.Y(n_562)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_533),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_480),
.A2(n_470),
.B1(n_438),
.B2(n_386),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_285),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_535),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_485),
.B(n_483),
.C(n_493),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_508),
.A2(n_386),
.B1(n_247),
.B2(n_245),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_476),
.A2(n_367),
.B1(n_37),
.B2(n_59),
.Y(n_539)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_539),
.Y(n_556)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_540),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_521),
.A2(n_501),
.B1(n_498),
.B2(n_487),
.Y(n_541)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_541),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_512),
.B(n_506),
.Y(n_543)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_543),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_490),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_544),
.B(n_529),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_526),
.B(n_503),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_546),
.B(n_522),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_531),
.B(n_498),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g581 ( 
.A(n_550),
.B(n_559),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_552),
.A2(n_555),
.B1(n_3),
.B2(n_5),
.Y(n_585)
);

OAI21xp33_ASAP7_75t_L g553 ( 
.A1(n_528),
.A2(n_499),
.B(n_479),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_553),
.B(n_561),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_554),
.B(n_563),
.C(n_215),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_534),
.A2(n_266),
.B1(n_215),
.B2(n_193),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_558),
.A2(n_525),
.B(n_519),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_531),
.B(n_238),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_511),
.B(n_235),
.Y(n_561)
);

XOR2x1_ASAP7_75t_L g563 ( 
.A(n_537),
.B(n_238),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_516),
.A2(n_215),
.B1(n_193),
.B2(n_136),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_565),
.Y(n_576)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_566),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_547),
.A2(n_518),
.B(n_536),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_567),
.A2(n_570),
.B(n_577),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_552),
.A2(n_515),
.B1(n_536),
.B2(n_527),
.Y(n_569)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_569),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_572),
.B(n_583),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_562),
.A2(n_513),
.B1(n_533),
.B2(n_510),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_573),
.B(n_540),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_558),
.A2(n_538),
.B(n_511),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_578),
.B(n_579),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_542),
.B(n_2),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_548),
.A2(n_136),
.B(n_3),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_580),
.A2(n_5),
.B(n_6),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_543),
.B(n_2),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_582),
.B(n_545),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_564),
.B(n_2),
.C(n_3),
.Y(n_583)
);

INVx13_ASAP7_75t_L g584 ( 
.A(n_545),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_584),
.A2(n_585),
.B1(n_556),
.B2(n_563),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g586 ( 
.A(n_546),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_586),
.B(n_551),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_568),
.A2(n_557),
.B1(n_556),
.B2(n_549),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_587),
.B(n_590),
.Y(n_605)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_588),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_577),
.B(n_564),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_592),
.B(n_595),
.Y(n_609)
);

FAx1_ASAP7_75t_SL g593 ( 
.A(n_566),
.B(n_560),
.CI(n_559),
.CON(n_593),
.SN(n_593)
);

BUFx24_ASAP7_75t_SL g619 ( 
.A(n_593),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_573),
.B(n_560),
.C(n_550),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_598),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_569),
.B(n_561),
.C(n_554),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_599),
.B(n_601),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_568),
.A2(n_541),
.B1(n_565),
.B2(n_7),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_600),
.B(n_580),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_586),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_602),
.B(n_582),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_SL g604 ( 
.A1(n_572),
.A2(n_583),
.B(n_578),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_604),
.A2(n_570),
.B(n_571),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_606),
.A2(n_599),
.B(n_593),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_607),
.B(n_576),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_597),
.B(n_575),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_611),
.B(n_612),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_603),
.B(n_574),
.C(n_581),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_595),
.B(n_574),
.C(n_571),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_613),
.B(n_614),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_592),
.B(n_596),
.C(n_594),
.Y(n_614)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_615),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_594),
.B(n_581),
.C(n_567),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_617),
.B(n_618),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_591),
.B(n_579),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g620 ( 
.A(n_610),
.B(n_575),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_620),
.B(n_629),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_622),
.B(n_627),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_616),
.A2(n_598),
.B1(n_600),
.B2(n_576),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_623),
.B(n_626),
.Y(n_637)
);

OAI21xp5_ASAP7_75t_SL g626 ( 
.A1(n_609),
.A2(n_584),
.B(n_589),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_SL g627 ( 
.A1(n_619),
.A2(n_589),
.B(n_590),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_614),
.A2(n_584),
.B(n_576),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_630),
.B(n_617),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_632),
.B(n_633),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_625),
.B(n_608),
.C(n_612),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_628),
.B(n_605),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_635),
.A2(n_636),
.B(n_5),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_621),
.B(n_607),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_631),
.A2(n_628),
.B(n_624),
.Y(n_639)
);

INVxp33_ASAP7_75t_L g642 ( 
.A(n_639),
.Y(n_642)
);

AOI21x1_ASAP7_75t_L g640 ( 
.A1(n_637),
.A2(n_629),
.B(n_9),
.Y(n_640)
);

AOI322xp5_ASAP7_75t_L g643 ( 
.A1(n_640),
.A2(n_641),
.A3(n_635),
.B1(n_11),
.B2(n_12),
.C1(n_14),
.C2(n_15),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_643),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_642),
.B(n_638),
.Y(n_645)
);

OAI221xp5_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_634),
.B1(n_11),
.B2(n_15),
.C(n_9),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_11),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_647),
.Y(n_648)
);


endmodule