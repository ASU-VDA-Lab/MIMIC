module fake_jpeg_12395_n_173 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVxp33_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_3),
.B(n_10),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx5_ASAP7_75t_SL g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

NAND2x1_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_35),
.Y(n_76)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_43),
.Y(n_70)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_45),
.B(n_46),
.Y(n_55)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_11),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_50),
.Y(n_58)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_52),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_69),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_67),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_18),
.B1(n_32),
.B2(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_65),
.B1(n_22),
.B2(n_17),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_18),
.B1(n_20),
.B2(n_13),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_20),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_75),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_16),
.B1(n_26),
.B2(n_22),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_74),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_14),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_38),
.B(n_28),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_7),
.C(n_8),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_89),
.B1(n_68),
.B2(n_64),
.Y(n_116)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_90),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_33),
.B(n_4),
.C(n_5),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_98),
.Y(n_115)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_92),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_97),
.Y(n_114)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_56),
.A2(n_60),
.B(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_72),
.Y(n_118)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_105),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_8),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_55),
.B1(n_65),
.B2(n_78),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_123),
.B1(n_103),
.B2(n_77),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_118),
.Y(n_133)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_79),
.C(n_57),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_111),
.C(n_104),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_57),
.C(n_68),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_98),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_64),
.B1(n_77),
.B2(n_73),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_84),
.B(n_87),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_115),
.B(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_105),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_128),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_123),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_139),
.B(n_122),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_131),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_85),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_128),
.C(n_111),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_83),
.B1(n_89),
.B2(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_137),
.A2(n_108),
.B1(n_117),
.B2(n_106),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_73),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_134),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_139),
.C(n_129),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_146),
.A2(n_132),
.B(n_109),
.C(n_138),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_125),
.B(n_124),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_126),
.B(n_136),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_133),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_149),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_150),
.B(n_151),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_142),
.C(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_162),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_144),
.C(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_160),
.B(n_161),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_102),
.B1(n_8),
.B2(n_100),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_153),
.B(n_150),
.C(n_143),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_117),
.B1(n_124),
.B2(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_110),
.C(n_137),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_167),
.B(n_168),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_163),
.C(n_169),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_167),
.Y(n_173)
);


endmodule