module fake_jpeg_3441_n_120 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_48),
.Y(n_50)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_32),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_40),
.B1(n_37),
.B2(n_38),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_57),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_4),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_51),
.C(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_80),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_41),
.C(n_18),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_1),
.B(n_3),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_79),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_3),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_92),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_5),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_6),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_6),
.B1(n_29),
.B2(n_9),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_103),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_8),
.C(n_10),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_19),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_11),
.B1(n_13),
.B2(n_16),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_102),
.B(n_17),
.Y(n_104)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_106),
.B1(n_100),
.B2(n_101),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_85),
.B(n_84),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_85),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_109),
.C(n_104),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_107),
.C(n_95),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_114),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_110),
.B(n_22),
.Y(n_116)
);

OAI31xp33_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_20),
.A3(n_24),
.B(n_25),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_26),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_27),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_28),
.Y(n_120)
);


endmodule