module fake_netlist_6_2758_n_3795 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_741, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_746, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3795);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_746;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3795;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1234;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1674;
wire n_1199;
wire n_3392;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_3152;
wire n_3579;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_3741;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_1009;
wire n_2405;
wire n_3706;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_1285;
wire n_873;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1772;
wire n_1232;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3316;
wire n_2212;
wire n_758;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_1798;
wire n_943;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_1094;
wire n_953;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_1088;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_3368;
wire n_917;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_1446;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_813;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_3732;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_3716;
wire n_1873;
wire n_905;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_3168;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_3247;
wire n_871;
wire n_3069;
wire n_922;
wire n_1760;
wire n_1335;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_2008;
wire n_2749;
wire n_3346;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3298;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_780;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_1214;
wire n_1801;
wire n_850;
wire n_1886;
wire n_928;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_3785;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_890;
wire n_2377;
wire n_2178;
wire n_3271;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_3500;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_3545;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_1634;
wire n_2078;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3431;
wire n_3209;
wire n_3450;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_963;
wire n_794;
wire n_2767;
wire n_3793;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1714;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_791;
wire n_1913;
wire n_3608;
wire n_837;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_2134;
wire n_1176;
wire n_1004;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_1817;
wire n_926;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_2231;
wire n_3609;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_3656;
wire n_2127;
wire n_1178;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_2424;
wire n_1604;
wire n_2296;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1398;
wire n_1048;
wire n_884;
wire n_1201;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_931;
wire n_1021;
wire n_3393;
wire n_811;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_1250;
wire n_958;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2323;
wire n_1220;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_2990;
wire n_1773;
wire n_1775;
wire n_1286;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3364;
wire n_3323;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3425;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_773;
wire n_3547;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_906;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3250;
wire n_3113;
wire n_3194;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_1847;
wire n_2052;
wire n_3634;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1397;
wire n_1037;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_3475;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3262;
wire n_3544;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_1406;
wire n_3790;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_806;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_1931;
wire n_2083;
wire n_1269;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_2128;
wire n_1650;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1325;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2888;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2923;
wire n_1804;
wire n_3711;
wire n_3776;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_3511;
wire n_2054;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_841;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1882;
wire n_1023;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_933;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_969;
wire n_2140;
wire n_988;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_769;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_3652;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_1408;
wire n_3567;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_863;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_1848;
wire n_1785;
wire n_1114;
wire n_763;
wire n_1147;
wire n_3268;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_957;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_3739;
wire n_2284;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_761;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3336;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_908;
wire n_2721;
wire n_2649;
wire n_944;
wire n_3556;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_2444;
wire n_839;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_779;
wire n_2205;
wire n_3699;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_829;
wire n_1156;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_859;
wire n_2033;
wire n_3086;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_3478;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_2221;
wire n_1170;
wire n_1819;
wire n_2055;
wire n_1260;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_2553;
wire n_1040;
wire n_915;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_3527;
wire n_2512;
wire n_3433;
wire n_1365;
wire n_1417;
wire n_2185;
wire n_2086;
wire n_1242;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_3504;
wire n_1449;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_341),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_7),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_687),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_16),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_116),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_528),
.Y(n_763)
);

BUFx8_ASAP7_75t_SL g764 ( 
.A(n_383),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_220),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_150),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_310),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_670),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_124),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_333),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_661),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_640),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_560),
.Y(n_773)
);

BUFx10_ASAP7_75t_L g774 ( 
.A(n_653),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_579),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_753),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_736),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_330),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_428),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_526),
.Y(n_780)
);

BUFx10_ASAP7_75t_L g781 ( 
.A(n_286),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_137),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_523),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_261),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_12),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_541),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_433),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_643),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_301),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_264),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_296),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_230),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_395),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_159),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_19),
.Y(n_795)
);

CKINVDCx14_ASAP7_75t_R g796 ( 
.A(n_248),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_461),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_704),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_559),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_702),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_259),
.Y(n_801)
);

CKINVDCx16_ASAP7_75t_R g802 ( 
.A(n_680),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_751),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_741),
.Y(n_804)
);

BUFx10_ASAP7_75t_L g805 ( 
.A(n_440),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_717),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_96),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_733),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_703),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_144),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_346),
.Y(n_811)
);

BUFx5_ASAP7_75t_L g812 ( 
.A(n_234),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_474),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_44),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_262),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_376),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_188),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_522),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_628),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_153),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_241),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_469),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_20),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_343),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_706),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_49),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_100),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_615),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_440),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_11),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_333),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_712),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_295),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_688),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_364),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_686),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_49),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_455),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_43),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_326),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_207),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_410),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_320),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_72),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_413),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_67),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_268),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_127),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_705),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_735),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_655),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_99),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_662),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_677),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_166),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_32),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_245),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_354),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_584),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_533),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_728),
.Y(n_861)
);

CKINVDCx16_ASAP7_75t_R g862 ( 
.A(n_343),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_361),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_611),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_241),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_349),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_125),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_88),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_707),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_624),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_726),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_701),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_389),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_303),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_721),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_469),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_499),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_539),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_148),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_156),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_376),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_12),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_3),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_597),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_421),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_320),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_262),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_125),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_757),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_342),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_247),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_671),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_386),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_327),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_593),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_393),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_711),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_166),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_738),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_668),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_454),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_642),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_245),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_534),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_617),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_211),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_734),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_310),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_384),
.Y(n_909)
);

BUFx2_ASAP7_75t_L g910 ( 
.A(n_404),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_744),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_138),
.Y(n_912)
);

CKINVDCx16_ASAP7_75t_R g913 ( 
.A(n_198),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_740),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_77),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_537),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_118),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_169),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_60),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_453),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_426),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_651),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_566),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_527),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_117),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_435),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_91),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_164),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_525),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_279),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_658),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_256),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_501),
.Y(n_933)
);

CKINVDCx16_ASAP7_75t_R g934 ( 
.A(n_732),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_532),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_454),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_218),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_380),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_510),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_404),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_134),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_380),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_417),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_323),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_531),
.Y(n_945)
);

BUFx5_ASAP7_75t_L g946 ( 
.A(n_718),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_693),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_729),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_283),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_261),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_339),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_87),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_375),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_240),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_654),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_229),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_284),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_511),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_120),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_194),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_109),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_441),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_102),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_524),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_109),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_209),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_107),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_207),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_722),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_251),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_568),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_17),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_44),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_472),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_117),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_632),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_131),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_644),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_752),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_564),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_126),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_322),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_453),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_30),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_549),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_439),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_192),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_124),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_192),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_673),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_299),
.B(n_89),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_221),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_567),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_723),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_431),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_562),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_268),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_672),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_258),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_209),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_212),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_147),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_487),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_421),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_554),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_332),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_477),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_163),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_517),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_719),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_378),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_94),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_15),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_275),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_535),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_692),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_392),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_198),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_73),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_621),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_739),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_518),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_163),
.Y(n_1023)
);

CKINVDCx14_ASAP7_75t_R g1024 ( 
.A(n_428),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_126),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_294),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_33),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_669),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_676),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_121),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_684),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_382),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_87),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_236),
.Y(n_1034)
);

INVxp67_ASAP7_75t_L g1035 ( 
.A(n_167),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_683),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_55),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_78),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_609),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_162),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_76),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_382),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_296),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_750),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_386),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_517),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_540),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_40),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_438),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_171),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_698),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_183),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_636),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_334),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_300),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_152),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_108),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_590),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_558),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_731),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_322),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_266),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_737),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_252),
.Y(n_1064)
);

BUFx10_ASAP7_75t_L g1065 ( 
.A(n_284),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_25),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_2),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_119),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_345),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_697),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_283),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_197),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_161),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_682),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_177),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_696),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_38),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_347),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_544),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_227),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_420),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_304),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_145),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_227),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_689),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_512),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_64),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_545),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_370),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_432),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_580),
.Y(n_1091)
);

INVx2_ASAP7_75t_SL g1092 ( 
.A(n_15),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_111),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_727),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_366),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_483),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_486),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_623),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_397),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_544),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_208),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_492),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_348),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_121),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_172),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_713),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_200),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_199),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_495),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_107),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_699),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_242),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_674),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_219),
.Y(n_1115)
);

BUFx10_ASAP7_75t_L g1116 ( 
.A(n_316),
.Y(n_1116)
);

INVxp67_ASAP7_75t_L g1117 ( 
.A(n_223),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_749),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_302),
.Y(n_1119)
);

CKINVDCx16_ASAP7_75t_R g1120 ( 
.A(n_754),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_208),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_487),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_582),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_652),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_565),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_156),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_488),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_9),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_171),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_552),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_690),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_530),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_311),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_110),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_714),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_657),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_52),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_2),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_503),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_220),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_234),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_197),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_69),
.Y(n_1143)
);

CKINVDCx16_ASAP7_75t_R g1144 ( 
.A(n_519),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_256),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_200),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_708),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_595),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_242),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_38),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_143),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_548),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_709),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_128),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_452),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_144),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_56),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_631),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_746),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_108),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_142),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_691),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_244),
.Y(n_1163)
);

CKINVDCx16_ASAP7_75t_R g1164 ( 
.A(n_513),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_470),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_492),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_159),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_292),
.Y(n_1168)
);

BUFx10_ASAP7_75t_L g1169 ( 
.A(n_538),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_436),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_285),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_319),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_457),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_55),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_259),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_725),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_641),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_439),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_493),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_634),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_74),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_539),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_236),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_418),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_321),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_358),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_360),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_131),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_161),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_383),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_418),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_347),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_604),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_240),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_747),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_267),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_346),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_271),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_260),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_80),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_334),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_720),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_232),
.Y(n_1203)
);

CKINVDCx16_ASAP7_75t_R g1204 ( 
.A(n_546),
.Y(n_1204)
);

CKINVDCx14_ASAP7_75t_R g1205 ( 
.A(n_408),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_536),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_120),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_141),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_43),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_187),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_323),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_330),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_228),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_685),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_575),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_681),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_294),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_529),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_83),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_28),
.Y(n_1220)
);

BUFx8_ASAP7_75t_SL g1221 ( 
.A(n_361),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_424),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_327),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_490),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_369),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_547),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_756),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_679),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_179),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_384),
.Y(n_1230)
);

CKINVDCx14_ASAP7_75t_R g1231 ( 
.A(n_152),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_182),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_645),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_98),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_136),
.Y(n_1235)
);

BUFx10_ASAP7_75t_L g1236 ( 
.A(n_287),
.Y(n_1236)
);

CKINVDCx20_ASAP7_75t_R g1237 ( 
.A(n_111),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_195),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_656),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_273),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_412),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_542),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_675),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_573),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_210),
.Y(n_1245)
);

CKINVDCx16_ASAP7_75t_R g1246 ( 
.A(n_205),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_90),
.Y(n_1247)
);

BUFx8_ASAP7_75t_SL g1248 ( 
.A(n_33),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_6),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_716),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_743),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_84),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_150),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_494),
.Y(n_1254)
);

BUFx8_ASAP7_75t_SL g1255 ( 
.A(n_700),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_710),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_35),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_305),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_665),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_56),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_508),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_478),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_715),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_397),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_145),
.Y(n_1265)
);

CKINVDCx14_ASAP7_75t_R g1266 ( 
.A(n_214),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_47),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_7),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_378),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_157),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_430),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_592),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_471),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_664),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_594),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_246),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_24),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_724),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_667),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_730),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_424),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_528),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_695),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_342),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_666),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_37),
.Y(n_1286)
);

BUFx8_ASAP7_75t_SL g1287 ( 
.A(n_694),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_225),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_357),
.Y(n_1289)
);

CKINVDCx16_ASAP7_75t_R g1290 ( 
.A(n_678),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_543),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_742),
.Y(n_1292)
);

INVxp67_ASAP7_75t_SL g1293 ( 
.A(n_893),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_812),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_812),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_812),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_812),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_812),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_893),
.Y(n_1299)
);

CKINVDCx14_ASAP7_75t_R g1300 ( 
.A(n_796),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_812),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_764),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_812),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_820),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_764),
.Y(n_1305)
);

INVxp33_ASAP7_75t_SL g1306 ( 
.A(n_846),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1221),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_820),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_894),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1221),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_894),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_832),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_903),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_903),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_835),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_941),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_941),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_954),
.Y(n_1318)
);

INVxp33_ASAP7_75t_SL g1319 ( 
.A(n_1155),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_954),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1183),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1183),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1240),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1240),
.Y(n_1324)
);

CKINVDCx16_ASAP7_75t_R g1325 ( 
.A(n_862),
.Y(n_1325)
);

INVxp33_ASAP7_75t_SL g1326 ( 
.A(n_991),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_760),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_835),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1248),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_832),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_835),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_835),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_839),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_839),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_839),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_839),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_865),
.Y(n_1337)
);

CKINVDCx14_ASAP7_75t_R g1338 ( 
.A(n_796),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_865),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_822),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_865),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_865),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_896),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_896),
.Y(n_1344)
);

INVxp33_ASAP7_75t_SL g1345 ( 
.A(n_991),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_896),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_896),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_986),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_986),
.Y(n_1349)
);

INVxp67_ASAP7_75t_L g1350 ( 
.A(n_910),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_986),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_986),
.Y(n_1352)
);

NOR2xp67_ASAP7_75t_L g1353 ( 
.A(n_789),
.B(n_0),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1248),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1007),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1007),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1007),
.Y(n_1357)
);

INVxp33_ASAP7_75t_SL g1358 ( 
.A(n_925),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_768),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1007),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_773),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1030),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1030),
.Y(n_1363)
);

INVxp33_ASAP7_75t_SL g1364 ( 
.A(n_1157),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_772),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1030),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1030),
.Y(n_1367)
);

INVxp33_ASAP7_75t_SL g1368 ( 
.A(n_1165),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1040),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1040),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1040),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1040),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1071),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1071),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1071),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1191),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_767),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1071),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1113),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1113),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1113),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1113),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_763),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_778),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_775),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_780),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_776),
.Y(n_1387)
);

INVxp67_ASAP7_75t_SL g1388 ( 
.A(n_767),
.Y(n_1388)
);

INVxp33_ASAP7_75t_L g1389 ( 
.A(n_770),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_770),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_799),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_800),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_791),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_792),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_793),
.Y(n_1395)
);

INVxp33_ASAP7_75t_SL g1396 ( 
.A(n_758),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_797),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_814),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1070),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_825),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_815),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_831),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_821),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_826),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_827),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_859),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_830),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1024),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_837),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_803),
.Y(n_1410)
);

INVxp33_ASAP7_75t_L g1411 ( 
.A(n_817),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_838),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_840),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_817),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_843),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_852),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1070),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_946),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_858),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_824),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_819),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_879),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_828),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_885),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_834),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_853),
.Y(n_1426)
);

INVxp67_ASAP7_75t_SL g1427 ( 
.A(n_824),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_887),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_888),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_898),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1359),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1327),
.Y(n_1432)
);

AND2x2_ASAP7_75t_SL g1433 ( 
.A(n_1325),
.B(n_913),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1361),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1402),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1330),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1315),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1365),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1294),
.A2(n_1059),
.B(n_948),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1331),
.Y(n_1440)
);

INVx5_ASAP7_75t_L g1441 ( 
.A(n_1408),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1342),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1330),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1360),
.Y(n_1444)
);

XNOR2x2_ASAP7_75t_L g1445 ( 
.A(n_1340),
.B(n_890),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1295),
.A2(n_1059),
.B(n_948),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1331),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1417),
.Y(n_1448)
);

INVx6_ASAP7_75t_L g1449 ( 
.A(n_1312),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1369),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_1300),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1417),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1373),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1293),
.B(n_851),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1339),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1387),
.B(n_1285),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1376),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1392),
.B(n_798),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1300),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1328),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1332),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1333),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1339),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1338),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1338),
.B(n_1024),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1293),
.B(n_955),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1326),
.A2(n_1231),
.B1(n_1266),
.B2(n_1205),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1410),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1343),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1334),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1335),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1336),
.Y(n_1472)
);

BUFx12f_ASAP7_75t_L g1473 ( 
.A(n_1302),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1343),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1378),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1299),
.B(n_1053),
.Y(n_1476)
);

INVx5_ASAP7_75t_L g1477 ( 
.A(n_1399),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1378),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_SL g1479 ( 
.A(n_1345),
.B(n_802),
.Y(n_1479)
);

CKINVDCx16_ASAP7_75t_R g1480 ( 
.A(n_1385),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1337),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1421),
.B(n_809),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1296),
.A2(n_1239),
.B(n_806),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1341),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1344),
.Y(n_1485)
);

BUFx6f_ASAP7_75t_L g1486 ( 
.A(n_1346),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1347),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1348),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1349),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1350),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1351),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1352),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1355),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1356),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1358),
.A2(n_1205),
.B1(n_1266),
.B2(n_1231),
.Y(n_1495)
);

BUFx8_ASAP7_75t_L g1496 ( 
.A(n_1304),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1299),
.B(n_1214),
.Y(n_1497)
);

CKINVDCx6p67_ASAP7_75t_R g1498 ( 
.A(n_1391),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1423),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1357),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1350),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1362),
.Y(n_1502)
);

INVx4_ASAP7_75t_L g1503 ( 
.A(n_1425),
.Y(n_1503)
);

INVx5_ASAP7_75t_L g1504 ( 
.A(n_1418),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1363),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1364),
.A2(n_1289),
.B1(n_1073),
.B2(n_876),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1389),
.B(n_1144),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1426),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1366),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1367),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1370),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1368),
.A2(n_1164),
.B1(n_1246),
.B2(n_1204),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1297),
.A2(n_1239),
.B(n_808),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1308),
.B(n_1309),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1371),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1305),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1311),
.B(n_1152),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1372),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1396),
.B(n_934),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1374),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1375),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1379),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1380),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1381),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1382),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1298),
.A2(n_1303),
.B(n_1301),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1383),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1313),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1384),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1388),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1307),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1386),
.Y(n_1532)
);

OAI22x1_ASAP7_75t_R g1533 ( 
.A1(n_1400),
.A2(n_1289),
.B1(n_1073),
.B2(n_886),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1388),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1390),
.A2(n_836),
.B(n_788),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1390),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1393),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1394),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1427),
.A2(n_850),
.B(n_849),
.Y(n_1539)
);

INVxp33_ASAP7_75t_SL g1540 ( 
.A(n_1310),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1314),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1329),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1306),
.A2(n_891),
.B1(n_901),
.B2(n_856),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1319),
.A2(n_1290),
.B1(n_1120),
.B2(n_1082),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1427),
.A2(n_871),
.B(n_854),
.Y(n_1545)
);

INVx3_ASAP7_75t_L g1546 ( 
.A(n_1316),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1377),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1395),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1317),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1377),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1318),
.B(n_1094),
.Y(n_1551)
);

INVx4_ASAP7_75t_L g1552 ( 
.A(n_1354),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1320),
.B(n_1152),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1397),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1414),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_L g1556 ( 
.A(n_1535),
.B(n_1401),
.C(n_1398),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1437),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1440),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1507),
.B(n_774),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1437),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1447),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1455),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1463),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1469),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1474),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1555),
.B(n_1389),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1475),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_SL g1568 ( 
.A(n_1512),
.B(n_908),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1437),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1435),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1442),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1478),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1555),
.B(n_1411),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1448),
.B(n_1411),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1442),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1541),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1549),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1526),
.B(n_946),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1537),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1537),
.Y(n_1580)
);

NAND2xp33_ASAP7_75t_SL g1581 ( 
.A(n_1544),
.B(n_967),
.Y(n_1581)
);

INVx4_ASAP7_75t_L g1582 ( 
.A(n_1443),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1442),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1449),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1444),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1490),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1444),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1526),
.B(n_946),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1436),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1479),
.A2(n_1014),
.B1(n_1022),
.B2(n_982),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1444),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1538),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1460),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1452),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1465),
.B(n_1321),
.Y(n_1595)
);

NAND2x1_ASAP7_75t_L g1596 ( 
.A(n_1439),
.B(n_771),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1538),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1527),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1527),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1460),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1460),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1439),
.B(n_946),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1530),
.B(n_1322),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1446),
.B(n_946),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1481),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1446),
.B(n_1539),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1527),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1532),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1457),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1535),
.B(n_946),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1481),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1433),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1532),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1481),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1497),
.B(n_1323),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1490),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1532),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1539),
.B(n_946),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1545),
.B(n_1158),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1501),
.B(n_1324),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1486),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1486),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1486),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_1488),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1548),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1449),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1451),
.B(n_774),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1548),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1548),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1488),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1554),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1554),
.Y(n_1632)
);

CKINVDCx11_ASAP7_75t_R g1633 ( 
.A(n_1432),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1488),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1492),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1554),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1529),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1492),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1545),
.B(n_875),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1514),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1514),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1501),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1484),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1551),
.A2(n_931),
.B(n_899),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1485),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1491),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1492),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1493),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1443),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1459),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1493),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1493),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1443),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1518),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1525),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1450),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1494),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1453),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1494),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1547),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1494),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1500),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1500),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1483),
.B(n_969),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1500),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1520),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1520),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1520),
.Y(n_1668)
);

OA21x2_ASAP7_75t_L g1669 ( 
.A1(n_1456),
.A2(n_996),
.B(n_985),
.Y(n_1669)
);

INVx1_ASAP7_75t_SL g1670 ( 
.A(n_1438),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1521),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1454),
.B(n_1414),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1521),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1483),
.B(n_1005),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_L g1675 ( 
.A(n_1534),
.B(n_1536),
.C(n_1513),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1521),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1523),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1523),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1513),
.B(n_1016),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1523),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1461),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1462),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1517),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1517),
.B(n_1403),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1528),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1454),
.B(n_1029),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1553),
.B(n_1404),
.Y(n_1687)
);

BUFx8_ASAP7_75t_L g1688 ( 
.A(n_1516),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1470),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1546),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1489),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1550),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1558),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1570),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1561),
.Y(n_1695)
);

AO21x2_ASAP7_75t_L g1696 ( 
.A1(n_1606),
.A2(n_1482),
.B(n_1458),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1566),
.B(n_1431),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1675),
.A2(n_1467),
.B1(n_1495),
.B2(n_1519),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1562),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1563),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1573),
.A2(n_1466),
.B1(n_1476),
.B2(n_1434),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1675),
.A2(n_1476),
.B1(n_1466),
.B2(n_1553),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1570),
.B(n_1431),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1584),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1574),
.B(n_1503),
.Y(n_1705)
);

CKINVDCx16_ASAP7_75t_R g1706 ( 
.A(n_1670),
.Y(n_1706)
);

AND2x6_ASAP7_75t_SL g1707 ( 
.A(n_1620),
.B(n_906),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1642),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1683),
.B(n_1503),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1586),
.B(n_1468),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1586),
.B(n_1672),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1616),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1683),
.B(n_1441),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1564),
.B(n_1499),
.Y(n_1714)
);

AO22x2_ASAP7_75t_L g1715 ( 
.A1(n_1559),
.A2(n_1533),
.B1(n_1054),
.B2(n_1055),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1683),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1681),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1615),
.B(n_1441),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1684),
.B(n_1441),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1594),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1686),
.A2(n_872),
.B1(n_897),
.B2(n_861),
.Y(n_1721)
);

INVx4_ASAP7_75t_L g1722 ( 
.A(n_1594),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1692),
.B(n_1508),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1565),
.B(n_1504),
.Y(n_1724)
);

BUFx10_ASAP7_75t_L g1725 ( 
.A(n_1684),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1567),
.B(n_1504),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1609),
.Y(n_1727)
);

AND3x2_ASAP7_75t_L g1728 ( 
.A(n_1612),
.B(n_1516),
.C(n_1531),
.Y(n_1728)
);

OR2x6_ASAP7_75t_L g1729 ( 
.A(n_1650),
.B(n_1473),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1572),
.Y(n_1730)
);

INVx4_ASAP7_75t_L g1731 ( 
.A(n_1601),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1692),
.Y(n_1732)
);

OAI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1686),
.A2(n_1406),
.B1(n_1353),
.B2(n_905),
.Y(n_1733)
);

BUFx10_ASAP7_75t_L g1734 ( 
.A(n_1687),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1639),
.A2(n_1036),
.B1(n_1063),
.B2(n_1039),
.Y(n_1735)
);

INVx4_ASAP7_75t_L g1736 ( 
.A(n_1601),
.Y(n_1736)
);

INVx6_ASAP7_75t_L g1737 ( 
.A(n_1688),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1687),
.B(n_1477),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1682),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1670),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1689),
.Y(n_1741)
);

INVxp33_ASAP7_75t_SL g1742 ( 
.A(n_1633),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1595),
.B(n_1464),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1643),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1645),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1660),
.B(n_1540),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1590),
.B(n_1480),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1594),
.B(n_1603),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1656),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1646),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1654),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1590),
.B(n_1498),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1619),
.B(n_1504),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1658),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1655),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1589),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1619),
.B(n_1471),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1576),
.B(n_1552),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1637),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1626),
.Y(n_1760)
);

INVx5_ASAP7_75t_L g1761 ( 
.A(n_1601),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1591),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1640),
.B(n_1641),
.Y(n_1763)
);

BUFx4f_ASAP7_75t_L g1764 ( 
.A(n_1669),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1603),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1577),
.B(n_1477),
.Y(n_1766)
);

INVx4_ASAP7_75t_L g1767 ( 
.A(n_1624),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1579),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1639),
.B(n_1472),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1580),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1592),
.B(n_1477),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1571),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1568),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1664),
.B(n_1674),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1685),
.B(n_1552),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1690),
.B(n_1598),
.Y(n_1776)
);

INVxp33_ASAP7_75t_L g1777 ( 
.A(n_1627),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1664),
.B(n_1487),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1591),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1691),
.Y(n_1780)
);

INVx5_ASAP7_75t_L g1781 ( 
.A(n_1624),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1597),
.B(n_1405),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1653),
.B(n_1420),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1591),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1557),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1556),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1581),
.Y(n_1787)
);

AND2x4_ASAP7_75t_L g1788 ( 
.A(n_1599),
.B(n_1407),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1607),
.B(n_1076),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1557),
.Y(n_1790)
);

INVx3_ASAP7_75t_L g1791 ( 
.A(n_1575),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1608),
.B(n_1613),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1674),
.B(n_1502),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1583),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1679),
.B(n_1505),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1556),
.A2(n_1135),
.B1(n_1180),
.B2(n_1118),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1560),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1624),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1560),
.Y(n_1799)
);

BUFx10_ASAP7_75t_L g1800 ( 
.A(n_1617),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1585),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1679),
.A2(n_1124),
.B1(n_1130),
.B2(n_1112),
.Y(n_1802)
);

INVxp33_ASAP7_75t_L g1803 ( 
.A(n_1669),
.Y(n_1803)
);

INVx3_ASAP7_75t_L g1804 ( 
.A(n_1587),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1625),
.Y(n_1805)
);

INVx5_ASAP7_75t_L g1806 ( 
.A(n_1630),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1688),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_1630),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1628),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1629),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1569),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1631),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1632),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1636),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1630),
.B(n_1233),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1606),
.B(n_1510),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1593),
.B(n_1409),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1649),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1638),
.B(n_1600),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1638),
.B(n_1250),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1578),
.B(n_1420),
.Y(n_1821)
);

AND2x6_ASAP7_75t_L g1822 ( 
.A(n_1610),
.B(n_771),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1569),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1623),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1659),
.B(n_1511),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1605),
.Y(n_1826)
);

INVx4_ASAP7_75t_L g1827 ( 
.A(n_1638),
.Y(n_1827)
);

INVx4_ASAP7_75t_L g1828 ( 
.A(n_1582),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1611),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1680),
.B(n_1542),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1614),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1662),
.B(n_1515),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1621),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1622),
.B(n_1412),
.Y(n_1834)
);

AND2x6_ASAP7_75t_L g1835 ( 
.A(n_1610),
.B(n_771),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_SL g1836 ( 
.A(n_1678),
.B(n_1256),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1663),
.A2(n_1274),
.B1(n_1123),
.B2(n_869),
.Y(n_1837)
);

AND3x2_ASAP7_75t_L g1838 ( 
.A(n_1634),
.B(n_1117),
.C(n_1035),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1635),
.B(n_1413),
.Y(n_1839)
);

INVx3_ASAP7_75t_L g1840 ( 
.A(n_1647),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1578),
.A2(n_1162),
.B1(n_1193),
.B2(n_1153),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1588),
.B(n_1445),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1651),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1588),
.A2(n_1216),
.B1(n_1243),
.B2(n_1202),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1652),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1618),
.A2(n_1263),
.B1(n_1272),
.B2(n_1244),
.Y(n_1846)
);

INVx2_ASAP7_75t_SL g1847 ( 
.A(n_1657),
.Y(n_1847)
);

INVx4_ASAP7_75t_L g1848 ( 
.A(n_1582),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1618),
.A2(n_1279),
.B1(n_1283),
.B2(n_1275),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1661),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1667),
.B(n_864),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1677),
.B(n_1543),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1623),
.Y(n_1853)
);

NAND2x1p5_ASAP7_75t_L g1854 ( 
.A(n_1716),
.B(n_1648),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1711),
.B(n_781),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1817),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1703),
.B(n_1668),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1817),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1834),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_L g1860 ( 
.A(n_1710),
.B(n_1506),
.Y(n_1860)
);

NOR2x1p5_ASAP7_75t_L g1861 ( 
.A(n_1752),
.B(n_759),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1701),
.B(n_1665),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1834),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1694),
.Y(n_1864)
);

INVxp67_ASAP7_75t_L g1865 ( 
.A(n_1712),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1842),
.B(n_1050),
.Y(n_1866)
);

NOR2xp67_ASAP7_75t_L g1867 ( 
.A(n_1746),
.B(n_1796),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1839),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1716),
.B(n_1666),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1774),
.B(n_1821),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1839),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1743),
.B(n_781),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1716),
.B(n_1671),
.Y(n_1873)
);

BUFx6f_ASAP7_75t_L g1874 ( 
.A(n_1784),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1702),
.B(n_1673),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1723),
.B(n_781),
.Y(n_1876)
);

NOR2xp67_ASAP7_75t_L g1877 ( 
.A(n_1722),
.B(n_1602),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1763),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1693),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1695),
.B(n_1648),
.Y(n_1880)
);

NAND3xp33_ASAP7_75t_L g1881 ( 
.A(n_1721),
.B(n_1496),
.C(n_1211),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1717),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1699),
.B(n_1676),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1700),
.B(n_1676),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1732),
.B(n_805),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1730),
.B(n_1602),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1786),
.B(n_1604),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1705),
.B(n_1604),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1696),
.B(n_1644),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1739),
.Y(n_1890)
);

NOR2xp67_ASAP7_75t_L g1891 ( 
.A(n_1756),
.B(n_1415),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1714),
.B(n_1045),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1802),
.B(n_1644),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1788),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1788),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1741),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1740),
.B(n_1046),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1735),
.B(n_1596),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1744),
.Y(n_1899)
);

INVx1_ASAP7_75t_SL g1900 ( 
.A(n_1708),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1742),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1698),
.B(n_1718),
.Y(n_1902)
);

NOR2x1p5_ASAP7_75t_L g1903 ( 
.A(n_1807),
.B(n_1747),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1841),
.B(n_1844),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1708),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1783),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1727),
.B(n_870),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1745),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1750),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1751),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_1697),
.B(n_1047),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1755),
.B(n_1292),
.Y(n_1912)
);

AND2x6_ASAP7_75t_SL g1913 ( 
.A(n_1729),
.B(n_912),
.Y(n_1913)
);

BUFx8_ASAP7_75t_L g1914 ( 
.A(n_1727),
.Y(n_1914)
);

INVxp33_ASAP7_75t_L g1915 ( 
.A(n_1852),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1782),
.Y(n_1916)
);

AND2x6_ASAP7_75t_L g1917 ( 
.A(n_1816),
.B(n_771),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1704),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1846),
.B(n_1524),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1782),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1787),
.B(n_884),
.Y(n_1921)
);

NOR2xp67_ASAP7_75t_L g1922 ( 
.A(n_1758),
.B(n_1837),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1849),
.B(n_1509),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1757),
.B(n_1522),
.Y(n_1924)
);

AOI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1773),
.A2(n_895),
.B1(n_900),
.B2(n_889),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1778),
.B(n_907),
.Y(n_1926)
);

INVxp67_ASAP7_75t_SL g1927 ( 
.A(n_1798),
.Y(n_1927)
);

OAI221xp5_ASAP7_75t_L g1928 ( 
.A1(n_1765),
.A2(n_1203),
.B1(n_1277),
.B2(n_1080),
.C(n_1077),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1733),
.B(n_914),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1793),
.B(n_922),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1749),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1795),
.B(n_923),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1769),
.B(n_947),
.Y(n_1933)
);

BUFx6f_ASAP7_75t_SL g1934 ( 
.A(n_1729),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1725),
.B(n_971),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1825),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1784),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1832),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1725),
.B(n_976),
.Y(n_1939)
);

INVx2_ASAP7_75t_SL g1940 ( 
.A(n_1706),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1822),
.B(n_1835),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1822),
.B(n_979),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1754),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_R g1944 ( 
.A(n_1720),
.B(n_1496),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1759),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1734),
.B(n_805),
.Y(n_1946)
);

A2O1A1Ixp33_ASAP7_75t_L g1947 ( 
.A1(n_1764),
.A2(n_1049),
.B(n_1092),
.C(n_794),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1803),
.A2(n_777),
.B1(n_892),
.B2(n_804),
.Y(n_1948)
);

NOR2x1p5_ASAP7_75t_L g1949 ( 
.A(n_1760),
.B(n_761),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1777),
.B(n_1048),
.Y(n_1950)
);

OAI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1780),
.A2(n_1100),
.B1(n_1101),
.B2(n_1084),
.Y(n_1951)
);

AOI22xp33_ASAP7_75t_L g1952 ( 
.A1(n_1822),
.A2(n_1835),
.B1(n_1715),
.B2(n_1809),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1805),
.Y(n_1953)
);

NAND2xp33_ASAP7_75t_L g1954 ( 
.A(n_1835),
.B(n_1798),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1734),
.B(n_980),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1810),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1794),
.B(n_990),
.Y(n_1957)
);

INVxp67_ASAP7_75t_L g1958 ( 
.A(n_1830),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1737),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1847),
.B(n_993),
.Y(n_1960)
);

NAND2xp33_ASAP7_75t_L g1961 ( 
.A(n_1798),
.B(n_994),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1808),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1812),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1813),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1762),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1814),
.B(n_998),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1779),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1808),
.B(n_1010),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1853),
.B(n_1021),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1824),
.B(n_1028),
.Y(n_1970)
);

NAND2xp33_ASAP7_75t_L g1971 ( 
.A(n_1808),
.B(n_1044),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1815),
.B(n_1145),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1820),
.B(n_1174),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1737),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1826),
.B(n_1051),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1761),
.B(n_1058),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1709),
.A2(n_1192),
.B1(n_1199),
.B2(n_1175),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1789),
.B(n_1206),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1836),
.B(n_805),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1761),
.B(n_1060),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1761),
.B(n_1074),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1748),
.B(n_810),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1831),
.B(n_1085),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1785),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1790),
.Y(n_1985)
);

AND2x4_ASAP7_75t_L g1986 ( 
.A(n_1768),
.B(n_1416),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1770),
.B(n_1235),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1833),
.A2(n_1850),
.B1(n_1843),
.B2(n_1776),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1801),
.Y(n_1989)
);

O2A1O1Ixp33_ASAP7_75t_L g1990 ( 
.A1(n_1851),
.A2(n_1247),
.B(n_1126),
.C(n_842),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1797),
.B(n_1799),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1811),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1823),
.B(n_1091),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1829),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1731),
.B(n_1099),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1772),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1781),
.B(n_1107),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1719),
.B(n_1713),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1775),
.B(n_1237),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1731),
.B(n_1114),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1736),
.B(n_1125),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1736),
.B(n_1131),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1784),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1800),
.B(n_1261),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1767),
.B(n_1136),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1767),
.B(n_1147),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1781),
.B(n_1148),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1818),
.B(n_1419),
.Y(n_2008)
);

INVx2_ASAP7_75t_SL g2009 ( 
.A(n_1838),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1781),
.B(n_1159),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1806),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1800),
.B(n_1255),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1840),
.B(n_1176),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1738),
.B(n_1422),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1845),
.B(n_1177),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1707),
.B(n_1287),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1806),
.B(n_1195),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1792),
.A2(n_1226),
.B1(n_1227),
.B2(n_1215),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1753),
.B(n_1228),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1724),
.A2(n_1259),
.B1(n_1280),
.B2(n_1251),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1791),
.B(n_777),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1728),
.B(n_1255),
.Y(n_2022)
);

AOI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_1715),
.A2(n_777),
.B1(n_892),
.B2(n_804),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1804),
.B(n_777),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1766),
.Y(n_2025)
);

OAI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1726),
.A2(n_929),
.B1(n_930),
.B2(n_924),
.C(n_919),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1905),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_1915),
.B(n_1828),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1867),
.B(n_1922),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1870),
.B(n_1848),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1899),
.Y(n_2031)
);

INVx4_ASAP7_75t_L g2032 ( 
.A(n_2011),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1909),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1879),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1908),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1910),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1936),
.B(n_1827),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1882),
.Y(n_2038)
);

NOR2x1_ASAP7_75t_L g2039 ( 
.A(n_1918),
.B(n_1819),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1866),
.B(n_1771),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1901),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1906),
.B(n_1806),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_1860),
.A2(n_774),
.B1(n_892),
.B2(n_804),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1958),
.B(n_1911),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1938),
.B(n_762),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1900),
.Y(n_2046)
);

INVx5_ASAP7_75t_L g2047 ( 
.A(n_2011),
.Y(n_2047)
);

AOI22x1_ASAP7_75t_L g2048 ( 
.A1(n_1931),
.A2(n_892),
.B1(n_902),
.B2(n_804),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1888),
.B(n_765),
.Y(n_2049)
);

BUFx2_ASAP7_75t_L g2050 ( 
.A(n_1914),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1864),
.B(n_1424),
.Y(n_2051)
);

INVxp67_ASAP7_75t_L g2052 ( 
.A(n_1940),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1887),
.B(n_766),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1953),
.Y(n_2054)
);

INVx4_ASAP7_75t_L g2055 ( 
.A(n_2011),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1956),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_2008),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1902),
.A2(n_1429),
.B1(n_1430),
.B2(n_1428),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1892),
.A2(n_779),
.B1(n_782),
.B2(n_769),
.Y(n_2059)
);

AOI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_1972),
.A2(n_784),
.B1(n_785),
.B2(n_783),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1963),
.Y(n_2061)
);

AND2x6_ASAP7_75t_SL g2062 ( 
.A(n_2016),
.B(n_933),
.Y(n_2062)
);

BUFx2_ASAP7_75t_L g2063 ( 
.A(n_1914),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1964),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_1959),
.Y(n_2065)
);

AND3x1_ASAP7_75t_L g2066 ( 
.A(n_1973),
.B(n_939),
.C(n_937),
.Y(n_2066)
);

NOR2x2_ASAP7_75t_L g2067 ( 
.A(n_1994),
.B(n_842),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1978),
.A2(n_1999),
.B1(n_1998),
.B2(n_1929),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1989),
.Y(n_2069)
);

NOR2x1p5_ASAP7_75t_L g2070 ( 
.A(n_1974),
.B(n_786),
.Y(n_2070)
);

NOR2xp67_ASAP7_75t_L g2071 ( 
.A(n_1865),
.B(n_550),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_1897),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1943),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1878),
.B(n_787),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_1986),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1890),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1886),
.B(n_790),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1926),
.B(n_795),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_1986),
.Y(n_2079)
);

BUFx12f_ASAP7_75t_L g2080 ( 
.A(n_1913),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1896),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1945),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1930),
.B(n_801),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_1874),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_1904),
.A2(n_902),
.B1(n_978),
.B2(n_911),
.Y(n_2085)
);

AND3x1_ASAP7_75t_L g2086 ( 
.A(n_1950),
.B(n_952),
.C(n_943),
.Y(n_2086)
);

BUFx6f_ASAP7_75t_L g2087 ( 
.A(n_1874),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1932),
.B(n_807),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_1855),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1933),
.B(n_811),
.Y(n_2090)
);

CKINVDCx20_ASAP7_75t_R g2091 ( 
.A(n_1944),
.Y(n_2091)
);

INVxp67_ASAP7_75t_L g2092 ( 
.A(n_1987),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1876),
.B(n_810),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_R g2094 ( 
.A(n_2004),
.B(n_813),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1924),
.B(n_816),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1880),
.Y(n_2096)
);

INVx5_ASAP7_75t_L g2097 ( 
.A(n_1874),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1883),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1872),
.B(n_818),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_SL g2100 ( 
.A(n_1934),
.B(n_1287),
.Y(n_2100)
);

OAI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1898),
.A2(n_829),
.B1(n_833),
.B2(n_823),
.Y(n_2101)
);

AND2x6_ASAP7_75t_L g2102 ( 
.A(n_1875),
.B(n_1278),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1884),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1984),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1934),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1858),
.Y(n_2106)
);

NAND2x1p5_ASAP7_75t_L g2107 ( 
.A(n_1937),
.B(n_902),
.Y(n_2107)
);

AND2x4_ASAP7_75t_L g2108 ( 
.A(n_1916),
.B(n_958),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1877),
.B(n_841),
.Y(n_2109)
);

AND2x4_ASAP7_75t_SL g2110 ( 
.A(n_1937),
.B(n_810),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_1937),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2023),
.B(n_844),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1985),
.Y(n_2113)
);

AND2x4_ASAP7_75t_L g2114 ( 
.A(n_1920),
.B(n_963),
.Y(n_2114)
);

O2A1O1Ixp33_ASAP7_75t_L g2115 ( 
.A1(n_1947),
.A2(n_972),
.B(n_974),
.C(n_964),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1992),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1912),
.B(n_845),
.Y(n_2117)
);

AND2x6_ASAP7_75t_L g2118 ( 
.A(n_1894),
.B(n_1895),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_2003),
.B(n_847),
.Y(n_2119)
);

BUFx4f_ASAP7_75t_L g2120 ( 
.A(n_2003),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_1977),
.B(n_848),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1979),
.B(n_855),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1982),
.B(n_860),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1859),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1856),
.B(n_863),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1863),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1951),
.B(n_866),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_1885),
.B(n_867),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_2003),
.B(n_868),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_1891),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1868),
.B(n_873),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1871),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1948),
.B(n_874),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1965),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1952),
.B(n_877),
.Y(n_2135)
);

BUFx12f_ASAP7_75t_L g2136 ( 
.A(n_1949),
.Y(n_2136)
);

OAI21xp5_ASAP7_75t_L g2137 ( 
.A1(n_1889),
.A2(n_992),
.B(n_989),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1967),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1946),
.B(n_1065),
.Y(n_2139)
);

AND2x4_ASAP7_75t_L g2140 ( 
.A(n_2025),
.B(n_1903),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2019),
.B(n_878),
.Y(n_2141)
);

INVx3_ASAP7_75t_L g2142 ( 
.A(n_1962),
.Y(n_2142)
);

NAND3xp33_ASAP7_75t_L g2143 ( 
.A(n_1925),
.B(n_881),
.C(n_880),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_2009),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1996),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1857),
.B(n_882),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1854),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1861),
.Y(n_2148)
);

AOI22xp5_ASAP7_75t_L g2149 ( 
.A1(n_1921),
.A2(n_883),
.B1(n_915),
.B2(n_904),
.Y(n_2149)
);

AND2x4_ASAP7_75t_L g2150 ( 
.A(n_2014),
.B(n_995),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1957),
.B(n_916),
.Y(n_2151)
);

INVxp67_ASAP7_75t_L g2152 ( 
.A(n_1907),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1960),
.B(n_917),
.Y(n_2153)
);

NOR3xp33_ASAP7_75t_SL g2154 ( 
.A(n_1881),
.B(n_920),
.C(n_918),
.Y(n_2154)
);

BUFx8_ASAP7_75t_L g2155 ( 
.A(n_2022),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1962),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1966),
.B(n_921),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_1935),
.Y(n_2158)
);

AOI22xp33_ASAP7_75t_L g2159 ( 
.A1(n_1862),
.A2(n_902),
.B1(n_978),
.B2(n_911),
.Y(n_2159)
);

OR2x6_ASAP7_75t_L g2160 ( 
.A(n_1939),
.B(n_857),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_1955),
.B(n_997),
.Y(n_2161)
);

NOR2xp67_ASAP7_75t_L g2162 ( 
.A(n_2012),
.B(n_551),
.Y(n_2162)
);

INVx5_ASAP7_75t_L g2163 ( 
.A(n_1917),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1991),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1988),
.Y(n_2165)
);

OAI22xp5_ASAP7_75t_SL g2166 ( 
.A1(n_1928),
.A2(n_949),
.B1(n_961),
.B2(n_932),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1927),
.B(n_926),
.Y(n_2167)
);

O2A1O1Ixp33_ASAP7_75t_L g2168 ( 
.A1(n_2026),
.A2(n_1011),
.B(n_1017),
.C(n_1006),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1995),
.B(n_927),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_1968),
.B(n_1026),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_L g2171 ( 
.A(n_1975),
.B(n_928),
.Y(n_2171)
);

AO22x1_ASAP7_75t_L g2172 ( 
.A1(n_1941),
.A2(n_936),
.B1(n_938),
.B2(n_935),
.Y(n_2172)
);

OR2x6_ASAP7_75t_L g2173 ( 
.A(n_1990),
.B(n_857),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_1869),
.B(n_1873),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1923),
.B(n_1065),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1919),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2021),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1969),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_1983),
.B(n_940),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2024),
.Y(n_2180)
);

NOR2xp67_ASAP7_75t_L g2181 ( 
.A(n_1942),
.B(n_553),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2046),
.Y(n_2182)
);

INVxp33_ASAP7_75t_L g2183 ( 
.A(n_2040),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_2065),
.Y(n_2184)
);

BUFx8_ASAP7_75t_L g2185 ( 
.A(n_2050),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2049),
.B(n_2053),
.Y(n_2186)
);

INVx3_ASAP7_75t_L g2187 ( 
.A(n_2047),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_2075),
.B(n_1976),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2034),
.Y(n_2189)
);

NOR2xp67_ASAP7_75t_L g2190 ( 
.A(n_2041),
.B(n_1970),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2068),
.B(n_2000),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2093),
.B(n_2020),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_2047),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2035),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2027),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2036),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2054),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2056),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2077),
.B(n_2001),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_2079),
.B(n_1980),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2061),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2030),
.B(n_2002),
.Y(n_2202)
);

BUFx3_ASAP7_75t_L g2203 ( 
.A(n_2140),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_SL g2204 ( 
.A(n_2072),
.B(n_2005),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_2171),
.B(n_2179),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_2087),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2164),
.B(n_2006),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2064),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2044),
.B(n_2013),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2069),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2092),
.B(n_1065),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2031),
.Y(n_2212)
);

NOR2xp67_ASAP7_75t_L g2213 ( 
.A(n_2089),
.B(n_1993),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2073),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_2057),
.B(n_2015),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2033),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2038),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2096),
.B(n_2018),
.Y(n_2218)
);

HB1xp67_ASAP7_75t_L g2219 ( 
.A(n_2052),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2098),
.B(n_2103),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2076),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2106),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2165),
.B(n_1981),
.Y(n_2223)
);

NAND2x1_ASAP7_75t_L g2224 ( 
.A(n_2118),
.B(n_1917),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2047),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2124),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2176),
.B(n_1997),
.Y(n_2227)
);

AND2x4_ASAP7_75t_L g2228 ( 
.A(n_2178),
.B(n_2007),
.Y(n_2228)
);

AND2x4_ASAP7_75t_L g2229 ( 
.A(n_2178),
.B(n_2010),
.Y(n_2229)
);

BUFx3_ASAP7_75t_L g2230 ( 
.A(n_2136),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_2039),
.B(n_2017),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2082),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2045),
.B(n_1961),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2078),
.B(n_1971),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2081),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2104),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2083),
.B(n_1917),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2139),
.B(n_2175),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_2028),
.B(n_1893),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2126),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2132),
.Y(n_2241)
);

NOR2xp33_ASAP7_75t_L g2242 ( 
.A(n_2029),
.B(n_944),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2113),
.Y(n_2243)
);

BUFx3_ASAP7_75t_L g2244 ( 
.A(n_2063),
.Y(n_2244)
);

AOI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2121),
.A2(n_1954),
.B1(n_1917),
.B2(n_950),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2116),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2134),
.Y(n_2247)
);

INVx4_ASAP7_75t_L g2248 ( 
.A(n_2097),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2088),
.B(n_1027),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_2090),
.B(n_945),
.Y(n_2250)
);

NOR2xp67_ASAP7_75t_L g2251 ( 
.A(n_2130),
.B(n_555),
.Y(n_2251)
);

CKINVDCx8_ASAP7_75t_R g2252 ( 
.A(n_2105),
.Y(n_2252)
);

INVx4_ASAP7_75t_L g2253 ( 
.A(n_2097),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2095),
.B(n_1032),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2150),
.B(n_1116),
.Y(n_2255)
);

BUFx2_ASAP7_75t_L g2256 ( 
.A(n_2097),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2152),
.A2(n_953),
.B1(n_956),
.B2(n_951),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2117),
.B(n_1034),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2138),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2145),
.Y(n_2260)
);

CKINVDCx11_ASAP7_75t_R g2261 ( 
.A(n_2080),
.Y(n_2261)
);

BUFx6f_ASAP7_75t_L g2262 ( 
.A(n_2087),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2037),
.B(n_2157),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2141),
.B(n_1038),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2169),
.B(n_1056),
.Y(n_2265)
);

BUFx6f_ASAP7_75t_L g2266 ( 
.A(n_2120),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_2122),
.B(n_957),
.Y(n_2267)
);

AOI22xp33_ASAP7_75t_SL g2268 ( 
.A1(n_2127),
.A2(n_1169),
.B1(n_1236),
.B2(n_1116),
.Y(n_2268)
);

AND2x6_ASAP7_75t_L g2269 ( 
.A(n_2177),
.B(n_911),
.Y(n_2269)
);

AND2x4_ASAP7_75t_L g2270 ( 
.A(n_2032),
.B(n_2055),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_L g2271 ( 
.A(n_2123),
.B(n_959),
.Y(n_2271)
);

INVx4_ASAP7_75t_L g2272 ( 
.A(n_2084),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2156),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2058),
.Y(n_2274)
);

OAI21x1_ASAP7_75t_L g2275 ( 
.A1(n_2180),
.A2(n_942),
.B(n_909),
.Y(n_2275)
);

AND3x1_ASAP7_75t_L g2276 ( 
.A(n_2154),
.B(n_1067),
.C(n_1062),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2151),
.B(n_1068),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2108),
.Y(n_2278)
);

NAND2xp33_ASAP7_75t_L g2279 ( 
.A(n_2118),
.B(n_911),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2114),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2094),
.B(n_2158),
.Y(n_2281)
);

NOR2xp33_ASAP7_75t_L g2282 ( 
.A(n_2153),
.B(n_962),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2142),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2099),
.B(n_2167),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2066),
.B(n_1116),
.Y(n_2285)
);

INVx4_ASAP7_75t_L g2286 ( 
.A(n_2111),
.Y(n_2286)
);

AOI21xp33_ASAP7_75t_L g2287 ( 
.A1(n_2112),
.A2(n_966),
.B(n_965),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_2158),
.B(n_1169),
.Y(n_2288)
);

AOI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2086),
.A2(n_970),
.B1(n_973),
.B2(n_968),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_2144),
.Y(n_2290)
);

BUFx3_ASAP7_75t_L g2291 ( 
.A(n_2091),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2147),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2125),
.Y(n_2293)
);

INVx4_ASAP7_75t_L g2294 ( 
.A(n_2118),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_2128),
.B(n_1169),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2135),
.B(n_1069),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2161),
.B(n_2060),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_2074),
.B(n_975),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_2174),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2107),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_R g2301 ( 
.A(n_2148),
.B(n_556),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2042),
.B(n_1072),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2131),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2146),
.Y(n_2304)
);

BUFx4f_ASAP7_75t_SL g2305 ( 
.A(n_2155),
.Y(n_2305)
);

BUFx8_ASAP7_75t_L g2306 ( 
.A(n_2170),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2173),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2173),
.Y(n_2308)
);

BUFx12f_ASAP7_75t_L g2309 ( 
.A(n_2070),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2109),
.Y(n_2310)
);

AND3x1_ASAP7_75t_SL g2311 ( 
.A(n_2067),
.B(n_1083),
.C(n_1081),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2051),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_2137),
.B(n_1088),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2101),
.B(n_1090),
.Y(n_2314)
);

AOI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2119),
.A2(n_981),
.B1(n_983),
.B2(n_977),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2059),
.B(n_2043),
.Y(n_2316)
);

NAND2xp33_ASAP7_75t_L g2317 ( 
.A(n_2102),
.B(n_978),
.Y(n_2317)
);

BUFx12f_ASAP7_75t_L g2318 ( 
.A(n_2062),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_2110),
.Y(n_2319)
);

INVx4_ASAP7_75t_L g2320 ( 
.A(n_2160),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2129),
.B(n_1095),
.Y(n_2321)
);

BUFx4f_ASAP7_75t_L g2322 ( 
.A(n_2160),
.Y(n_2322)
);

BUFx3_ASAP7_75t_L g2323 ( 
.A(n_2149),
.Y(n_2323)
);

BUFx2_ASAP7_75t_L g2324 ( 
.A(n_2102),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2071),
.B(n_2133),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2115),
.Y(n_2326)
);

BUFx12f_ASAP7_75t_L g2327 ( 
.A(n_2100),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2162),
.B(n_1236),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2102),
.B(n_1096),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2181),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_2143),
.Y(n_2331)
);

AND2x6_ASAP7_75t_L g2332 ( 
.A(n_2163),
.B(n_978),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_2166),
.B(n_1236),
.Y(n_2333)
);

INVx5_ASAP7_75t_L g2334 ( 
.A(n_2163),
.Y(n_2334)
);

OAI22xp5_ASAP7_75t_L g2335 ( 
.A1(n_2085),
.A2(n_987),
.B1(n_999),
.B2(n_984),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2172),
.B(n_2168),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2205),
.B(n_1000),
.Y(n_2337)
);

AOI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2191),
.A2(n_2163),
.B(n_2159),
.Y(n_2338)
);

O2A1O1Ixp5_ASAP7_75t_L g2339 ( 
.A1(n_2239),
.A2(n_1098),
.B(n_1104),
.C(n_1097),
.Y(n_2339)
);

AND2x2_ASAP7_75t_SL g2340 ( 
.A(n_2279),
.B(n_909),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2201),
.Y(n_2341)
);

OAI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_2323),
.A2(n_2186),
.B1(n_2263),
.B2(n_2316),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2210),
.Y(n_2343)
);

OAI21x1_ASAP7_75t_L g2344 ( 
.A1(n_2275),
.A2(n_2048),
.B(n_960),
.Y(n_2344)
);

OAI21x1_ASAP7_75t_L g2345 ( 
.A1(n_2224),
.A2(n_960),
.B(n_942),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2220),
.B(n_1001),
.Y(n_2346)
);

A2O1A1Ixp33_ASAP7_75t_L g2347 ( 
.A1(n_2250),
.A2(n_1008),
.B(n_1189),
.C(n_988),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_L g2348 ( 
.A1(n_2224),
.A2(n_1008),
.B(n_988),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2331),
.B(n_1264),
.Y(n_2349)
);

INVx3_ASAP7_75t_L g2350 ( 
.A(n_2266),
.Y(n_2350)
);

AOI21x1_ASAP7_75t_L g2351 ( 
.A1(n_2237),
.A2(n_1108),
.B(n_1106),
.Y(n_2351)
);

OAI21x1_ASAP7_75t_L g2352 ( 
.A1(n_2325),
.A2(n_1189),
.B(n_1110),
.Y(n_2352)
);

INVxp67_ASAP7_75t_SL g2353 ( 
.A(n_2195),
.Y(n_2353)
);

INVx2_ASAP7_75t_SL g2354 ( 
.A(n_2266),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2189),
.Y(n_2355)
);

OAI21x1_ASAP7_75t_L g2356 ( 
.A1(n_2202),
.A2(n_1119),
.B(n_1109),
.Y(n_2356)
);

AO31x2_ASAP7_75t_L g2357 ( 
.A1(n_2324),
.A2(n_1133),
.A3(n_1134),
.B(n_1127),
.Y(n_2357)
);

A2O1A1Ixp33_ASAP7_75t_L g2358 ( 
.A1(n_2282),
.A2(n_1139),
.B(n_1141),
.C(n_1138),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2293),
.B(n_1002),
.Y(n_2359)
);

OAI21x1_ASAP7_75t_L g2360 ( 
.A1(n_2330),
.A2(n_1146),
.B(n_1142),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2194),
.Y(n_2361)
);

INVx2_ASAP7_75t_SL g2362 ( 
.A(n_2290),
.Y(n_2362)
);

CKINVDCx5p33_ASAP7_75t_R g2363 ( 
.A(n_2305),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2284),
.B(n_1003),
.Y(n_2364)
);

OAI21x1_ASAP7_75t_SL g2365 ( 
.A1(n_2223),
.A2(n_1271),
.B(n_1270),
.Y(n_2365)
);

AOI21x1_ASAP7_75t_L g2366 ( 
.A1(n_2324),
.A2(n_1160),
.B(n_1151),
.Y(n_2366)
);

INVx5_ASAP7_75t_L g2367 ( 
.A(n_2248),
.Y(n_2367)
);

OAI21x1_ASAP7_75t_L g2368 ( 
.A1(n_2199),
.A2(n_1163),
.B(n_1161),
.Y(n_2368)
);

OAI22xp5_ASAP7_75t_L g2369 ( 
.A1(n_2268),
.A2(n_2322),
.B1(n_2183),
.B2(n_2233),
.Y(n_2369)
);

OAI21xp5_ASAP7_75t_L g2370 ( 
.A1(n_2267),
.A2(n_2271),
.B(n_2313),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2196),
.Y(n_2371)
);

NOR2xp67_ASAP7_75t_L g2372 ( 
.A(n_2310),
.B(n_557),
.Y(n_2372)
);

AOI21x1_ASAP7_75t_L g2373 ( 
.A1(n_2336),
.A2(n_1172),
.B(n_1166),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2303),
.B(n_1004),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_SL g2375 ( 
.A(n_2252),
.B(n_1264),
.Y(n_2375)
);

OAI21x1_ASAP7_75t_L g2376 ( 
.A1(n_2234),
.A2(n_1196),
.B(n_1187),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2212),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2304),
.B(n_1009),
.Y(n_2378)
);

BUFx3_ASAP7_75t_L g2379 ( 
.A(n_2184),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2207),
.A2(n_1031),
.B(n_1020),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2218),
.A2(n_1031),
.B(n_1020),
.Y(n_2381)
);

OAI21x1_ASAP7_75t_L g2382 ( 
.A1(n_2329),
.A2(n_1201),
.B(n_1198),
.Y(n_2382)
);

AO31x2_ASAP7_75t_L g2383 ( 
.A1(n_2326),
.A2(n_1208),
.A3(n_1209),
.B(n_1207),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2197),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2198),
.Y(n_2385)
);

BUFx3_ASAP7_75t_L g2386 ( 
.A(n_2290),
.Y(n_2386)
);

AOI21xp5_ASAP7_75t_L g2387 ( 
.A1(n_2317),
.A2(n_1031),
.B(n_1020),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2238),
.B(n_1012),
.Y(n_2388)
);

AOI21x1_ASAP7_75t_L g2389 ( 
.A1(n_2204),
.A2(n_1217),
.B(n_1213),
.Y(n_2389)
);

OAI21x1_ASAP7_75t_L g2390 ( 
.A1(n_2227),
.A2(n_1224),
.B(n_1219),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_2270),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_2331),
.B(n_2297),
.Y(n_2392)
);

BUFx8_ASAP7_75t_L g2393 ( 
.A(n_2327),
.Y(n_2393)
);

AOI21xp33_ASAP7_75t_L g2394 ( 
.A1(n_2314),
.A2(n_1234),
.B(n_1230),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2209),
.B(n_1013),
.Y(n_2395)
);

OAI21x1_ASAP7_75t_SL g2396 ( 
.A1(n_2294),
.A2(n_1291),
.B(n_1249),
.Y(n_2396)
);

OAI21x1_ASAP7_75t_L g2397 ( 
.A1(n_2232),
.A2(n_1252),
.B(n_1245),
.Y(n_2397)
);

OAI21x1_ASAP7_75t_L g2398 ( 
.A1(n_2235),
.A2(n_1276),
.B(n_1265),
.Y(n_2398)
);

AOI21xp33_ASAP7_75t_L g2399 ( 
.A1(n_2296),
.A2(n_1018),
.B(n_1015),
.Y(n_2399)
);

OAI21x1_ASAP7_75t_L g2400 ( 
.A1(n_2214),
.A2(n_1031),
.B(n_1020),
.Y(n_2400)
);

OAI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2299),
.A2(n_2192),
.B1(n_2312),
.B2(n_2242),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2249),
.B(n_1019),
.Y(n_2402)
);

OAI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2265),
.A2(n_1273),
.B(n_1269),
.Y(n_2403)
);

CKINVDCx20_ASAP7_75t_R g2404 ( 
.A(n_2261),
.Y(n_2404)
);

OAI21xp33_ASAP7_75t_L g2405 ( 
.A1(n_2298),
.A2(n_1025),
.B(n_1023),
.Y(n_2405)
);

OAI21xp5_ASAP7_75t_L g2406 ( 
.A1(n_2264),
.A2(n_1284),
.B(n_1282),
.Y(n_2406)
);

INVx3_ASAP7_75t_L g2407 ( 
.A(n_2270),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2277),
.B(n_1033),
.Y(n_2408)
);

OAI21x1_ASAP7_75t_L g2409 ( 
.A1(n_2208),
.A2(n_1278),
.B(n_563),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_2182),
.B(n_1037),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2258),
.B(n_1041),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_2231),
.B(n_1264),
.Y(n_2412)
);

OAI21x1_ASAP7_75t_L g2413 ( 
.A1(n_2222),
.A2(n_1278),
.B(n_569),
.Y(n_2413)
);

NAND3xp33_ASAP7_75t_L g2414 ( 
.A(n_2333),
.B(n_1043),
.C(n_1042),
.Y(n_2414)
);

OAI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_2254),
.A2(n_1258),
.B(n_1257),
.Y(n_2415)
);

OAI21x1_ASAP7_75t_L g2416 ( 
.A1(n_2226),
.A2(n_1278),
.B(n_570),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2211),
.B(n_1052),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2278),
.B(n_1057),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2240),
.Y(n_2419)
);

AOI21x1_ASAP7_75t_L g2420 ( 
.A1(n_2274),
.A2(n_571),
.B(n_561),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2280),
.B(n_1061),
.Y(n_2421)
);

A2O1A1Ixp33_ASAP7_75t_L g2422 ( 
.A1(n_2287),
.A2(n_1066),
.B(n_1075),
.C(n_1064),
.Y(n_2422)
);

AOI21xp5_ASAP7_75t_L g2423 ( 
.A1(n_2334),
.A2(n_2245),
.B(n_2215),
.Y(n_2423)
);

AND2x2_ASAP7_75t_SL g2424 ( 
.A(n_2276),
.B(n_0),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_L g2425 ( 
.A(n_2219),
.B(n_1078),
.Y(n_2425)
);

BUFx3_ASAP7_75t_L g2426 ( 
.A(n_2203),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_2272),
.Y(n_2427)
);

AOI221xp5_ASAP7_75t_L g2428 ( 
.A1(n_2285),
.A2(n_1087),
.B1(n_1089),
.B2(n_1086),
.C(n_1079),
.Y(n_2428)
);

BUFx6f_ASAP7_75t_SL g2429 ( 
.A(n_2230),
.Y(n_2429)
);

AOI22xp5_ASAP7_75t_L g2430 ( 
.A1(n_2295),
.A2(n_1102),
.B1(n_1103),
.B2(n_1093),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2228),
.B(n_2229),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2228),
.B(n_1105),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2241),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2229),
.B(n_1111),
.Y(n_2434)
);

INVx1_ASAP7_75t_SL g2435 ( 
.A(n_2291),
.Y(n_2435)
);

INVxp67_ASAP7_75t_L g2436 ( 
.A(n_2281),
.Y(n_2436)
);

AO21x2_ASAP7_75t_L g2437 ( 
.A1(n_2251),
.A2(n_574),
.B(n_572),
.Y(n_2437)
);

OAI22x1_ASAP7_75t_L g2438 ( 
.A1(n_2307),
.A2(n_1121),
.B1(n_1122),
.B2(n_1115),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2328),
.B(n_1128),
.Y(n_2439)
);

INVxp67_ASAP7_75t_SL g2440 ( 
.A(n_2292),
.Y(n_2440)
);

OAI21xp5_ASAP7_75t_SL g2441 ( 
.A1(n_2289),
.A2(n_1132),
.B(n_1129),
.Y(n_2441)
);

NAND3x1_ASAP7_75t_L g2442 ( 
.A(n_2319),
.B(n_1),
.C(n_3),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2334),
.A2(n_577),
.B(n_576),
.Y(n_2443)
);

OAI21x1_ASAP7_75t_L g2444 ( 
.A1(n_2308),
.A2(n_581),
.B(n_578),
.Y(n_2444)
);

NAND2xp33_ASAP7_75t_L g2445 ( 
.A(n_2334),
.B(n_1137),
.Y(n_2445)
);

OAI21x1_ASAP7_75t_L g2446 ( 
.A1(n_2273),
.A2(n_585),
.B(n_583),
.Y(n_2446)
);

BUFx3_ASAP7_75t_L g2447 ( 
.A(n_2206),
.Y(n_2447)
);

AND2x2_ASAP7_75t_SL g2448 ( 
.A(n_2320),
.B(n_4),
.Y(n_2448)
);

NAND2x1p5_ASAP7_75t_L g2449 ( 
.A(n_2253),
.B(n_586),
.Y(n_2449)
);

BUFx2_ASAP7_75t_L g2450 ( 
.A(n_2206),
.Y(n_2450)
);

OAI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_2213),
.A2(n_1288),
.B(n_1143),
.Y(n_2451)
);

INVx2_ASAP7_75t_SL g2452 ( 
.A(n_2262),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2217),
.B(n_1140),
.Y(n_2453)
);

CKINVDCx11_ASAP7_75t_R g2454 ( 
.A(n_2318),
.Y(n_2454)
);

AND2x6_ASAP7_75t_SL g2455 ( 
.A(n_2255),
.B(n_1149),
.Y(n_2455)
);

AO31x2_ASAP7_75t_L g2456 ( 
.A1(n_2243),
.A2(n_6),
.A3(n_4),
.B(n_5),
.Y(n_2456)
);

INVx1_ASAP7_75t_SL g2457 ( 
.A(n_2244),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2231),
.B(n_1238),
.Y(n_2458)
);

OAI21x1_ASAP7_75t_L g2459 ( 
.A1(n_2247),
.A2(n_588),
.B(n_587),
.Y(n_2459)
);

INVxp67_ASAP7_75t_SL g2460 ( 
.A(n_2216),
.Y(n_2460)
);

AOI21x1_ASAP7_75t_L g2461 ( 
.A1(n_2321),
.A2(n_591),
.B(n_589),
.Y(n_2461)
);

OAI21x1_ASAP7_75t_L g2462 ( 
.A1(n_2300),
.A2(n_598),
.B(n_596),
.Y(n_2462)
);

BUFx3_ASAP7_75t_L g2463 ( 
.A(n_2262),
.Y(n_2463)
);

AOI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_2256),
.A2(n_600),
.B(n_599),
.Y(n_2464)
);

AO31x2_ASAP7_75t_L g2465 ( 
.A1(n_2335),
.A2(n_9),
.A3(n_5),
.B(n_8),
.Y(n_2465)
);

OAI21x1_ASAP7_75t_L g2466 ( 
.A1(n_2221),
.A2(n_602),
.B(n_601),
.Y(n_2466)
);

AOI21x1_ASAP7_75t_L g2467 ( 
.A1(n_2190),
.A2(n_605),
.B(n_603),
.Y(n_2467)
);

BUFx6f_ASAP7_75t_L g2468 ( 
.A(n_2256),
.Y(n_2468)
);

OAI21x1_ASAP7_75t_L g2469 ( 
.A1(n_2236),
.A2(n_607),
.B(n_606),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2246),
.A2(n_610),
.B(n_608),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2302),
.B(n_1150),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2259),
.B(n_1154),
.Y(n_2472)
);

OAI21x1_ASAP7_75t_L g2473 ( 
.A1(n_2260),
.A2(n_613),
.B(n_612),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_2288),
.B(n_1156),
.Y(n_2474)
);

BUFx3_ASAP7_75t_L g2475 ( 
.A(n_2185),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2306),
.B(n_1167),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2306),
.B(n_1168),
.Y(n_2477)
);

OAI21xp5_ASAP7_75t_L g2478 ( 
.A1(n_2257),
.A2(n_1286),
.B(n_1171),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2302),
.B(n_1170),
.Y(n_2479)
);

OAI21x1_ASAP7_75t_L g2480 ( 
.A1(n_2283),
.A2(n_616),
.B(n_614),
.Y(n_2480)
);

AO31x2_ASAP7_75t_L g2481 ( 
.A1(n_2269),
.A2(n_2332),
.A3(n_2286),
.B(n_2311),
.Y(n_2481)
);

NAND2x1p5_ASAP7_75t_L g2482 ( 
.A(n_2187),
.B(n_2193),
.Y(n_2482)
);

A2O1A1Ixp33_ASAP7_75t_L g2483 ( 
.A1(n_2188),
.A2(n_1178),
.B(n_1179),
.C(n_1173),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2377),
.Y(n_2484)
);

INVx4_ASAP7_75t_L g2485 ( 
.A(n_2363),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2431),
.B(n_2188),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_SL g2487 ( 
.A(n_2370),
.B(n_2200),
.Y(n_2487)
);

INVx3_ASAP7_75t_L g2488 ( 
.A(n_2379),
.Y(n_2488)
);

BUFx3_ASAP7_75t_L g2489 ( 
.A(n_2447),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2355),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2342),
.B(n_2200),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2401),
.B(n_2315),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2361),
.Y(n_2493)
);

BUFx6f_ASAP7_75t_L g2494 ( 
.A(n_2463),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2371),
.Y(n_2495)
);

A2O1A1Ixp33_ASAP7_75t_SL g2496 ( 
.A1(n_2337),
.A2(n_2474),
.B(n_2381),
.C(n_2478),
.Y(n_2496)
);

HB1xp67_ASAP7_75t_L g2497 ( 
.A(n_2353),
.Y(n_2497)
);

OR2x6_ASAP7_75t_SL g2498 ( 
.A(n_2369),
.B(n_1181),
.Y(n_2498)
);

BUFx6f_ASAP7_75t_L g2499 ( 
.A(n_2386),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2341),
.Y(n_2500)
);

AOI21xp5_ASAP7_75t_L g2501 ( 
.A1(n_2340),
.A2(n_2269),
.B(n_2332),
.Y(n_2501)
);

OAI22xp5_ASAP7_75t_L g2502 ( 
.A1(n_2436),
.A2(n_2225),
.B1(n_2309),
.B2(n_1184),
.Y(n_2502)
);

OAI22xp5_ASAP7_75t_L g2503 ( 
.A1(n_2392),
.A2(n_1185),
.B1(n_1186),
.B2(n_1182),
.Y(n_2503)
);

AOI21xp33_ASAP7_75t_L g2504 ( 
.A1(n_2405),
.A2(n_2185),
.B(n_2269),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2468),
.B(n_2332),
.Y(n_2505)
);

BUFx12f_ASAP7_75t_L g2506 ( 
.A(n_2454),
.Y(n_2506)
);

CKINVDCx5p33_ASAP7_75t_R g2507 ( 
.A(n_2404),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2468),
.B(n_618),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2384),
.Y(n_2509)
);

BUFx3_ASAP7_75t_L g2510 ( 
.A(n_2450),
.Y(n_2510)
);

CKINVDCx5p33_ASAP7_75t_R g2511 ( 
.A(n_2393),
.Y(n_2511)
);

NOR2x1_ASAP7_75t_SL g2512 ( 
.A(n_2437),
.B(n_2373),
.Y(n_2512)
);

OAI22xp33_ASAP7_75t_L g2513 ( 
.A1(n_2375),
.A2(n_1268),
.B1(n_1281),
.B2(n_1267),
.Y(n_2513)
);

OR2x6_ASAP7_75t_L g2514 ( 
.A(n_2449),
.B(n_2301),
.Y(n_2514)
);

AOI21xp5_ASAP7_75t_L g2515 ( 
.A1(n_2338),
.A2(n_1190),
.B(n_1188),
.Y(n_2515)
);

NOR2xp33_ASAP7_75t_L g2516 ( 
.A(n_2435),
.B(n_1194),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2385),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2440),
.B(n_2343),
.Y(n_2518)
);

A2O1A1Ixp33_ASAP7_75t_SL g2519 ( 
.A1(n_2394),
.A2(n_1200),
.B(n_1210),
.C(n_1197),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2468),
.B(n_619),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2460),
.B(n_1225),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2419),
.Y(n_2522)
);

OR2x2_ASAP7_75t_L g2523 ( 
.A(n_2433),
.B(n_8),
.Y(n_2523)
);

BUFx2_ASAP7_75t_L g2524 ( 
.A(n_2352),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2424),
.B(n_620),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2364),
.B(n_1241),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_2482),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2383),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_L g2529 ( 
.A(n_2458),
.B(n_1212),
.Y(n_2529)
);

AOI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_2414),
.A2(n_1220),
.B1(n_1222),
.B2(n_1218),
.Y(n_2530)
);

BUFx2_ASAP7_75t_L g2531 ( 
.A(n_2383),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2395),
.B(n_1262),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2357),
.B(n_622),
.Y(n_2533)
);

INVx1_ASAP7_75t_SL g2534 ( 
.A(n_2457),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2346),
.B(n_1223),
.Y(n_2535)
);

AND2x4_ASAP7_75t_L g2536 ( 
.A(n_2391),
.B(n_625),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_L g2537 ( 
.A(n_2349),
.B(n_1229),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2383),
.Y(n_2538)
);

O2A1O1Ixp5_ASAP7_75t_SL g2539 ( 
.A1(n_2412),
.A2(n_1242),
.B(n_1253),
.C(n_1232),
.Y(n_2539)
);

INVx3_ASAP7_75t_L g2540 ( 
.A(n_2426),
.Y(n_2540)
);

A2O1A1Ixp33_ASAP7_75t_L g2541 ( 
.A1(n_2399),
.A2(n_1260),
.B(n_1254),
.C(n_13),
.Y(n_2541)
);

NAND2x1p5_ASAP7_75t_L g2542 ( 
.A(n_2367),
.B(n_626),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2456),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2350),
.Y(n_2544)
);

HB1xp67_ASAP7_75t_L g2545 ( 
.A(n_2407),
.Y(n_2545)
);

O2A1O1Ixp5_ASAP7_75t_SL g2546 ( 
.A1(n_2451),
.A2(n_2403),
.B(n_2415),
.C(n_2406),
.Y(n_2546)
);

BUFx3_ASAP7_75t_L g2547 ( 
.A(n_2354),
.Y(n_2547)
);

INVxp67_ASAP7_75t_SL g2548 ( 
.A(n_2423),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2397),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2372),
.B(n_10),
.Y(n_2550)
);

OAI22xp5_ASAP7_75t_L g2551 ( 
.A1(n_2483),
.A2(n_2432),
.B1(n_2434),
.B2(n_2430),
.Y(n_2551)
);

INVx1_ASAP7_75t_SL g2552 ( 
.A(n_2410),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2359),
.B(n_10),
.Y(n_2553)
);

BUFx3_ASAP7_75t_L g2554 ( 
.A(n_2362),
.Y(n_2554)
);

HB1xp67_ASAP7_75t_L g2555 ( 
.A(n_2356),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2456),
.Y(n_2556)
);

INVx4_ASAP7_75t_L g2557 ( 
.A(n_2367),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2441),
.A2(n_2471),
.B1(n_2448),
.B2(n_2445),
.Y(n_2558)
);

INVx3_ASAP7_75t_SL g2559 ( 
.A(n_2475),
.Y(n_2559)
);

NAND2x1_ASAP7_75t_L g2560 ( 
.A(n_2365),
.B(n_627),
.Y(n_2560)
);

OAI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2439),
.A2(n_2442),
.B1(n_2479),
.B2(n_2422),
.Y(n_2561)
);

OR2x2_ASAP7_75t_L g2562 ( 
.A(n_2357),
.B(n_11),
.Y(n_2562)
);

AOI21xp5_ASAP7_75t_L g2563 ( 
.A1(n_2380),
.A2(n_2387),
.B(n_2470),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2398),
.Y(n_2564)
);

AOI21xp5_ASAP7_75t_L g2565 ( 
.A1(n_2443),
.A2(n_630),
.B(n_629),
.Y(n_2565)
);

OR2x6_ASAP7_75t_L g2566 ( 
.A(n_2464),
.B(n_633),
.Y(n_2566)
);

INVx3_ASAP7_75t_L g2567 ( 
.A(n_2427),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2456),
.Y(n_2568)
);

AOI21xp5_ASAP7_75t_L g2569 ( 
.A1(n_2344),
.A2(n_637),
.B(n_635),
.Y(n_2569)
);

AOI22xp33_ASAP7_75t_L g2570 ( 
.A1(n_2438),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_2393),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2357),
.B(n_638),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2347),
.B(n_639),
.Y(n_2573)
);

CKINVDCx8_ASAP7_75t_R g2574 ( 
.A(n_2455),
.Y(n_2574)
);

AOI21xp5_ASAP7_75t_L g2575 ( 
.A1(n_2400),
.A2(n_2368),
.B(n_2376),
.Y(n_2575)
);

OR2x6_ASAP7_75t_L g2576 ( 
.A(n_2396),
.B(n_646),
.Y(n_2576)
);

AOI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_2345),
.A2(n_648),
.B(n_647),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2452),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2389),
.Y(n_2579)
);

INVx2_ASAP7_75t_SL g2580 ( 
.A(n_2367),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2428),
.A2(n_18),
.B1(n_14),
.B2(n_17),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2465),
.B(n_649),
.Y(n_2582)
);

BUFx3_ASAP7_75t_L g2583 ( 
.A(n_2476),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2465),
.Y(n_2584)
);

INVx2_ASAP7_75t_SL g2585 ( 
.A(n_2477),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2374),
.B(n_18),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_SL g2587 ( 
.A(n_2366),
.B(n_2402),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2408),
.B(n_650),
.Y(n_2588)
);

AND2x4_ASAP7_75t_L g2589 ( 
.A(n_2497),
.B(n_2444),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2518),
.B(n_2465),
.Y(n_2590)
);

HB1xp67_ASAP7_75t_L g2591 ( 
.A(n_2522),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2500),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2486),
.B(n_2481),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2490),
.Y(n_2594)
);

OR2x6_ASAP7_75t_SL g2595 ( 
.A(n_2511),
.B(n_2388),
.Y(n_2595)
);

O2A1O1Ixp33_ASAP7_75t_SL g2596 ( 
.A1(n_2496),
.A2(n_2358),
.B(n_2378),
.C(n_2417),
.Y(n_2596)
);

NAND2xp33_ASAP7_75t_L g2597 ( 
.A(n_2541),
.B(n_2411),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2493),
.B(n_2481),
.Y(n_2598)
);

NOR2xp33_ASAP7_75t_L g2599 ( 
.A(n_2534),
.B(n_2425),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2491),
.B(n_2453),
.Y(n_2600)
);

AND2x4_ASAP7_75t_L g2601 ( 
.A(n_2495),
.B(n_2462),
.Y(n_2601)
);

AND2x4_ASAP7_75t_L g2602 ( 
.A(n_2509),
.B(n_2480),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2548),
.B(n_2472),
.Y(n_2603)
);

INVx2_ASAP7_75t_SL g2604 ( 
.A(n_2489),
.Y(n_2604)
);

O2A1O1Ixp5_ASAP7_75t_L g2605 ( 
.A1(n_2565),
.A2(n_2420),
.B(n_2351),
.C(n_2467),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2517),
.B(n_2418),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2487),
.B(n_2481),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2528),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2538),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2484),
.Y(n_2610)
);

AOI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2563),
.A2(n_2390),
.B(n_2339),
.Y(n_2611)
);

OR2x2_ASAP7_75t_L g2612 ( 
.A(n_2531),
.B(n_2421),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2531),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2545),
.B(n_2409),
.Y(n_2614)
);

INVx3_ASAP7_75t_L g2615 ( 
.A(n_2557),
.Y(n_2615)
);

BUFx2_ASAP7_75t_L g2616 ( 
.A(n_2510),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2582),
.B(n_2413),
.Y(n_2617)
);

OAI22xp5_ASAP7_75t_L g2618 ( 
.A1(n_2498),
.A2(n_2429),
.B1(n_2461),
.B2(n_2360),
.Y(n_2618)
);

HB1xp67_ASAP7_75t_L g2619 ( 
.A(n_2584),
.Y(n_2619)
);

O2A1O1Ixp33_ASAP7_75t_L g2620 ( 
.A1(n_2561),
.A2(n_2382),
.B(n_2416),
.C(n_2459),
.Y(n_2620)
);

AOI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_2566),
.A2(n_2348),
.B(n_2446),
.Y(n_2621)
);

A2O1A1Ixp33_ASAP7_75t_L g2622 ( 
.A1(n_2558),
.A2(n_2537),
.B(n_2529),
.C(n_2588),
.Y(n_2622)
);

INVx2_ASAP7_75t_SL g2623 ( 
.A(n_2494),
.Y(n_2623)
);

BUFx3_ASAP7_75t_L g2624 ( 
.A(n_2494),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2525),
.B(n_2466),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2527),
.B(n_2469),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2552),
.B(n_19),
.Y(n_2627)
);

O2A1O1Ixp33_ASAP7_75t_L g2628 ( 
.A1(n_2587),
.A2(n_22),
.B(n_20),
.C(n_21),
.Y(n_2628)
);

INVxp67_ASAP7_75t_L g2629 ( 
.A(n_2578),
.Y(n_2629)
);

INVxp67_ASAP7_75t_L g2630 ( 
.A(n_2554),
.Y(n_2630)
);

BUFx5_ASAP7_75t_L g2631 ( 
.A(n_2543),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2533),
.B(n_2473),
.Y(n_2632)
);

NOR2xp67_ASAP7_75t_L g2633 ( 
.A(n_2567),
.B(n_21),
.Y(n_2633)
);

A2O1A1Ixp33_ASAP7_75t_L g2634 ( 
.A1(n_2504),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2556),
.Y(n_2635)
);

CKINVDCx11_ASAP7_75t_R g2636 ( 
.A(n_2506),
.Y(n_2636)
);

BUFx3_ASAP7_75t_L g2637 ( 
.A(n_2499),
.Y(n_2637)
);

A2O1A1Ixp33_ASAP7_75t_L g2638 ( 
.A1(n_2581),
.A2(n_26),
.B(n_23),
.C(n_25),
.Y(n_2638)
);

INVx2_ASAP7_75t_SL g2639 ( 
.A(n_2499),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2568),
.B(n_26),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2555),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2572),
.B(n_27),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2549),
.Y(n_2643)
);

CKINVDCx6p67_ASAP7_75t_R g2644 ( 
.A(n_2559),
.Y(n_2644)
);

A2O1A1Ixp33_ASAP7_75t_SL g2645 ( 
.A1(n_2515),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_2645)
);

OA21x2_ASAP7_75t_L g2646 ( 
.A1(n_2575),
.A2(n_29),
.B(n_30),
.Y(n_2646)
);

A2O1A1Ixp33_ASAP7_75t_L g2647 ( 
.A1(n_2492),
.A2(n_34),
.B(n_31),
.C(n_32),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2523),
.B(n_31),
.Y(n_2648)
);

OR2x6_ASAP7_75t_SL g2649 ( 
.A(n_2571),
.B(n_34),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2580),
.B(n_755),
.Y(n_2650)
);

HB1xp67_ASAP7_75t_L g2651 ( 
.A(n_2524),
.Y(n_2651)
);

O2A1O1Ixp5_ASAP7_75t_L g2652 ( 
.A1(n_2501),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2564),
.Y(n_2653)
);

NAND2x1p5_ASAP7_75t_L g2654 ( 
.A(n_2505),
.B(n_659),
.Y(n_2654)
);

A2O1A1Ixp33_ASAP7_75t_L g2655 ( 
.A1(n_2551),
.A2(n_2570),
.B(n_2553),
.C(n_2586),
.Y(n_2655)
);

HB1xp67_ASAP7_75t_L g2656 ( 
.A(n_2524),
.Y(n_2656)
);

O2A1O1Ixp5_ASAP7_75t_L g2657 ( 
.A1(n_2560),
.A2(n_40),
.B(n_36),
.C(n_39),
.Y(n_2657)
);

BUFx2_ASAP7_75t_L g2658 ( 
.A(n_2540),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2585),
.B(n_39),
.Y(n_2659)
);

INVxp33_ASAP7_75t_SL g2660 ( 
.A(n_2507),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2579),
.Y(n_2661)
);

A2O1A1Ixp33_ASAP7_75t_SL g2662 ( 
.A1(n_2516),
.A2(n_45),
.B(n_41),
.C(n_42),
.Y(n_2662)
);

AOI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_2566),
.A2(n_663),
.B(n_660),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2562),
.Y(n_2664)
);

AND2x4_ASAP7_75t_L g2665 ( 
.A(n_2505),
.B(n_745),
.Y(n_2665)
);

OA21x2_ASAP7_75t_L g2666 ( 
.A1(n_2569),
.A2(n_2577),
.B(n_2550),
.Y(n_2666)
);

BUFx6f_ASAP7_75t_L g2667 ( 
.A(n_2544),
.Y(n_2667)
);

OAI21xp5_ASAP7_75t_L g2668 ( 
.A1(n_2622),
.A2(n_2546),
.B(n_2573),
.Y(n_2668)
);

BUFx3_ASAP7_75t_L g2669 ( 
.A(n_2644),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2594),
.Y(n_2670)
);

HB1xp67_ASAP7_75t_L g2671 ( 
.A(n_2619),
.Y(n_2671)
);

HB1xp67_ASAP7_75t_L g2672 ( 
.A(n_2651),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2591),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2593),
.B(n_2616),
.Y(n_2674)
);

OA21x2_ASAP7_75t_L g2675 ( 
.A1(n_2608),
.A2(n_2521),
.B(n_2532),
.Y(n_2675)
);

OAI21x1_ASAP7_75t_L g2676 ( 
.A1(n_2611),
.A2(n_2542),
.B(n_2539),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2592),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2610),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2615),
.Y(n_2679)
);

BUFx6f_ASAP7_75t_L g2680 ( 
.A(n_2667),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2609),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2661),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2661),
.Y(n_2683)
);

OR2x6_ASAP7_75t_L g2684 ( 
.A(n_2621),
.B(n_2589),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2658),
.B(n_2583),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2635),
.Y(n_2686)
);

AND2x4_ASAP7_75t_L g2687 ( 
.A(n_2589),
.B(n_2488),
.Y(n_2687)
);

INVx3_ASAP7_75t_L g2688 ( 
.A(n_2615),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2664),
.Y(n_2689)
);

HB1xp67_ASAP7_75t_L g2690 ( 
.A(n_2656),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2641),
.Y(n_2691)
);

OR2x6_ASAP7_75t_L g2692 ( 
.A(n_2607),
.B(n_2514),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2590),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2598),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2613),
.Y(n_2695)
);

AND2x4_ASAP7_75t_L g2696 ( 
.A(n_2601),
.B(n_2547),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2643),
.Y(n_2697)
);

INVx2_ASAP7_75t_SL g2698 ( 
.A(n_2604),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2653),
.Y(n_2699)
);

AND2x4_ASAP7_75t_L g2700 ( 
.A(n_2601),
.B(n_2508),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2612),
.Y(n_2701)
);

INVx3_ASAP7_75t_L g2702 ( 
.A(n_2602),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2631),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2631),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2631),
.Y(n_2705)
);

INVx2_ASAP7_75t_SL g2706 ( 
.A(n_2624),
.Y(n_2706)
);

OAI21x1_ASAP7_75t_L g2707 ( 
.A1(n_2605),
.A2(n_2512),
.B(n_2502),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2631),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2606),
.B(n_2526),
.Y(n_2709)
);

AND2x4_ASAP7_75t_L g2710 ( 
.A(n_2602),
.B(n_2614),
.Y(n_2710)
);

OAI21x1_ASAP7_75t_L g2711 ( 
.A1(n_2620),
.A2(n_2503),
.B(n_2535),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2626),
.Y(n_2712)
);

NAND2x1p5_ASAP7_75t_L g2713 ( 
.A(n_2666),
.B(n_2508),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2640),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2630),
.B(n_2544),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2646),
.Y(n_2716)
);

NOR2xp67_ASAP7_75t_R g2717 ( 
.A(n_2637),
.B(n_2485),
.Y(n_2717)
);

OA21x2_ASAP7_75t_L g2718 ( 
.A1(n_2652),
.A2(n_2657),
.B(n_2603),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2646),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2667),
.Y(n_2720)
);

BUFx2_ASAP7_75t_L g2721 ( 
.A(n_2625),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2617),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2595),
.B(n_2629),
.Y(n_2723)
);

HB1xp67_ASAP7_75t_L g2724 ( 
.A(n_2600),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2667),
.Y(n_2725)
);

OAI21xp5_ASAP7_75t_L g2726 ( 
.A1(n_2655),
.A2(n_2576),
.B(n_2513),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2632),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_SL g2728 ( 
.A(n_2618),
.B(n_2520),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2666),
.B(n_2520),
.Y(n_2729)
);

BUFx3_ASAP7_75t_L g2730 ( 
.A(n_2636),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2659),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2627),
.Y(n_2732)
);

AO31x2_ASAP7_75t_L g2733 ( 
.A1(n_2647),
.A2(n_2576),
.A3(n_2519),
.B(n_2514),
.Y(n_2733)
);

AND2x4_ASAP7_75t_L g2734 ( 
.A(n_2623),
.B(n_2536),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2639),
.Y(n_2735)
);

BUFx2_ASAP7_75t_L g2736 ( 
.A(n_2650),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2648),
.Y(n_2737)
);

OA21x2_ASAP7_75t_L g2738 ( 
.A1(n_2634),
.A2(n_2530),
.B(n_2536),
.Y(n_2738)
);

NOR2xp33_ASAP7_75t_L g2739 ( 
.A(n_2596),
.B(n_2574),
.Y(n_2739)
);

OAI21x1_ASAP7_75t_L g2740 ( 
.A1(n_2663),
.A2(n_2628),
.B(n_2654),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2710),
.B(n_2665),
.Y(n_2741)
);

HB1xp67_ASAP7_75t_L g2742 ( 
.A(n_2671),
.Y(n_2742)
);

OR2x2_ASAP7_75t_L g2743 ( 
.A(n_2701),
.B(n_2642),
.Y(n_2743)
);

INVxp67_ASAP7_75t_L g2744 ( 
.A(n_2675),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2689),
.Y(n_2745)
);

INVx3_ASAP7_75t_L g2746 ( 
.A(n_2687),
.Y(n_2746)
);

INVx4_ASAP7_75t_L g2747 ( 
.A(n_2730),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2674),
.B(n_2721),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2724),
.B(n_2599),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2724),
.B(n_2649),
.Y(n_2750)
);

BUFx3_ASAP7_75t_L g2751 ( 
.A(n_2730),
.Y(n_2751)
);

HB1xp67_ASAP7_75t_L g2752 ( 
.A(n_2672),
.Y(n_2752)
);

OR2x2_ASAP7_75t_L g2753 ( 
.A(n_2693),
.B(n_2633),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2710),
.B(n_2650),
.Y(n_2754)
);

INVxp33_ASAP7_75t_L g2755 ( 
.A(n_2685),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2671),
.Y(n_2756)
);

AOI22xp33_ASAP7_75t_L g2757 ( 
.A1(n_2668),
.A2(n_2597),
.B1(n_2665),
.B2(n_2660),
.Y(n_2757)
);

INVx1_ASAP7_75t_SL g2758 ( 
.A(n_2672),
.Y(n_2758)
);

INVx3_ASAP7_75t_L g2759 ( 
.A(n_2687),
.Y(n_2759)
);

NAND2x1_ASAP7_75t_L g2760 ( 
.A(n_2684),
.B(n_2662),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2670),
.Y(n_2761)
);

INVxp67_ASAP7_75t_L g2762 ( 
.A(n_2675),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2681),
.Y(n_2763)
);

INVx4_ASAP7_75t_L g2764 ( 
.A(n_2669),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2691),
.B(n_2645),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2673),
.B(n_2638),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2690),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2690),
.Y(n_2768)
);

OR2x2_ASAP7_75t_L g2769 ( 
.A(n_2722),
.B(n_41),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2677),
.B(n_42),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2682),
.Y(n_2771)
);

HB1xp67_ASAP7_75t_L g2772 ( 
.A(n_2682),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2683),
.Y(n_2773)
);

AND2x4_ASAP7_75t_SL g2774 ( 
.A(n_2734),
.B(n_748),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2712),
.Y(n_2775)
);

NOR2x1_ASAP7_75t_L g2776 ( 
.A(n_2669),
.B(n_45),
.Y(n_2776)
);

INVx4_ASAP7_75t_L g2777 ( 
.A(n_2680),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2683),
.Y(n_2778)
);

NOR2xp67_ASAP7_75t_L g2779 ( 
.A(n_2702),
.B(n_46),
.Y(n_2779)
);

INVx3_ASAP7_75t_L g2780 ( 
.A(n_2696),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2686),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2678),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2742),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2772),
.Y(n_2784)
);

INVx3_ASAP7_75t_L g2785 ( 
.A(n_2746),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2746),
.B(n_2702),
.Y(n_2786)
);

BUFx2_ASAP7_75t_L g2787 ( 
.A(n_2764),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2772),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2749),
.B(n_2714),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2759),
.B(n_2723),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2759),
.B(n_2684),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2780),
.B(n_2684),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2742),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2753),
.B(n_2732),
.Y(n_2794)
);

OR2x2_ASAP7_75t_L g2795 ( 
.A(n_2743),
.B(n_2758),
.Y(n_2795)
);

HB1xp67_ASAP7_75t_L g2796 ( 
.A(n_2752),
.Y(n_2796)
);

INVx3_ASAP7_75t_L g2797 ( 
.A(n_2780),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2756),
.Y(n_2798)
);

OR2x2_ASAP7_75t_L g2799 ( 
.A(n_2758),
.B(n_2727),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2748),
.B(n_2692),
.Y(n_2800)
);

INVxp67_ASAP7_75t_SL g2801 ( 
.A(n_2744),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2763),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2761),
.Y(n_2803)
);

INVx4_ASAP7_75t_L g2804 ( 
.A(n_2747),
.Y(n_2804)
);

INVx2_ASAP7_75t_SL g2805 ( 
.A(n_2764),
.Y(n_2805)
);

INVx5_ASAP7_75t_L g2806 ( 
.A(n_2747),
.Y(n_2806)
);

BUFx2_ASAP7_75t_L g2807 ( 
.A(n_2777),
.Y(n_2807)
);

NAND2x1_ASAP7_75t_L g2808 ( 
.A(n_2767),
.B(n_2692),
.Y(n_2808)
);

INVxp67_ASAP7_75t_SL g2809 ( 
.A(n_2744),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2771),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2755),
.B(n_2692),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2768),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2781),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2773),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2778),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2762),
.Y(n_2816)
);

AND2x2_ASAP7_75t_L g2817 ( 
.A(n_2750),
.B(n_2696),
.Y(n_2817)
);

INVx2_ASAP7_75t_SL g2818 ( 
.A(n_2751),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2762),
.B(n_2694),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2813),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2802),
.Y(n_2821)
);

AOI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2790),
.A2(n_2739),
.B1(n_2668),
.B2(n_2726),
.Y(n_2822)
);

OR2x2_ASAP7_75t_L g2823 ( 
.A(n_2795),
.B(n_2765),
.Y(n_2823)
);

AND2x2_ASAP7_75t_L g2824 ( 
.A(n_2790),
.B(n_2754),
.Y(n_2824)
);

AND2x4_ASAP7_75t_L g2825 ( 
.A(n_2806),
.B(n_2741),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2798),
.Y(n_2826)
);

HB1xp67_ASAP7_75t_L g2827 ( 
.A(n_2796),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2797),
.Y(n_2828)
);

AND2x4_ASAP7_75t_SL g2829 ( 
.A(n_2804),
.B(n_2741),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2812),
.Y(n_2830)
);

HB1xp67_ASAP7_75t_L g2831 ( 
.A(n_2816),
.Y(n_2831)
);

OR2x2_ASAP7_75t_L g2832 ( 
.A(n_2794),
.B(n_2765),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2801),
.B(n_2809),
.Y(n_2833)
);

INVx2_ASAP7_75t_L g2834 ( 
.A(n_2797),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2816),
.B(n_2819),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2815),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2803),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2800),
.B(n_2731),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2783),
.Y(n_2839)
);

INVxp67_ASAP7_75t_SL g2840 ( 
.A(n_2784),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2819),
.B(n_2745),
.Y(n_2841)
);

INVxp67_ASAP7_75t_SL g2842 ( 
.A(n_2784),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2793),
.Y(n_2843)
);

HB1xp67_ASAP7_75t_L g2844 ( 
.A(n_2788),
.Y(n_2844)
);

INVx2_ASAP7_75t_SL g2845 ( 
.A(n_2806),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2810),
.Y(n_2846)
);

INVx2_ASAP7_75t_SL g2847 ( 
.A(n_2806),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2810),
.Y(n_2848)
);

HB1xp67_ASAP7_75t_L g2849 ( 
.A(n_2788),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2800),
.B(n_2777),
.Y(n_2850)
);

NOR2xp67_ASAP7_75t_L g2851 ( 
.A(n_2806),
.B(n_2804),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2797),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2814),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2814),
.B(n_2782),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2785),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2789),
.B(n_2770),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2820),
.Y(n_2857)
);

NAND4xp25_ASAP7_75t_SL g2858 ( 
.A(n_2822),
.B(n_2776),
.C(n_2757),
.D(n_2726),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2850),
.B(n_2824),
.Y(n_2859)
);

AO21x2_ASAP7_75t_L g2860 ( 
.A1(n_2851),
.A2(n_2770),
.B(n_2779),
.Y(n_2860)
);

INVx1_ASAP7_75t_SL g2861 ( 
.A(n_2829),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2832),
.B(n_2787),
.Y(n_2862)
);

AOI221xp5_ASAP7_75t_L g2863 ( 
.A1(n_2833),
.A2(n_2739),
.B1(n_2766),
.B2(n_2760),
.C(n_2728),
.Y(n_2863)
);

AO21x2_ASAP7_75t_L g2864 ( 
.A1(n_2833),
.A2(n_2792),
.B(n_2791),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2856),
.B(n_2804),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2828),
.Y(n_2866)
);

AND2x4_ASAP7_75t_SL g2867 ( 
.A(n_2825),
.B(n_2805),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2856),
.B(n_2806),
.Y(n_2868)
);

INVx4_ASAP7_75t_L g2869 ( 
.A(n_2845),
.Y(n_2869)
);

AOI33xp33_ASAP7_75t_L g2870 ( 
.A1(n_2839),
.A2(n_2818),
.A3(n_2737),
.B1(n_2716),
.B2(n_2719),
.B3(n_2805),
.Y(n_2870)
);

HB1xp67_ASAP7_75t_L g2871 ( 
.A(n_2831),
.Y(n_2871)
);

OAI21x1_ASAP7_75t_L g2872 ( 
.A1(n_2835),
.A2(n_2808),
.B(n_2785),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2821),
.Y(n_2873)
);

BUFx3_ASAP7_75t_L g2874 ( 
.A(n_2847),
.Y(n_2874)
);

OAI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2823),
.A2(n_2818),
.B1(n_2728),
.B2(n_2807),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2834),
.Y(n_2876)
);

INVx2_ASAP7_75t_SL g2877 ( 
.A(n_2825),
.Y(n_2877)
);

AOI221xp5_ASAP7_75t_L g2878 ( 
.A1(n_2827),
.A2(n_2766),
.B1(n_2709),
.B2(n_2729),
.C(n_2769),
.Y(n_2878)
);

OAI21x1_ASAP7_75t_L g2879 ( 
.A1(n_2835),
.A2(n_2785),
.B(n_2792),
.Y(n_2879)
);

AOI222xp33_ASAP7_75t_L g2880 ( 
.A1(n_2843),
.A2(n_2811),
.B1(n_2711),
.B2(n_2729),
.C1(n_2817),
.C2(n_2717),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2852),
.Y(n_2881)
);

INVx3_ASAP7_75t_L g2882 ( 
.A(n_2855),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2838),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2836),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2844),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2826),
.B(n_2817),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2830),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2837),
.B(n_2811),
.Y(n_2888)
);

HB1xp67_ASAP7_75t_L g2889 ( 
.A(n_2844),
.Y(n_2889)
);

AOI21x1_ASAP7_75t_L g2890 ( 
.A1(n_2849),
.A2(n_2786),
.B(n_2791),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2846),
.Y(n_2891)
);

NOR2xp33_ASAP7_75t_L g2892 ( 
.A(n_2861),
.B(n_2841),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2889),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2889),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2859),
.B(n_2867),
.Y(n_2895)
);

OR2x2_ASAP7_75t_L g2896 ( 
.A(n_2862),
.B(n_2841),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2869),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2871),
.Y(n_2898)
);

INVxp67_ASAP7_75t_L g2899 ( 
.A(n_2871),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2867),
.B(n_2877),
.Y(n_2900)
);

OR2x2_ASAP7_75t_L g2901 ( 
.A(n_2888),
.B(n_2868),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2885),
.Y(n_2902)
);

OR2x6_ASAP7_75t_SL g2903 ( 
.A(n_2875),
.B(n_2735),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2886),
.B(n_2786),
.Y(n_2904)
);

AND2x2_ASAP7_75t_L g2905 ( 
.A(n_2886),
.B(n_2883),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2865),
.B(n_2840),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2869),
.B(n_2840),
.Y(n_2907)
);

OR2x2_ASAP7_75t_L g2908 ( 
.A(n_2864),
.B(n_2854),
.Y(n_2908)
);

AND3x2_ASAP7_75t_L g2909 ( 
.A(n_2863),
.B(n_2842),
.C(n_2717),
.Y(n_2909)
);

AND2x4_ASAP7_75t_SL g2910 ( 
.A(n_2865),
.B(n_2698),
.Y(n_2910)
);

OR2x2_ASAP7_75t_L g2911 ( 
.A(n_2864),
.B(n_2854),
.Y(n_2911)
);

OR2x2_ASAP7_75t_L g2912 ( 
.A(n_2874),
.B(n_2842),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2885),
.Y(n_2913)
);

INVx6_ASAP7_75t_L g2914 ( 
.A(n_2874),
.Y(n_2914)
);

NOR2x1p5_ASAP7_75t_L g2915 ( 
.A(n_2890),
.B(n_2848),
.Y(n_2915)
);

AND2x4_ASAP7_75t_SL g2916 ( 
.A(n_2882),
.B(n_2706),
.Y(n_2916)
);

INVx2_ASAP7_75t_SL g2917 ( 
.A(n_2860),
.Y(n_2917)
);

NOR2xp33_ASAP7_75t_L g2918 ( 
.A(n_2858),
.B(n_2715),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2891),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2891),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2857),
.Y(n_2921)
);

INVx3_ASAP7_75t_L g2922 ( 
.A(n_2860),
.Y(n_2922)
);

NOR2xp33_ASAP7_75t_L g2923 ( 
.A(n_2873),
.B(n_2853),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2884),
.Y(n_2924)
);

AOI22xp33_ASAP7_75t_L g2925 ( 
.A1(n_2863),
.A2(n_2738),
.B1(n_2718),
.B2(n_2740),
.Y(n_2925)
);

AOI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2878),
.A2(n_2738),
.B1(n_2718),
.B2(n_2700),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2887),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2876),
.B(n_2725),
.Y(n_2928)
);

NOR2x1_ASAP7_75t_R g2929 ( 
.A(n_2882),
.B(n_2736),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2881),
.B(n_2799),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2878),
.B(n_2775),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2866),
.B(n_2720),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2866),
.B(n_2720),
.Y(n_2933)
);

OR2x2_ASAP7_75t_L g2934 ( 
.A(n_2879),
.B(n_2733),
.Y(n_2934)
);

AOI21xp5_ASAP7_75t_L g2935 ( 
.A1(n_2880),
.A2(n_2707),
.B(n_2713),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2870),
.B(n_2733),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2870),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2893),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2893),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2895),
.B(n_2900),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2894),
.Y(n_2941)
);

HB1xp67_ASAP7_75t_L g2942 ( 
.A(n_2907),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2898),
.Y(n_2943)
);

HB1xp67_ASAP7_75t_L g2944 ( 
.A(n_2917),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2897),
.B(n_2872),
.Y(n_2945)
);

A2O1A1Ixp33_ASAP7_75t_L g2946 ( 
.A1(n_2937),
.A2(n_2676),
.B(n_2774),
.C(n_2700),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2919),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2937),
.B(n_2733),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2920),
.Y(n_2949)
);

HB1xp67_ASAP7_75t_L g2950 ( 
.A(n_2912),
.Y(n_2950)
);

INVx2_ASAP7_75t_L g2951 ( 
.A(n_2914),
.Y(n_2951)
);

HB1xp67_ASAP7_75t_L g2952 ( 
.A(n_2922),
.Y(n_2952)
);

OR2x2_ASAP7_75t_L g2953 ( 
.A(n_2896),
.B(n_2695),
.Y(n_2953)
);

INVx2_ASAP7_75t_L g2954 ( 
.A(n_2914),
.Y(n_2954)
);

OR2x2_ASAP7_75t_L g2955 ( 
.A(n_2906),
.B(n_2679),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2899),
.Y(n_2956)
);

NOR2x1p5_ASAP7_75t_SL g2957 ( 
.A(n_2908),
.B(n_2704),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2904),
.B(n_2680),
.Y(n_2958)
);

NOR2xp33_ASAP7_75t_L g2959 ( 
.A(n_2918),
.B(n_2734),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2916),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2892),
.B(n_2679),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2905),
.B(n_2688),
.Y(n_2962)
);

OR2x2_ASAP7_75t_L g2963 ( 
.A(n_2901),
.B(n_2688),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2910),
.B(n_2680),
.Y(n_2964)
);

NAND4xp25_ASAP7_75t_SL g2965 ( 
.A(n_2926),
.B(n_2705),
.C(n_2708),
.D(n_2703),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2902),
.Y(n_2966)
);

AND2x2_ASAP7_75t_L g2967 ( 
.A(n_2928),
.B(n_2713),
.Y(n_2967)
);

OAI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_2925),
.A2(n_46),
.B(n_47),
.Y(n_2968)
);

OAI22xp5_ASAP7_75t_L g2969 ( 
.A1(n_2903),
.A2(n_2708),
.B1(n_2699),
.B2(n_2697),
.Y(n_2969)
);

INVx1_ASAP7_75t_SL g2970 ( 
.A(n_2922),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2913),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2923),
.B(n_48),
.Y(n_2972)
);

AND2x2_ASAP7_75t_L g2973 ( 
.A(n_2930),
.B(n_48),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2929),
.Y(n_2974)
);

NAND3xp33_ASAP7_75t_L g2975 ( 
.A(n_2909),
.B(n_50),
.C(n_51),
.Y(n_2975)
);

OR2x6_ASAP7_75t_L g2976 ( 
.A(n_2915),
.B(n_50),
.Y(n_2976)
);

AND2x2_ASAP7_75t_L g2977 ( 
.A(n_2932),
.B(n_2933),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2921),
.B(n_51),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2924),
.B(n_52),
.Y(n_2979)
);

INVxp67_ASAP7_75t_L g2980 ( 
.A(n_2911),
.Y(n_2980)
);

OR2x2_ASAP7_75t_L g2981 ( 
.A(n_2931),
.B(n_53),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2927),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2934),
.B(n_53),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2936),
.B(n_54),
.Y(n_2984)
);

NAND2x1_ASAP7_75t_L g2985 ( 
.A(n_2935),
.B(n_54),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2893),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2893),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2893),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2893),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2893),
.Y(n_2990)
);

HB1xp67_ASAP7_75t_L g2991 ( 
.A(n_2907),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2897),
.B(n_57),
.Y(n_2992)
);

NAND2xp33_ASAP7_75t_SL g2993 ( 
.A(n_2895),
.B(n_57),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2893),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2897),
.B(n_58),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2893),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2897),
.B(n_58),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2893),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2893),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2893),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2897),
.B(n_59),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2893),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2893),
.Y(n_3003)
);

NOR2x1p5_ASAP7_75t_SL g3004 ( 
.A(n_2912),
.B(n_59),
.Y(n_3004)
);

HB1xp67_ASAP7_75t_L g3005 ( 
.A(n_2942),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2940),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2951),
.B(n_60),
.Y(n_3007)
);

AOI21xp5_ASAP7_75t_L g3008 ( 
.A1(n_2968),
.A2(n_61),
.B(n_62),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2954),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2950),
.Y(n_3010)
);

HB1xp67_ASAP7_75t_L g3011 ( 
.A(n_2991),
.Y(n_3011)
);

OR2x2_ASAP7_75t_L g3012 ( 
.A(n_2981),
.B(n_61),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2960),
.B(n_62),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2974),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2952),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2958),
.B(n_63),
.Y(n_3016)
);

OR2x2_ASAP7_75t_L g3017 ( 
.A(n_2956),
.B(n_63),
.Y(n_3017)
);

AND2x4_ASAP7_75t_L g3018 ( 
.A(n_3004),
.B(n_64),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2977),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2973),
.B(n_65),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2964),
.B(n_65),
.Y(n_3021)
);

NOR3xp33_ASAP7_75t_L g3022 ( 
.A(n_2975),
.B(n_66),
.C(n_67),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2984),
.B(n_66),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2976),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2944),
.Y(n_3025)
);

OAI33xp33_ASAP7_75t_L g3026 ( 
.A1(n_2980),
.A2(n_70),
.A3(n_72),
.B1(n_68),
.B2(n_69),
.B3(n_71),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2938),
.Y(n_3027)
);

AND2x2_ASAP7_75t_L g3028 ( 
.A(n_2959),
.B(n_68),
.Y(n_3028)
);

NOR4xp25_ASAP7_75t_SL g3029 ( 
.A(n_2993),
.B(n_2986),
.C(n_2987),
.D(n_2939),
.Y(n_3029)
);

NAND2xp33_ASAP7_75t_R g3030 ( 
.A(n_2976),
.B(n_70),
.Y(n_3030)
);

NOR2xp67_ASAP7_75t_L g3031 ( 
.A(n_2975),
.B(n_71),
.Y(n_3031)
);

HB1xp67_ASAP7_75t_L g3032 ( 
.A(n_2976),
.Y(n_3032)
);

BUFx2_ASAP7_75t_SL g3033 ( 
.A(n_2943),
.Y(n_3033)
);

NAND2xp33_ASAP7_75t_SL g3034 ( 
.A(n_2985),
.B(n_73),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2983),
.B(n_74),
.Y(n_3035)
);

OR2x2_ASAP7_75t_L g3036 ( 
.A(n_2992),
.B(n_75),
.Y(n_3036)
);

OR2x2_ASAP7_75t_L g3037 ( 
.A(n_2995),
.B(n_75),
.Y(n_3037)
);

OR2x2_ASAP7_75t_L g3038 ( 
.A(n_2997),
.B(n_76),
.Y(n_3038)
);

OR2x2_ASAP7_75t_L g3039 ( 
.A(n_3001),
.B(n_77),
.Y(n_3039)
);

NOR3xp33_ASAP7_75t_L g3040 ( 
.A(n_2968),
.B(n_78),
.C(n_79),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2978),
.B(n_79),
.Y(n_3041)
);

INVxp67_ASAP7_75t_L g3042 ( 
.A(n_2945),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2988),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_L g3044 ( 
.A(n_2979),
.B(n_80),
.Y(n_3044)
);

NAND3xp33_ASAP7_75t_L g3045 ( 
.A(n_2948),
.B(n_81),
.C(n_82),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2941),
.B(n_81),
.Y(n_3046)
);

NAND2xp33_ASAP7_75t_SL g3047 ( 
.A(n_2972),
.B(n_82),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2962),
.B(n_83),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2989),
.Y(n_3049)
);

OR2x6_ASAP7_75t_L g3050 ( 
.A(n_2990),
.B(n_2994),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2996),
.B(n_84),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2998),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2999),
.Y(n_3053)
);

OAI221xp5_ASAP7_75t_L g3054 ( 
.A1(n_2946),
.A2(n_88),
.B1(n_85),
.B2(n_86),
.C(n_89),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2961),
.B(n_85),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_3000),
.Y(n_3056)
);

NAND3xp33_ASAP7_75t_L g3057 ( 
.A(n_2966),
.B(n_2971),
.C(n_3002),
.Y(n_3057)
);

AND2x2_ASAP7_75t_L g3058 ( 
.A(n_2955),
.B(n_86),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_3003),
.B(n_90),
.Y(n_3059)
);

AND2x2_ASAP7_75t_L g3060 ( 
.A(n_2967),
.B(n_91),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2963),
.B(n_92),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2947),
.B(n_92),
.Y(n_3062)
);

OR2x4_ASAP7_75t_L g3063 ( 
.A(n_2982),
.B(n_93),
.Y(n_3063)
);

HB1xp67_ASAP7_75t_L g3064 ( 
.A(n_2970),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2970),
.Y(n_3065)
);

AOI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2965),
.A2(n_93),
.B(n_94),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_2949),
.B(n_95),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2953),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_2969),
.B(n_95),
.Y(n_3069)
);

AND4x1_ASAP7_75t_L g3070 ( 
.A(n_2957),
.B(n_98),
.C(n_96),
.D(n_97),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2950),
.Y(n_3071)
);

INVxp67_ASAP7_75t_SL g3072 ( 
.A(n_2942),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2950),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2950),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_2940),
.B(n_97),
.Y(n_3075)
);

NOR2x1_ASAP7_75t_L g3076 ( 
.A(n_2975),
.B(n_99),
.Y(n_3076)
);

AND2x2_ASAP7_75t_L g3077 ( 
.A(n_2940),
.B(n_100),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2940),
.B(n_101),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2950),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_2940),
.B(n_101),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2942),
.B(n_102),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2942),
.B(n_103),
.Y(n_3082)
);

INVx2_ASAP7_75t_SL g3083 ( 
.A(n_2951),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2950),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2940),
.B(n_103),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2942),
.B(n_104),
.Y(n_3086)
);

AND2x4_ASAP7_75t_L g3087 ( 
.A(n_2940),
.B(n_104),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2942),
.B(n_105),
.Y(n_3088)
);

NAND2xp33_ASAP7_75t_R g3089 ( 
.A(n_2976),
.B(n_105),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2950),
.Y(n_3090)
);

OAI211xp5_ASAP7_75t_L g3091 ( 
.A1(n_2975),
.A2(n_112),
.B(n_106),
.C(n_110),
.Y(n_3091)
);

OR2x2_ASAP7_75t_L g3092 ( 
.A(n_2942),
.B(n_106),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2950),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2942),
.B(n_112),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2942),
.B(n_113),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2952),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2952),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_3006),
.B(n_113),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_3005),
.Y(n_3099)
);

OAI22xp5_ASAP7_75t_L g3100 ( 
.A1(n_3029),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_3011),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_3072),
.Y(n_3102)
);

OR2x2_ASAP7_75t_L g3103 ( 
.A(n_3010),
.B(n_114),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_3064),
.Y(n_3104)
);

NAND3xp33_ASAP7_75t_L g3105 ( 
.A(n_3022),
.B(n_115),
.C(n_118),
.Y(n_3105)
);

OR2x2_ASAP7_75t_L g3106 ( 
.A(n_3071),
.B(n_119),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_3031),
.B(n_122),
.Y(n_3107)
);

NOR2xp33_ASAP7_75t_L g3108 ( 
.A(n_3024),
.B(n_122),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_3032),
.B(n_123),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_SL g3110 ( 
.A(n_3018),
.B(n_123),
.Y(n_3110)
);

OR2x2_ASAP7_75t_L g3111 ( 
.A(n_3073),
.B(n_127),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_3050),
.Y(n_3112)
);

OR2x2_ASAP7_75t_L g3113 ( 
.A(n_3074),
.B(n_128),
.Y(n_3113)
);

OR2x2_ASAP7_75t_L g3114 ( 
.A(n_3079),
.B(n_129),
.Y(n_3114)
);

INVxp67_ASAP7_75t_L g3115 ( 
.A(n_3030),
.Y(n_3115)
);

NOR2xp33_ASAP7_75t_SL g3116 ( 
.A(n_3076),
.B(n_129),
.Y(n_3116)
);

OR2x6_ASAP7_75t_L g3117 ( 
.A(n_3083),
.B(n_130),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_3050),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_3018),
.B(n_130),
.Y(n_3119)
);

AND2x2_ASAP7_75t_L g3120 ( 
.A(n_3075),
.B(n_132),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_3077),
.B(n_132),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_3078),
.B(n_133),
.Y(n_3122)
);

OR2x2_ASAP7_75t_L g3123 ( 
.A(n_3084),
.B(n_133),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_3087),
.B(n_134),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_3080),
.B(n_135),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_3085),
.B(n_135),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_3087),
.B(n_136),
.Y(n_3127)
);

NOR2xp33_ASAP7_75t_L g3128 ( 
.A(n_3063),
.B(n_137),
.Y(n_3128)
);

INVxp67_ASAP7_75t_SL g3129 ( 
.A(n_3089),
.Y(n_3129)
);

INVxp67_ASAP7_75t_L g3130 ( 
.A(n_3034),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_3097),
.Y(n_3131)
);

AND2x4_ASAP7_75t_L g3132 ( 
.A(n_3090),
.B(n_138),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_3014),
.B(n_139),
.Y(n_3133)
);

AOI221xp5_ASAP7_75t_L g3134 ( 
.A1(n_3054),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.C(n_142),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_3096),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_3096),
.Y(n_3136)
);

AOI21xp5_ASAP7_75t_L g3137 ( 
.A1(n_3008),
.A2(n_140),
.B(n_143),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_SL g3138 ( 
.A(n_3070),
.B(n_146),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_3097),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_3093),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_3065),
.Y(n_3141)
);

AND2x2_ASAP7_75t_L g3142 ( 
.A(n_3009),
.B(n_146),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3015),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_3019),
.B(n_147),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_3092),
.Y(n_3145)
);

INVxp67_ASAP7_75t_L g3146 ( 
.A(n_3033),
.Y(n_3146)
);

NOR2x1_ASAP7_75t_L g3147 ( 
.A(n_3045),
.B(n_148),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_3025),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_L g3149 ( 
.A(n_3042),
.B(n_149),
.Y(n_3149)
);

NOR3xp33_ASAP7_75t_L g3150 ( 
.A(n_3047),
.B(n_149),
.C(n_151),
.Y(n_3150)
);

OR2x2_ASAP7_75t_L g3151 ( 
.A(n_3081),
.B(n_3082),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3017),
.Y(n_3152)
);

AOI211xp5_ASAP7_75t_L g3153 ( 
.A1(n_3040),
.A2(n_154),
.B(n_151),
.C(n_153),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3020),
.Y(n_3154)
);

INVx1_ASAP7_75t_SL g3155 ( 
.A(n_3016),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_3035),
.Y(n_3156)
);

INVx1_ASAP7_75t_SL g3157 ( 
.A(n_3007),
.Y(n_3157)
);

INVx1_ASAP7_75t_SL g3158 ( 
.A(n_3012),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_3067),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_3013),
.B(n_154),
.Y(n_3160)
);

INVxp67_ASAP7_75t_L g3161 ( 
.A(n_3021),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3086),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_3060),
.B(n_155),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_3028),
.B(n_155),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_3055),
.B(n_157),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_3048),
.B(n_3061),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_3091),
.B(n_158),
.Y(n_3167)
);

OR2x2_ASAP7_75t_L g3168 ( 
.A(n_3088),
.B(n_158),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_3094),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_3095),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_3058),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_3068),
.B(n_160),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_3041),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_3023),
.B(n_160),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3044),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_3027),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_3036),
.B(n_3037),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_3038),
.B(n_162),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_3039),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3062),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_3043),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_3049),
.Y(n_3182)
);

AND5x1_ASAP7_75t_L g3183 ( 
.A(n_3066),
.B(n_167),
.C(n_164),
.D(n_165),
.E(n_168),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_3046),
.B(n_165),
.Y(n_3184)
);

OR2x2_ASAP7_75t_L g3185 ( 
.A(n_3051),
.B(n_168),
.Y(n_3185)
);

NOR2xp33_ASAP7_75t_L g3186 ( 
.A(n_3026),
.B(n_169),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_3052),
.Y(n_3187)
);

AND2x2_ASAP7_75t_L g3188 ( 
.A(n_3053),
.B(n_170),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3056),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_3059),
.B(n_170),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_3057),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_L g3192 ( 
.A(n_3069),
.B(n_172),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_3006),
.Y(n_3193)
);

NAND4xp25_ASAP7_75t_L g3194 ( 
.A(n_3014),
.B(n_175),
.C(n_173),
.D(n_174),
.Y(n_3194)
);

AND2x2_ASAP7_75t_L g3195 ( 
.A(n_3006),
.B(n_173),
.Y(n_3195)
);

CKINVDCx16_ASAP7_75t_R g3196 ( 
.A(n_3030),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_3072),
.B(n_174),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3005),
.Y(n_3198)
);

AOI22xp33_ASAP7_75t_SL g3199 ( 
.A1(n_3054),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_3199)
);

NOR2xp33_ASAP7_75t_L g3200 ( 
.A(n_3024),
.B(n_176),
.Y(n_3200)
);

AND2x2_ASAP7_75t_L g3201 ( 
.A(n_3006),
.B(n_178),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_3006),
.B(n_178),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_3006),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_3072),
.B(n_179),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3005),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_3005),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_3006),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3005),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3005),
.Y(n_3209)
);

CKINVDCx16_ASAP7_75t_R g3210 ( 
.A(n_3030),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_3006),
.Y(n_3211)
);

HB1xp67_ASAP7_75t_L g3212 ( 
.A(n_3005),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3005),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3005),
.Y(n_3214)
);

AND2x2_ASAP7_75t_L g3215 ( 
.A(n_3006),
.B(n_180),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_3006),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3072),
.B(n_180),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_3005),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_3072),
.B(n_181),
.Y(n_3219)
);

OR2x2_ASAP7_75t_L g3220 ( 
.A(n_3072),
.B(n_181),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3005),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3005),
.Y(n_3222)
);

AND4x1_ASAP7_75t_L g3223 ( 
.A(n_3076),
.B(n_184),
.C(n_182),
.D(n_183),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_3006),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3005),
.Y(n_3225)
);

NOR2x1_ASAP7_75t_L g3226 ( 
.A(n_3076),
.B(n_184),
.Y(n_3226)
);

INVx4_ASAP7_75t_L g3227 ( 
.A(n_3007),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_3072),
.B(n_185),
.Y(n_3228)
);

HB1xp67_ASAP7_75t_L g3229 ( 
.A(n_3005),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3072),
.B(n_185),
.Y(n_3230)
);

OR2x2_ASAP7_75t_L g3231 ( 
.A(n_3072),
.B(n_186),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3005),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_3006),
.B(n_186),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3072),
.B(n_187),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_3006),
.B(n_188),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3005),
.Y(n_3236)
);

INVx3_ASAP7_75t_L g3237 ( 
.A(n_3050),
.Y(n_3237)
);

NOR2xp33_ASAP7_75t_L g3238 ( 
.A(n_3024),
.B(n_189),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_3006),
.B(n_189),
.Y(n_3239)
);

AOI22xp33_ASAP7_75t_L g3240 ( 
.A1(n_3014),
.A2(n_193),
.B1(n_190),
.B2(n_191),
.Y(n_3240)
);

AND2x2_ASAP7_75t_L g3241 ( 
.A(n_3006),
.B(n_190),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_3072),
.B(n_191),
.Y(n_3242)
);

INVxp67_ASAP7_75t_L g3243 ( 
.A(n_3030),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_3005),
.Y(n_3244)
);

AND2x2_ASAP7_75t_L g3245 ( 
.A(n_3006),
.B(n_193),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_3006),
.B(n_194),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_3006),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_3006),
.B(n_195),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_3005),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_3006),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3072),
.B(n_196),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_3006),
.B(n_196),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_3006),
.B(n_199),
.Y(n_3253)
);

OAI21xp33_ASAP7_75t_L g3254 ( 
.A1(n_3129),
.A2(n_201),
.B(n_202),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3212),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_3196),
.B(n_3210),
.Y(n_3256)
);

INVx1_ASAP7_75t_SL g3257 ( 
.A(n_3226),
.Y(n_3257)
);

AOI222xp33_ASAP7_75t_L g3258 ( 
.A1(n_3100),
.A2(n_203),
.B1(n_205),
.B2(n_201),
.C1(n_202),
.C2(n_204),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3229),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3117),
.Y(n_3260)
);

AOI221xp5_ASAP7_75t_L g3261 ( 
.A1(n_3191),
.A2(n_3115),
.B1(n_3243),
.B2(n_3130),
.C(n_3104),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3117),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_3227),
.B(n_203),
.Y(n_3263)
);

NOR2x1_ASAP7_75t_L g3264 ( 
.A(n_3237),
.B(n_204),
.Y(n_3264)
);

O2A1O1Ixp33_ASAP7_75t_L g3265 ( 
.A1(n_3116),
.A2(n_211),
.B(n_206),
.C(n_210),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3209),
.Y(n_3266)
);

AND2x2_ASAP7_75t_L g3267 ( 
.A(n_3227),
.B(n_206),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3209),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3237),
.B(n_3146),
.Y(n_3269)
);

INVxp67_ASAP7_75t_L g3270 ( 
.A(n_3110),
.Y(n_3270)
);

OAI21xp33_ASAP7_75t_SL g3271 ( 
.A1(n_3102),
.A2(n_212),
.B(n_213),
.Y(n_3271)
);

INVx1_ASAP7_75t_SL g3272 ( 
.A(n_3155),
.Y(n_3272)
);

AOI221xp5_ASAP7_75t_L g3273 ( 
.A1(n_3101),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.C(n_216),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3220),
.Y(n_3274)
);

AOI221xp5_ASAP7_75t_L g3275 ( 
.A1(n_3198),
.A2(n_3208),
.B1(n_3213),
.B2(n_3206),
.C(n_3205),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3099),
.B(n_215),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_3166),
.B(n_216),
.Y(n_3277)
);

INVxp67_ASAP7_75t_L g3278 ( 
.A(n_3138),
.Y(n_3278)
);

AOI222xp33_ASAP7_75t_L g3279 ( 
.A1(n_3141),
.A2(n_219),
.B1(n_222),
.B2(n_217),
.C1(n_218),
.C2(n_221),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3231),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_3112),
.A2(n_223),
.B1(n_217),
.B2(n_222),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3214),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_3118),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3218),
.B(n_224),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_3157),
.B(n_224),
.Y(n_3285)
);

AOI221xp5_ASAP7_75t_L g3286 ( 
.A1(n_3221),
.A2(n_228),
.B1(n_225),
.B2(n_226),
.C(n_229),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_L g3287 ( 
.A(n_3223),
.B(n_226),
.Y(n_3287)
);

INVx1_ASAP7_75t_SL g3288 ( 
.A(n_3158),
.Y(n_3288)
);

A2O1A1Ixp33_ASAP7_75t_L g3289 ( 
.A1(n_3186),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3222),
.B(n_231),
.Y(n_3290)
);

OAI21xp33_ASAP7_75t_L g3291 ( 
.A1(n_3225),
.A2(n_3236),
.B(n_3232),
.Y(n_3291)
);

INVxp67_ASAP7_75t_L g3292 ( 
.A(n_3128),
.Y(n_3292)
);

AOI21xp33_ASAP7_75t_SL g3293 ( 
.A1(n_3244),
.A2(n_233),
.B(n_235),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_3132),
.Y(n_3294)
);

AOI22xp5_ASAP7_75t_L g3295 ( 
.A1(n_3161),
.A2(n_237),
.B1(n_233),
.B2(n_235),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3249),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3137),
.A2(n_237),
.B(n_238),
.Y(n_3297)
);

OAI322xp33_ASAP7_75t_L g3298 ( 
.A1(n_3140),
.A2(n_238),
.A3(n_239),
.B1(n_243),
.B2(n_244),
.C1(n_246),
.C2(n_247),
.Y(n_3298)
);

INVx1_ASAP7_75t_SL g3299 ( 
.A(n_3160),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_3171),
.B(n_239),
.Y(n_3300)
);

AOI32xp33_ASAP7_75t_L g3301 ( 
.A1(n_3147),
.A2(n_249),
.A3(n_243),
.B1(n_248),
.B2(n_250),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3178),
.B(n_249),
.Y(n_3302)
);

A2O1A1Ixp33_ASAP7_75t_SL g3303 ( 
.A1(n_3131),
.A2(n_252),
.B(n_250),
.C(n_251),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3132),
.Y(n_3304)
);

INVx2_ASAP7_75t_SL g3305 ( 
.A(n_3142),
.Y(n_3305)
);

OAI22xp5_ASAP7_75t_L g3306 ( 
.A1(n_3199),
.A2(n_3105),
.B1(n_3167),
.B2(n_3153),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3163),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_3145),
.B(n_3159),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3119),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_3165),
.B(n_253),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3120),
.Y(n_3311)
);

OAI21xp5_ASAP7_75t_SL g3312 ( 
.A1(n_3193),
.A2(n_253),
.B(n_254),
.Y(n_3312)
);

AOI221xp5_ASAP7_75t_L g3313 ( 
.A1(n_3148),
.A2(n_3143),
.B1(n_3135),
.B2(n_3139),
.C(n_3136),
.Y(n_3313)
);

HB1xp67_ASAP7_75t_L g3314 ( 
.A(n_3197),
.Y(n_3314)
);

AOI211xp5_ASAP7_75t_L g3315 ( 
.A1(n_3134),
.A2(n_257),
.B(n_254),
.C(n_255),
.Y(n_3315)
);

AOI222xp33_ASAP7_75t_L g3316 ( 
.A1(n_3149),
.A2(n_258),
.B1(n_263),
.B2(n_255),
.C1(n_257),
.C2(n_260),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3121),
.Y(n_3317)
);

AOI221xp5_ASAP7_75t_SL g3318 ( 
.A1(n_3203),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.C(n_266),
.Y(n_3318)
);

AND2x2_ASAP7_75t_L g3319 ( 
.A(n_3207),
.B(n_265),
.Y(n_3319)
);

OAI221xp5_ASAP7_75t_L g3320 ( 
.A1(n_3211),
.A2(n_270),
.B1(n_267),
.B2(n_269),
.C(n_271),
.Y(n_3320)
);

NOR2xp67_ASAP7_75t_L g3321 ( 
.A(n_3152),
.B(n_3216),
.Y(n_3321)
);

NAND3xp33_ASAP7_75t_L g3322 ( 
.A(n_3224),
.B(n_269),
.C(n_270),
.Y(n_3322)
);

AOI22xp5_ASAP7_75t_L g3323 ( 
.A1(n_3247),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_3323)
);

NAND2x1p5_ASAP7_75t_L g3324 ( 
.A(n_3122),
.B(n_3125),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3126),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_3250),
.B(n_272),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_3103),
.Y(n_3327)
);

OR2x2_ASAP7_75t_L g3328 ( 
.A(n_3109),
.B(n_3204),
.Y(n_3328)
);

INVxp67_ASAP7_75t_L g3329 ( 
.A(n_3192),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_3106),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3124),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3127),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3174),
.B(n_274),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3133),
.B(n_275),
.Y(n_3334)
);

NOR2x1p5_ASAP7_75t_L g3335 ( 
.A(n_3177),
.B(n_276),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_3098),
.B(n_276),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3144),
.Y(n_3337)
);

OAI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_3240),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_3338)
);

OAI31xp33_ASAP7_75t_L g3339 ( 
.A1(n_3150),
.A2(n_280),
.A3(n_277),
.B(n_278),
.Y(n_3339)
);

OAI22xp5_ASAP7_75t_L g3340 ( 
.A1(n_3151),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3195),
.Y(n_3341)
);

OR2x2_ASAP7_75t_L g3342 ( 
.A(n_3217),
.B(n_281),
.Y(n_3342)
);

OAI21xp33_ASAP7_75t_L g3343 ( 
.A1(n_3154),
.A2(n_282),
.B(n_285),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_3201),
.B(n_286),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3202),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3215),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_3111),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_3113),
.Y(n_3348)
);

INVxp67_ASAP7_75t_L g3349 ( 
.A(n_3108),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3233),
.B(n_287),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3235),
.Y(n_3351)
);

AOI321xp33_ASAP7_75t_L g3352 ( 
.A1(n_3179),
.A2(n_290),
.A3(n_292),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_3352)
);

AOI222xp33_ASAP7_75t_L g3353 ( 
.A1(n_3180),
.A2(n_290),
.B1(n_293),
.B2(n_288),
.C1(n_289),
.C2(n_291),
.Y(n_3353)
);

AOI22xp5_ASAP7_75t_L g3354 ( 
.A1(n_3200),
.A2(n_297),
.B1(n_293),
.B2(n_295),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3239),
.Y(n_3355)
);

OAI22xp5_ASAP7_75t_L g3356 ( 
.A1(n_3156),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_3356)
);

OAI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3219),
.A2(n_298),
.B(n_300),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3241),
.Y(n_3358)
);

XNOR2xp5_ASAP7_75t_L g3359 ( 
.A(n_3194),
.B(n_301),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3245),
.B(n_302),
.Y(n_3360)
);

OR2x2_ASAP7_75t_L g3361 ( 
.A(n_3228),
.B(n_303),
.Y(n_3361)
);

AOI21xp33_ASAP7_75t_L g3362 ( 
.A1(n_3162),
.A2(n_304),
.B(n_305),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3246),
.Y(n_3363)
);

OA21x2_ASAP7_75t_L g3364 ( 
.A1(n_3230),
.A2(n_306),
.B(n_307),
.Y(n_3364)
);

OAI21xp5_ASAP7_75t_SL g3365 ( 
.A1(n_3169),
.A2(n_306),
.B(n_307),
.Y(n_3365)
);

AOI22xp33_ASAP7_75t_L g3366 ( 
.A1(n_3173),
.A2(n_311),
.B1(n_308),
.B2(n_309),
.Y(n_3366)
);

OAI31xp33_ASAP7_75t_SL g3367 ( 
.A1(n_3181),
.A2(n_312),
.A3(n_308),
.B(n_309),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3248),
.B(n_312),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3252),
.Y(n_3369)
);

AOI221xp5_ASAP7_75t_L g3370 ( 
.A1(n_3187),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.C(n_316),
.Y(n_3370)
);

AOI222xp33_ASAP7_75t_L g3371 ( 
.A1(n_3170),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.C1(n_317),
.C2(n_318),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3114),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3253),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3175),
.B(n_317),
.Y(n_3374)
);

AOI221xp5_ASAP7_75t_L g3375 ( 
.A1(n_3189),
.A2(n_321),
.B1(n_318),
.B2(n_319),
.C(n_324),
.Y(n_3375)
);

HB1xp67_ASAP7_75t_L g3376 ( 
.A(n_3234),
.Y(n_3376)
);

INVxp67_ASAP7_75t_L g3377 ( 
.A(n_3238),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3107),
.B(n_324),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_SL g3379 ( 
.A(n_3257),
.B(n_3242),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_3324),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3256),
.B(n_3188),
.Y(n_3381)
);

INVx1_ASAP7_75t_SL g3382 ( 
.A(n_3288),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3294),
.B(n_3251),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3304),
.B(n_3182),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3260),
.B(n_3164),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_SL g3386 ( 
.A(n_3271),
.B(n_3123),
.Y(n_3386)
);

AND2x2_ASAP7_75t_L g3387 ( 
.A(n_3272),
.B(n_3172),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3264),
.Y(n_3388)
);

AND2x4_ASAP7_75t_L g3389 ( 
.A(n_3321),
.B(n_3176),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3263),
.Y(n_3390)
);

NOR2xp33_ASAP7_75t_L g3391 ( 
.A(n_3278),
.B(n_3168),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3262),
.B(n_3190),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3287),
.B(n_3184),
.Y(n_3393)
);

OAI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_3289),
.A2(n_3176),
.B(n_3185),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3267),
.B(n_3183),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3258),
.B(n_325),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3299),
.B(n_325),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_SL g3398 ( 
.A(n_3367),
.B(n_3255),
.Y(n_3398)
);

INVx1_ASAP7_75t_SL g3399 ( 
.A(n_3277),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3259),
.B(n_326),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3336),
.B(n_328),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3269),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3344),
.B(n_328),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_SL g3404 ( 
.A(n_3270),
.B(n_329),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3285),
.Y(n_3405)
);

AND2x4_ASAP7_75t_L g3406 ( 
.A(n_3335),
.B(n_329),
.Y(n_3406)
);

OR2x2_ASAP7_75t_L g3407 ( 
.A(n_3283),
.B(n_331),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3350),
.B(n_3274),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3307),
.B(n_331),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_3311),
.B(n_332),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_3325),
.Y(n_3411)
);

AOI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_3297),
.A2(n_335),
.B(n_336),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3280),
.B(n_335),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3300),
.Y(n_3414)
);

INVxp67_ASAP7_75t_L g3415 ( 
.A(n_3308),
.Y(n_3415)
);

HB1xp67_ASAP7_75t_L g3416 ( 
.A(n_3364),
.Y(n_3416)
);

HB1xp67_ASAP7_75t_L g3417 ( 
.A(n_3364),
.Y(n_3417)
);

BUFx2_ASAP7_75t_L g3418 ( 
.A(n_3266),
.Y(n_3418)
);

INVxp67_ASAP7_75t_L g3419 ( 
.A(n_3378),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3261),
.B(n_336),
.Y(n_3420)
);

INVxp67_ASAP7_75t_L g3421 ( 
.A(n_3319),
.Y(n_3421)
);

NOR3xp33_ASAP7_75t_L g3422 ( 
.A(n_3291),
.B(n_337),
.C(n_338),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_SL g3423 ( 
.A(n_3301),
.B(n_337),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3305),
.B(n_338),
.Y(n_3424)
);

OR2x2_ASAP7_75t_L g3425 ( 
.A(n_3317),
.B(n_339),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3326),
.Y(n_3426)
);

OAI31xp33_ASAP7_75t_L g3427 ( 
.A1(n_3303),
.A2(n_344),
.A3(n_340),
.B(n_341),
.Y(n_3427)
);

NOR2xp67_ASAP7_75t_L g3428 ( 
.A(n_3293),
.B(n_340),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3318),
.B(n_344),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3310),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3342),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3337),
.B(n_345),
.Y(n_3432)
);

OR2x2_ASAP7_75t_L g3433 ( 
.A(n_3341),
.B(n_348),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3268),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3345),
.B(n_349),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3346),
.B(n_350),
.Y(n_3436)
);

AND2x2_ASAP7_75t_L g3437 ( 
.A(n_3351),
.B(n_350),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3302),
.Y(n_3438)
);

OAI21xp5_ASAP7_75t_L g3439 ( 
.A1(n_3275),
.A2(n_351),
.B(n_352),
.Y(n_3439)
);

HB1xp67_ASAP7_75t_L g3440 ( 
.A(n_3327),
.Y(n_3440)
);

OR2x2_ASAP7_75t_L g3441 ( 
.A(n_3355),
.B(n_351),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3358),
.B(n_352),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3333),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3363),
.B(n_353),
.Y(n_3444)
);

NAND2x1_ASAP7_75t_L g3445 ( 
.A(n_3330),
.B(n_353),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3360),
.Y(n_3446)
);

NOR2xp33_ASAP7_75t_SL g3447 ( 
.A(n_3339),
.B(n_354),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3369),
.B(n_355),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3373),
.B(n_355),
.Y(n_3449)
);

OR2x2_ASAP7_75t_L g3450 ( 
.A(n_3276),
.B(n_356),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3316),
.B(n_356),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3279),
.B(n_357),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_SL g3453 ( 
.A(n_3352),
.B(n_3265),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3374),
.B(n_358),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3254),
.B(n_359),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3368),
.Y(n_3456)
);

AND2x4_ASAP7_75t_SL g3457 ( 
.A(n_3347),
.B(n_359),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3334),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3361),
.Y(n_3459)
);

OR2x2_ASAP7_75t_L g3460 ( 
.A(n_3348),
.B(n_360),
.Y(n_3460)
);

OR2x2_ASAP7_75t_L g3461 ( 
.A(n_3372),
.B(n_362),
.Y(n_3461)
);

INVxp67_ASAP7_75t_SL g3462 ( 
.A(n_3359),
.Y(n_3462)
);

AND2x4_ASAP7_75t_L g3463 ( 
.A(n_3282),
.B(n_3296),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3284),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3353),
.B(n_362),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3292),
.B(n_363),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3290),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3328),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3371),
.B(n_363),
.Y(n_3469)
);

INVxp67_ASAP7_75t_L g3470 ( 
.A(n_3314),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3376),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3309),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3309),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3331),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3332),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3349),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3312),
.B(n_364),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3365),
.B(n_365),
.Y(n_3478)
);

OR2x2_ASAP7_75t_L g3479 ( 
.A(n_3306),
.B(n_365),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_3377),
.B(n_366),
.Y(n_3480)
);

INVxp67_ASAP7_75t_L g3481 ( 
.A(n_3320),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3322),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3315),
.B(n_3313),
.Y(n_3483)
);

INVx3_ASAP7_75t_L g3484 ( 
.A(n_3362),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3356),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3329),
.B(n_367),
.Y(n_3486)
);

INVxp67_ASAP7_75t_L g3487 ( 
.A(n_3340),
.Y(n_3487)
);

AND2x2_ASAP7_75t_L g3488 ( 
.A(n_3357),
.B(n_367),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3323),
.Y(n_3489)
);

INVxp67_ASAP7_75t_L g3490 ( 
.A(n_3338),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3295),
.Y(n_3491)
);

AND2x4_ASAP7_75t_L g3492 ( 
.A(n_3354),
.B(n_368),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_SL g3493 ( 
.A(n_3273),
.B(n_368),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3343),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3286),
.B(n_369),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3281),
.B(n_370),
.Y(n_3496)
);

NAND2x1p5_ASAP7_75t_L g3497 ( 
.A(n_3298),
.B(n_371),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3366),
.B(n_371),
.Y(n_3498)
);

INVxp67_ASAP7_75t_SL g3499 ( 
.A(n_3370),
.Y(n_3499)
);

HB1xp67_ASAP7_75t_L g3500 ( 
.A(n_3375),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3256),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3324),
.B(n_372),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3257),
.B(n_372),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3283),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3257),
.B(n_373),
.Y(n_3505)
);

AND2x2_ASAP7_75t_L g3506 ( 
.A(n_3324),
.B(n_374),
.Y(n_3506)
);

OR2x2_ASAP7_75t_L g3507 ( 
.A(n_3256),
.B(n_377),
.Y(n_3507)
);

NAND3xp33_ASAP7_75t_L g3508 ( 
.A(n_3261),
.B(n_377),
.C(n_379),
.Y(n_3508)
);

OAI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_3256),
.A2(n_385),
.B1(n_379),
.B2(n_381),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3257),
.B(n_381),
.Y(n_3510)
);

OAI211xp5_ASAP7_75t_L g3511 ( 
.A1(n_3261),
.A2(n_388),
.B(n_385),
.C(n_387),
.Y(n_3511)
);

INVxp67_ASAP7_75t_L g3512 ( 
.A(n_3264),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3256),
.Y(n_3513)
);

INVx3_ASAP7_75t_L g3514 ( 
.A(n_3294),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3256),
.Y(n_3515)
);

NAND3xp33_ASAP7_75t_SL g3516 ( 
.A(n_3257),
.B(n_387),
.C(n_388),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3257),
.B(n_389),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3257),
.B(n_390),
.Y(n_3518)
);

XOR2xp5_ASAP7_75t_L g3519 ( 
.A(n_3359),
.B(n_390),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_SL g3520 ( 
.A(n_3257),
.B(n_391),
.Y(n_3520)
);

INVx1_ASAP7_75t_SL g3521 ( 
.A(n_3257),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3257),
.B(n_391),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3257),
.B(n_392),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3324),
.B(n_393),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3256),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3256),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_SL g3527 ( 
.A(n_3257),
.B(n_394),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3257),
.B(n_394),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3257),
.B(n_395),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3256),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3256),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3256),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3256),
.Y(n_3533)
);

AOI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3256),
.A2(n_396),
.B(n_398),
.Y(n_3534)
);

NAND2xp5_ASAP7_75t_L g3535 ( 
.A(n_3257),
.B(n_396),
.Y(n_3535)
);

AOI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3256),
.A2(n_398),
.B(n_399),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3256),
.Y(n_3537)
);

NAND3xp33_ASAP7_75t_L g3538 ( 
.A(n_3512),
.B(n_399),
.C(n_400),
.Y(n_3538)
);

NAND3xp33_ASAP7_75t_L g3539 ( 
.A(n_3388),
.B(n_400),
.C(n_401),
.Y(n_3539)
);

OAI21xp33_ASAP7_75t_L g3540 ( 
.A1(n_3382),
.A2(n_401),
.B(n_402),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3386),
.A2(n_402),
.B(n_403),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3514),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3416),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3417),
.Y(n_3544)
);

INVx4_ASAP7_75t_L g3545 ( 
.A(n_3514),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3389),
.Y(n_3546)
);

INVx2_ASAP7_75t_SL g3547 ( 
.A(n_3457),
.Y(n_3547)
);

AND2x4_ASAP7_75t_L g3548 ( 
.A(n_3389),
.B(n_403),
.Y(n_3548)
);

OR2x2_ASAP7_75t_L g3549 ( 
.A(n_3516),
.B(n_405),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3502),
.Y(n_3550)
);

XOR2x2_ASAP7_75t_L g3551 ( 
.A(n_3519),
.B(n_405),
.Y(n_3551)
);

NOR2xp33_ASAP7_75t_R g3552 ( 
.A(n_3404),
.B(n_406),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3506),
.Y(n_3553)
);

AND2x4_ASAP7_75t_L g3554 ( 
.A(n_3524),
.B(n_406),
.Y(n_3554)
);

INVxp67_ASAP7_75t_SL g3555 ( 
.A(n_3428),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3406),
.Y(n_3556)
);

NOR4xp25_ASAP7_75t_SL g3557 ( 
.A(n_3398),
.B(n_409),
.C(n_407),
.D(n_408),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3406),
.Y(n_3558)
);

AND2x2_ASAP7_75t_L g3559 ( 
.A(n_3521),
.B(n_407),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3445),
.Y(n_3560)
);

OAI321xp33_ASAP7_75t_L g3561 ( 
.A1(n_3483),
.A2(n_3415),
.A3(n_3501),
.B1(n_3525),
.B2(n_3515),
.C(n_3513),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3399),
.B(n_3390),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_3380),
.Y(n_3563)
);

O2A1O1Ixp33_ASAP7_75t_L g3564 ( 
.A1(n_3427),
.A2(n_411),
.B(n_409),
.C(n_410),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3440),
.Y(n_3565)
);

AND2x2_ASAP7_75t_L g3566 ( 
.A(n_3411),
.B(n_411),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_SL g3567 ( 
.A(n_3463),
.B(n_412),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3418),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3507),
.Y(n_3569)
);

NOR3xp33_ASAP7_75t_L g3570 ( 
.A(n_3526),
.B(n_413),
.C(n_414),
.Y(n_3570)
);

HB1xp67_ASAP7_75t_L g3571 ( 
.A(n_3463),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3503),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3381),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3505),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_3379),
.A2(n_414),
.B(n_415),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3409),
.B(n_3410),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3510),
.Y(n_3577)
);

AOI322xp5_ASAP7_75t_L g3578 ( 
.A1(n_3453),
.A2(n_415),
.A3(n_416),
.B1(n_417),
.B2(n_419),
.C1(n_420),
.C2(n_422),
.Y(n_3578)
);

XOR2x2_ASAP7_75t_L g3579 ( 
.A(n_3497),
.B(n_416),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3517),
.Y(n_3580)
);

AND2x2_ASAP7_75t_SL g3581 ( 
.A(n_3422),
.B(n_419),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3518),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3405),
.B(n_422),
.Y(n_3583)
);

INVx2_ASAP7_75t_SL g3584 ( 
.A(n_3407),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_SL g3585 ( 
.A(n_3447),
.B(n_423),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3522),
.Y(n_3586)
);

INVx1_ASAP7_75t_SL g3587 ( 
.A(n_3523),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3528),
.Y(n_3588)
);

OR2x2_ASAP7_75t_L g3589 ( 
.A(n_3395),
.B(n_423),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3387),
.B(n_425),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3529),
.Y(n_3591)
);

AOI22xp5_ASAP7_75t_L g3592 ( 
.A1(n_3530),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3535),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3425),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3384),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3433),
.Y(n_3596)
);

INVx2_ASAP7_75t_L g3597 ( 
.A(n_3441),
.Y(n_3597)
);

BUFx2_ASAP7_75t_L g3598 ( 
.A(n_3394),
.Y(n_3598)
);

INVxp33_ASAP7_75t_L g3599 ( 
.A(n_3391),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3531),
.B(n_427),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3437),
.Y(n_3601)
);

NOR2xp33_ASAP7_75t_L g3602 ( 
.A(n_3511),
.B(n_429),
.Y(n_3602)
);

AOI221xp5_ASAP7_75t_L g3603 ( 
.A1(n_3439),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.C(n_432),
.Y(n_3603)
);

BUFx2_ASAP7_75t_L g3604 ( 
.A(n_3444),
.Y(n_3604)
);

NOR3xp33_ASAP7_75t_SL g3605 ( 
.A(n_3532),
.B(n_433),
.C(n_434),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3408),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3533),
.B(n_434),
.Y(n_3607)
);

NOR4xp25_ASAP7_75t_SL g3608 ( 
.A(n_3423),
.B(n_437),
.C(n_435),
.D(n_436),
.Y(n_3608)
);

AOI221x1_ASAP7_75t_L g3609 ( 
.A1(n_3534),
.A2(n_437),
.B1(n_438),
.B2(n_441),
.C(n_442),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3460),
.Y(n_3610)
);

NOR3xp33_ASAP7_75t_L g3611 ( 
.A(n_3537),
.B(n_442),
.C(n_443),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3397),
.Y(n_3612)
);

CKINVDCx5p33_ASAP7_75t_R g3613 ( 
.A(n_3402),
.Y(n_3613)
);

INVx1_ASAP7_75t_SL g3614 ( 
.A(n_3479),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3383),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_3461),
.Y(n_3616)
);

INVx1_ASAP7_75t_SL g3617 ( 
.A(n_3520),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3414),
.B(n_443),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3426),
.B(n_444),
.Y(n_3619)
);

NOR2x1_ASAP7_75t_L g3620 ( 
.A(n_3508),
.B(n_444),
.Y(n_3620)
);

AND2x2_ASAP7_75t_L g3621 ( 
.A(n_3488),
.B(n_3485),
.Y(n_3621)
);

INVx4_ASAP7_75t_L g3622 ( 
.A(n_3476),
.Y(n_3622)
);

INVx1_ASAP7_75t_SL g3623 ( 
.A(n_3527),
.Y(n_3623)
);

AOI22xp5_ASAP7_75t_L g3624 ( 
.A1(n_3499),
.A2(n_447),
.B1(n_445),
.B2(n_446),
.Y(n_3624)
);

NOR4xp25_ASAP7_75t_L g3625 ( 
.A(n_3420),
.B(n_3487),
.C(n_3490),
.D(n_3482),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3401),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3421),
.B(n_445),
.Y(n_3627)
);

AND2x2_ASAP7_75t_L g3628 ( 
.A(n_3496),
.B(n_446),
.Y(n_3628)
);

INVx2_ASAP7_75t_SL g3629 ( 
.A(n_3471),
.Y(n_3629)
);

XNOR2xp5_ASAP7_75t_L g3630 ( 
.A(n_3500),
.B(n_447),
.Y(n_3630)
);

INVx2_ASAP7_75t_SL g3631 ( 
.A(n_3434),
.Y(n_3631)
);

XNOR2x1_ASAP7_75t_L g3632 ( 
.A(n_3494),
.B(n_448),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3403),
.Y(n_3633)
);

OAI211xp5_ASAP7_75t_SL g3634 ( 
.A1(n_3562),
.A2(n_3470),
.B(n_3481),
.C(n_3385),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3571),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3546),
.B(n_3536),
.Y(n_3636)
);

NOR2x1p5_ASAP7_75t_SL g3637 ( 
.A(n_3543),
.B(n_3491),
.Y(n_3637)
);

NOR3xp33_ASAP7_75t_L g3638 ( 
.A(n_3561),
.B(n_3392),
.C(n_3393),
.Y(n_3638)
);

NOR2x1_ASAP7_75t_SL g3639 ( 
.A(n_3545),
.B(n_3468),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3545),
.Y(n_3640)
);

NOR3xp33_ASAP7_75t_L g3641 ( 
.A(n_3598),
.B(n_3622),
.C(n_3558),
.Y(n_3641)
);

NOR2x1_ASAP7_75t_L g3642 ( 
.A(n_3544),
.B(n_3424),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3556),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3547),
.B(n_3412),
.Y(n_3644)
);

AOI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_3555),
.A2(n_3451),
.B(n_3429),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3560),
.B(n_3492),
.Y(n_3646)
);

NOR3xp33_ASAP7_75t_L g3647 ( 
.A(n_3622),
.B(n_3462),
.C(n_3484),
.Y(n_3647)
);

NOR3xp33_ASAP7_75t_L g3648 ( 
.A(n_3585),
.B(n_3484),
.C(n_3419),
.Y(n_3648)
);

AND4x1_ASAP7_75t_L g3649 ( 
.A(n_3625),
.B(n_3459),
.C(n_3438),
.D(n_3430),
.Y(n_3649)
);

NAND3x1_ASAP7_75t_L g3650 ( 
.A(n_3620),
.B(n_3478),
.C(n_3477),
.Y(n_3650)
);

NAND4xp75_ASAP7_75t_L g3651 ( 
.A(n_3565),
.B(n_3475),
.C(n_3474),
.D(n_3473),
.Y(n_3651)
);

A2O1A1Ixp33_ASAP7_75t_L g3652 ( 
.A1(n_3564),
.A2(n_3452),
.B(n_3469),
.C(n_3465),
.Y(n_3652)
);

AO21x1_ASAP7_75t_L g3653 ( 
.A1(n_3541),
.A2(n_3396),
.B(n_3400),
.Y(n_3653)
);

NOR4xp25_ASAP7_75t_L g3654 ( 
.A(n_3617),
.B(n_3472),
.C(n_3489),
.D(n_3467),
.Y(n_3654)
);

OAI22xp5_ASAP7_75t_L g3655 ( 
.A1(n_3599),
.A2(n_3495),
.B1(n_3455),
.B2(n_3498),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3559),
.Y(n_3656)
);

NOR3x1_ASAP7_75t_L g3657 ( 
.A(n_3604),
.B(n_3493),
.C(n_3413),
.Y(n_3657)
);

NOR2xp33_ASAP7_75t_L g3658 ( 
.A(n_3542),
.B(n_3454),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3554),
.B(n_3492),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3548),
.Y(n_3660)
);

OAI22xp5_ASAP7_75t_L g3661 ( 
.A1(n_3563),
.A2(n_3466),
.B1(n_3480),
.B2(n_3431),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_3568),
.B(n_3432),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3554),
.B(n_3443),
.Y(n_3663)
);

NOR2xp33_ASAP7_75t_L g3664 ( 
.A(n_3614),
.B(n_3435),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_SL g3665 ( 
.A(n_3552),
.B(n_3436),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3548),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3590),
.Y(n_3667)
);

NOR3x1_ASAP7_75t_L g3668 ( 
.A(n_3629),
.B(n_3448),
.C(n_3442),
.Y(n_3668)
);

INVx3_ASAP7_75t_L g3669 ( 
.A(n_3553),
.Y(n_3669)
);

AOI221xp5_ASAP7_75t_L g3670 ( 
.A1(n_3623),
.A2(n_3464),
.B1(n_3446),
.B2(n_3458),
.C(n_3456),
.Y(n_3670)
);

AOI211xp5_ASAP7_75t_L g3671 ( 
.A1(n_3589),
.A2(n_3509),
.B(n_3449),
.C(n_3486),
.Y(n_3671)
);

NAND5xp2_ASAP7_75t_L g3672 ( 
.A(n_3573),
.B(n_3504),
.C(n_3450),
.D(n_450),
.E(n_451),
.Y(n_3672)
);

OAI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_3575),
.A2(n_448),
.B(n_449),
.Y(n_3673)
);

NOR3xp33_ASAP7_75t_L g3674 ( 
.A(n_3606),
.B(n_449),
.C(n_450),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3630),
.Y(n_3675)
);

AND2x2_ASAP7_75t_L g3676 ( 
.A(n_3621),
.B(n_3550),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_SL g3677 ( 
.A(n_3549),
.B(n_451),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3566),
.Y(n_3678)
);

NAND4xp25_ASAP7_75t_L g3679 ( 
.A(n_3576),
.B(n_3601),
.C(n_3587),
.D(n_3595),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3618),
.Y(n_3680)
);

NAND3xp33_ASAP7_75t_SL g3681 ( 
.A(n_3557),
.B(n_452),
.C(n_455),
.Y(n_3681)
);

OAI221xp5_ASAP7_75t_L g3682 ( 
.A1(n_3631),
.A2(n_456),
.B1(n_457),
.B2(n_458),
.C(n_459),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3619),
.Y(n_3683)
);

NOR2xp67_ASAP7_75t_L g3684 ( 
.A(n_3539),
.B(n_456),
.Y(n_3684)
);

NOR2x1_ASAP7_75t_L g3685 ( 
.A(n_3538),
.B(n_458),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3608),
.B(n_459),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3627),
.Y(n_3687)
);

INVx1_ASAP7_75t_SL g3688 ( 
.A(n_3551),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_SL g3689 ( 
.A(n_3581),
.B(n_460),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3628),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3600),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_SL g3692 ( 
.A(n_3605),
.B(n_460),
.Y(n_3692)
);

NAND3xp33_ASAP7_75t_L g3693 ( 
.A(n_3609),
.B(n_461),
.C(n_462),
.Y(n_3693)
);

AOI22xp5_ASAP7_75t_L g3694 ( 
.A1(n_3613),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.Y(n_3694)
);

NOR2xp33_ASAP7_75t_L g3695 ( 
.A(n_3540),
.B(n_3567),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3632),
.Y(n_3696)
);

NAND4xp25_ASAP7_75t_L g3697 ( 
.A(n_3647),
.B(n_3569),
.C(n_3615),
.D(n_3577),
.Y(n_3697)
);

NOR3xp33_ASAP7_75t_L g3698 ( 
.A(n_3634),
.B(n_3584),
.C(n_3594),
.Y(n_3698)
);

NOR3xp33_ASAP7_75t_L g3699 ( 
.A(n_3679),
.B(n_3616),
.C(n_3610),
.Y(n_3699)
);

NOR2xp67_ASAP7_75t_L g3700 ( 
.A(n_3681),
.B(n_3596),
.Y(n_3700)
);

AOI221xp5_ASAP7_75t_L g3701 ( 
.A1(n_3654),
.A2(n_3591),
.B1(n_3588),
.B2(n_3574),
.C(n_3593),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3639),
.Y(n_3702)
);

NAND4xp75_ASAP7_75t_L g3703 ( 
.A(n_3637),
.B(n_3580),
.C(n_3586),
.D(n_3582),
.Y(n_3703)
);

AOI32xp33_ASAP7_75t_L g3704 ( 
.A1(n_3635),
.A2(n_3612),
.A3(n_3597),
.B1(n_3626),
.B2(n_3633),
.Y(n_3704)
);

NOR3xp33_ASAP7_75t_L g3705 ( 
.A(n_3641),
.B(n_3607),
.C(n_3572),
.Y(n_3705)
);

NAND4xp25_ASAP7_75t_L g3706 ( 
.A(n_3638),
.B(n_3603),
.C(n_3602),
.D(n_3583),
.Y(n_3706)
);

NAND4xp25_ASAP7_75t_SL g3707 ( 
.A(n_3670),
.B(n_3578),
.C(n_3611),
.D(n_3570),
.Y(n_3707)
);

AOI22xp5_ASAP7_75t_L g3708 ( 
.A1(n_3688),
.A2(n_3579),
.B1(n_3624),
.B2(n_3592),
.Y(n_3708)
);

NOR2x1_ASAP7_75t_L g3709 ( 
.A(n_3651),
.B(n_463),
.Y(n_3709)
);

NAND3xp33_ASAP7_75t_L g3710 ( 
.A(n_3693),
.B(n_464),
.C(n_465),
.Y(n_3710)
);

AOI211xp5_ASAP7_75t_L g3711 ( 
.A1(n_3672),
.A2(n_465),
.B(n_466),
.C(n_467),
.Y(n_3711)
);

OAI21xp33_ASAP7_75t_L g3712 ( 
.A1(n_3695),
.A2(n_466),
.B(n_467),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_SL g3713 ( 
.A(n_3686),
.B(n_468),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3660),
.B(n_468),
.Y(n_3714)
);

NOR3x1_ASAP7_75t_L g3715 ( 
.A(n_3673),
.B(n_470),
.C(n_471),
.Y(n_3715)
);

NOR2xp33_ASAP7_75t_L g3716 ( 
.A(n_3666),
.B(n_472),
.Y(n_3716)
);

AOI21xp33_ASAP7_75t_SL g3717 ( 
.A1(n_3659),
.A2(n_473),
.B(n_474),
.Y(n_3717)
);

AOI221xp5_ASAP7_75t_L g3718 ( 
.A1(n_3643),
.A2(n_473),
.B1(n_475),
.B2(n_476),
.C(n_477),
.Y(n_3718)
);

NOR4xp25_ASAP7_75t_L g3719 ( 
.A(n_3652),
.B(n_475),
.C(n_476),
.D(n_478),
.Y(n_3719)
);

NAND2xp33_ASAP7_75t_L g3720 ( 
.A(n_3674),
.B(n_479),
.Y(n_3720)
);

NAND4xp75_ASAP7_75t_L g3721 ( 
.A(n_3668),
.B(n_479),
.C(n_480),
.D(n_481),
.Y(n_3721)
);

OAI21xp33_ASAP7_75t_SL g3722 ( 
.A1(n_3640),
.A2(n_480),
.B(n_481),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3646),
.Y(n_3723)
);

NAND4xp25_ASAP7_75t_L g3724 ( 
.A(n_3657),
.B(n_482),
.C(n_483),
.D(n_484),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3676),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3669),
.B(n_3667),
.Y(n_3726)
);

NAND3xp33_ASAP7_75t_SL g3727 ( 
.A(n_3649),
.B(n_482),
.C(n_484),
.Y(n_3727)
);

NOR2x1p5_ASAP7_75t_L g3728 ( 
.A(n_3669),
.B(n_485),
.Y(n_3728)
);

NOR3xp33_ASAP7_75t_SL g3729 ( 
.A(n_3655),
.B(n_485),
.C(n_486),
.Y(n_3729)
);

NOR2x1_ASAP7_75t_L g3730 ( 
.A(n_3642),
.B(n_488),
.Y(n_3730)
);

NAND5xp2_ASAP7_75t_L g3731 ( 
.A(n_3645),
.B(n_489),
.C(n_490),
.D(n_491),
.E(n_493),
.Y(n_3731)
);

AOI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3648),
.A2(n_489),
.B1(n_491),
.B2(n_494),
.Y(n_3732)
);

NAND3xp33_ASAP7_75t_SL g3733 ( 
.A(n_3671),
.B(n_495),
.C(n_496),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3730),
.Y(n_3734)
);

AOI21xp5_ASAP7_75t_SL g3735 ( 
.A1(n_3713),
.A2(n_3689),
.B(n_3636),
.Y(n_3735)
);

AND2x2_ASAP7_75t_L g3736 ( 
.A(n_3725),
.B(n_3690),
.Y(n_3736)
);

INVxp67_ASAP7_75t_L g3737 ( 
.A(n_3731),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3728),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3700),
.B(n_3680),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3726),
.Y(n_3740)
);

AOI22x1_ASAP7_75t_L g3741 ( 
.A1(n_3702),
.A2(n_3687),
.B1(n_3656),
.B2(n_3683),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3719),
.B(n_3691),
.Y(n_3742)
);

OAI322xp33_ASAP7_75t_L g3743 ( 
.A1(n_3708),
.A2(n_3662),
.A3(n_3644),
.B1(n_3675),
.B2(n_3696),
.C1(n_3664),
.C2(n_3665),
.Y(n_3743)
);

NOR3xp33_ASAP7_75t_L g3744 ( 
.A(n_3706),
.B(n_3661),
.C(n_3663),
.Y(n_3744)
);

NAND2x1p5_ASAP7_75t_L g3745 ( 
.A(n_3709),
.B(n_3678),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3720),
.A2(n_3677),
.B(n_3692),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3714),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3721),
.Y(n_3748)
);

NOR2xp33_ASAP7_75t_L g3749 ( 
.A(n_3727),
.B(n_3653),
.Y(n_3749)
);

NAND3xp33_ASAP7_75t_L g3750 ( 
.A(n_3711),
.B(n_3685),
.C(n_3658),
.Y(n_3750)
);

NOR2x1_ASAP7_75t_L g3751 ( 
.A(n_3703),
.B(n_3682),
.Y(n_3751)
);

OAI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_3710),
.A2(n_3684),
.B1(n_3650),
.B2(n_3694),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3745),
.Y(n_3753)
);

NOR2x1_ASAP7_75t_L g3754 ( 
.A(n_3734),
.B(n_3724),
.Y(n_3754)
);

AOI21xp33_ASAP7_75t_SL g3755 ( 
.A1(n_3749),
.A2(n_3698),
.B(n_3699),
.Y(n_3755)
);

OAI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3751),
.A2(n_3722),
.B(n_3733),
.Y(n_3756)
);

NAND3xp33_ASAP7_75t_L g3757 ( 
.A(n_3744),
.B(n_3729),
.C(n_3701),
.Y(n_3757)
);

NOR2xp33_ASAP7_75t_L g3758 ( 
.A(n_3737),
.B(n_3712),
.Y(n_3758)
);

OAI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_3750),
.A2(n_3746),
.B(n_3739),
.Y(n_3759)
);

INVx1_ASAP7_75t_SL g3760 ( 
.A(n_3742),
.Y(n_3760)
);

NAND4xp75_ASAP7_75t_L g3761 ( 
.A(n_3736),
.B(n_3723),
.C(n_3715),
.D(n_3732),
.Y(n_3761)
);

OA21x2_ASAP7_75t_L g3762 ( 
.A1(n_3741),
.A2(n_3697),
.B(n_3705),
.Y(n_3762)
);

NAND4xp25_ASAP7_75t_L g3763 ( 
.A(n_3748),
.B(n_3704),
.C(n_3716),
.D(n_3718),
.Y(n_3763)
);

NOR3x2_ASAP7_75t_L g3764 ( 
.A(n_3735),
.B(n_3717),
.C(n_3707),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3738),
.Y(n_3765)
);

NAND3xp33_ASAP7_75t_L g3766 ( 
.A(n_3755),
.B(n_3740),
.C(n_3752),
.Y(n_3766)
);

NAND2x1p5_ASAP7_75t_L g3767 ( 
.A(n_3753),
.B(n_3747),
.Y(n_3767)
);

OAI22xp33_ASAP7_75t_SL g3768 ( 
.A1(n_3760),
.A2(n_3765),
.B1(n_3756),
.B2(n_3754),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3762),
.B(n_3743),
.Y(n_3769)
);

AOI22xp5_ASAP7_75t_L g3770 ( 
.A1(n_3757),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_3770)
);

NOR2xp67_ASAP7_75t_L g3771 ( 
.A(n_3763),
.B(n_497),
.Y(n_3771)
);

NOR2xp33_ASAP7_75t_L g3772 ( 
.A(n_3761),
.B(n_498),
.Y(n_3772)
);

INVxp67_ASAP7_75t_L g3773 ( 
.A(n_3758),
.Y(n_3773)
);

NAND3xp33_ASAP7_75t_SL g3774 ( 
.A(n_3759),
.B(n_499),
.C(n_500),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3764),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3769),
.Y(n_3776)
);

XNOR2xp5_ASAP7_75t_L g3777 ( 
.A(n_3766),
.B(n_3762),
.Y(n_3777)
);

INVx3_ASAP7_75t_L g3778 ( 
.A(n_3767),
.Y(n_3778)
);

NOR3xp33_ASAP7_75t_SL g3779 ( 
.A(n_3772),
.B(n_500),
.C(n_501),
.Y(n_3779)
);

AO22x1_ASAP7_75t_L g3780 ( 
.A1(n_3775),
.A2(n_502),
.B1(n_503),
.B2(n_504),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3778),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3777),
.A2(n_3768),
.B(n_3774),
.Y(n_3782)
);

OAI22xp5_ASAP7_75t_L g3783 ( 
.A1(n_3776),
.A2(n_3771),
.B1(n_3770),
.B2(n_3773),
.Y(n_3783)
);

AOI221xp5_ASAP7_75t_SL g3784 ( 
.A1(n_3779),
.A2(n_502),
.B1(n_504),
.B2(n_505),
.C(n_506),
.Y(n_3784)
);

AOI221x1_ASAP7_75t_L g3785 ( 
.A1(n_3782),
.A2(n_3783),
.B1(n_3781),
.B2(n_3784),
.C(n_3780),
.Y(n_3785)
);

AOI22xp5_ASAP7_75t_L g3786 ( 
.A1(n_3785),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_3786)
);

OAI21xp33_ASAP7_75t_L g3787 ( 
.A1(n_3786),
.A2(n_507),
.B(n_508),
.Y(n_3787)
);

AOI22xp5_ASAP7_75t_L g3788 ( 
.A1(n_3787),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.Y(n_3788)
);

BUFx2_ASAP7_75t_L g3789 ( 
.A(n_3788),
.Y(n_3789)
);

OAI22xp5_ASAP7_75t_L g3790 ( 
.A1(n_3789),
.A2(n_509),
.B1(n_512),
.B2(n_513),
.Y(n_3790)
);

AOI22xp5_ASAP7_75t_L g3791 ( 
.A1(n_3790),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_3791)
);

INVxp67_ASAP7_75t_SL g3792 ( 
.A(n_3791),
.Y(n_3792)
);

OR2x6_ASAP7_75t_L g3793 ( 
.A(n_3792),
.B(n_514),
.Y(n_3793)
);

AOI221xp5_ASAP7_75t_L g3794 ( 
.A1(n_3793),
.A2(n_515),
.B1(n_516),
.B2(n_518),
.C(n_519),
.Y(n_3794)
);

AOI211xp5_ASAP7_75t_L g3795 ( 
.A1(n_3794),
.A2(n_520),
.B(n_521),
.C(n_522),
.Y(n_3795)
);


endmodule