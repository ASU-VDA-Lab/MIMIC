module fake_jpeg_4338_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_43),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_41),
.B(n_42),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_46),
.Y(n_79)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_60),
.Y(n_91)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_62),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_50),
.B(n_52),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g58 ( 
.A(n_19),
.Y(n_58)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_38),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_15),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_59),
.Y(n_109)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_67),
.Y(n_124)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_39),
.B1(n_36),
.B2(n_34),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_68),
.A2(n_71),
.B1(n_89),
.B2(n_90),
.Y(n_142)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_75),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_39),
.B1(n_36),
.B2(n_23),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_29),
.B1(n_23),
.B2(n_32),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_73),
.A2(n_74),
.B1(n_93),
.B2(n_95),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_54),
.A2(n_26),
.B1(n_32),
.B2(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_85),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_78),
.A2(n_80),
.B1(n_82),
.B2(n_86),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_30),
.B1(n_31),
.B2(n_25),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_28),
.B1(n_37),
.B2(n_33),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g140 ( 
.A1(n_81),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_37),
.B1(n_24),
.B2(n_33),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_91),
.Y(n_115)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_28),
.B1(n_37),
.B2(n_33),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_31),
.B1(n_25),
.B2(n_28),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_24),
.B1(n_31),
.B2(n_25),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_38),
.B1(n_19),
.B2(n_21),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_40),
.A2(n_38),
.B1(n_19),
.B2(n_21),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_96),
.B(n_98),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_40),
.A2(n_38),
.B1(n_19),
.B2(n_21),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_107),
.B1(n_8),
.B2(n_13),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_57),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_106),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_44),
.A2(n_38),
.B1(n_35),
.B2(n_2),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_9),
.B(n_13),
.C(n_12),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_11),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_55),
.A2(n_63),
.B1(n_59),
.B2(n_3),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_46),
.Y(n_111)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_78),
.B(n_11),
.Y(n_146)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_115),
.B(n_133),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_116),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_0),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_118),
.A2(n_135),
.B(n_143),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_64),
.B1(n_72),
.B2(n_92),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_81),
.A2(n_14),
.B1(n_7),
.B2(n_10),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_66),
.B1(n_72),
.B2(n_67),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_132),
.Y(n_161)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_128),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_1),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_69),
.B(n_7),
.Y(n_133)
);

OR2x4_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_10),
.Y(n_135)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_88),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_105),
.B1(n_76),
.B2(n_80),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_102),
.B(n_1),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_83),
.B(n_3),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_3),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_147),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_156),
.Y(n_189)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_152),
.Y(n_181)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_151),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_136),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_153),
.B(n_154),
.Y(n_211)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_82),
.B1(n_110),
.B2(n_86),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_155),
.A2(n_158),
.B1(n_163),
.B2(n_113),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_103),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_112),
.B(n_85),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_65),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_142),
.B1(n_140),
.B2(n_130),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_159),
.B(n_162),
.Y(n_204)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_141),
.B1(n_138),
.B2(n_118),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_164),
.B(n_167),
.Y(n_212)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_166),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_75),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_174),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_143),
.B1(n_65),
.B2(n_88),
.Y(n_199)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_111),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_87),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_87),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_129),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_188),
.B1(n_194),
.B2(n_199),
.Y(n_223)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_201),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_118),
.B1(n_116),
.B2(n_126),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_143),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_190),
.A2(n_207),
.B(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_193),
.B(n_195),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_99),
.B1(n_114),
.B2(n_117),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_87),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_178),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_64),
.C(n_77),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_151),
.C(n_148),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_214),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_117),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_150),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_206),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_77),
.Y(n_206)
);

OR2x6_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_121),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_12),
.B1(n_121),
.B2(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_209),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_165),
.A2(n_146),
.B1(n_157),
.B2(n_174),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_213),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_150),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_229),
.C(n_238),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_SL g217 ( 
.A(n_189),
.B(n_146),
.C(n_160),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_222),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_237),
.B(n_207),
.Y(n_252)
);

AOI221xp5_ASAP7_75t_L g219 ( 
.A1(n_213),
.A2(n_160),
.B1(n_159),
.B2(n_178),
.C(n_173),
.Y(n_219)
);

NOR4xp25_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_185),
.C(n_190),
.D(n_209),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_227),
.Y(n_250)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_228),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_186),
.B(n_152),
.C(n_180),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_235),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_203),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_173),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_236),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_192),
.B(n_189),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_169),
.C(n_162),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_169),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_182),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_215),
.A2(n_188),
.B1(n_207),
.B2(n_199),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_244),
.A2(n_220),
.B1(n_223),
.B2(n_226),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_207),
.B1(n_201),
.B2(n_190),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_252),
.B(n_255),
.Y(n_271)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_210),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_225),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_256),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_254),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_259),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_222),
.Y(n_264)
);

NAND2xp33_ASAP7_75t_SL g259 ( 
.A(n_218),
.B(n_204),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_252),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_255),
.C(n_257),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_215),
.B(n_237),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_233),
.C(n_235),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_262),
.B(n_263),
.C(n_273),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_233),
.C(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_251),
.B1(n_248),
.B2(n_211),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_244),
.A2(n_231),
.B(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_216),
.C(n_229),
.Y(n_273)
);

OA22x2_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_194),
.B1(n_217),
.B2(n_232),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_271),
.B1(n_266),
.B2(n_260),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_230),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_241),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_270),
.B(n_249),
.Y(n_276)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_260),
.B(n_261),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_279),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_284),
.B1(n_274),
.B2(n_258),
.Y(n_298)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_267),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_285),
.C(n_287),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_185),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_221),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_241),
.B1(n_243),
.B2(n_246),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_212),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_262),
.C(n_263),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_292),
.B(n_294),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_273),
.C(n_271),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_285),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_260),
.C(n_268),
.Y(n_294)
);

AOI22x1_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_274),
.B1(n_253),
.B2(n_254),
.Y(n_295)
);

OAI321xp33_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_278),
.A3(n_289),
.B1(n_254),
.B2(n_242),
.C(n_224),
.Y(n_308)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_288),
.A2(n_274),
.B1(n_253),
.B2(n_236),
.Y(n_299)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_300),
.B(n_301),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_283),
.A2(n_181),
.B1(n_184),
.B2(n_191),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_307),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_287),
.Y(n_307)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_308),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_203),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_309),
.B(n_291),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_295),
.B1(n_294),
.B2(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_310),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_311),
.A2(n_313),
.B1(n_290),
.B2(n_242),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_297),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_307),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_318),
.A3(n_315),
.B1(n_303),
.B2(n_312),
.C1(n_310),
.C2(n_317),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_316),
.A2(n_304),
.A3(n_309),
.B1(n_290),
.B2(n_187),
.C1(n_202),
.C2(n_162),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_321),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_172),
.C(n_179),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_172),
.Y(n_324)
);


endmodule