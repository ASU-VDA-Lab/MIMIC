module real_jpeg_1015_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_43;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_40;
wire n_39;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_0),
.B(n_13),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_0),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_0),
.B(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

OR2x4_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_1),
.B(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_2),
.A2(n_14),
.B(n_15),
.Y(n_13)
);

AO21x1_ASAP7_75t_L g22 ( 
.A1(n_2),
.A2(n_23),
.B(n_24),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_2),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_4),
.Y(n_15)
);

OAI221xp5_ASAP7_75t_L g39 ( 
.A1(n_3),
.A2(n_13),
.B1(n_40),
.B2(n_42),
.C(n_43),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_10),
.Y(n_9)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

AOI211xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_11),
.B(n_16),
.C(n_39),
.Y(n_7)
);

INVx1_ASAP7_75t_SL g8 ( 
.A(n_9),
.Y(n_8)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_10),
.B(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

OAI221xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.C(n_28),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_19),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);


endmodule