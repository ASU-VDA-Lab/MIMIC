module fake_jpeg_22960_n_220 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_220);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx9p33_ASAP7_75t_R g67 ( 
.A(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_44),
.Y(n_47)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_17),
.Y(n_55)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_32),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_50),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_39),
.B1(n_37),
.B2(n_44),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_60),
.B1(n_66),
.B2(n_24),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_61),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_59),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_26),
.B1(n_31),
.B2(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_68),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_35),
.A2(n_32),
.B1(n_26),
.B2(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_22),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_2),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_22),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_98),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_77),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_25),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_86),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_39),
.B1(n_37),
.B2(n_50),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_62),
.B1(n_67),
.B2(n_18),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_25),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_29),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_21),
.Y(n_90)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_92),
.Y(n_115)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_45),
.B1(n_62),
.B2(n_33),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_24),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_100),
.Y(n_116)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_99),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_41),
.A3(n_36),
.B1(n_18),
.B2(n_25),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_41),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_108),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_16),
.B(n_23),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_126),
.B(n_82),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_41),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_82),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_110),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_71),
.B(n_45),
.Y(n_117)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_48),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_75),
.B(n_13),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_3),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_7),
.B(n_8),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_48),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_76),
.B(n_11),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_36),
.B(n_5),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_98),
.A3(n_87),
.B1(n_96),
.B2(n_74),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_87),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_130),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_135),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_138),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_73),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_73),
.B(n_67),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_142),
.B(n_144),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_85),
.B1(n_78),
.B2(n_11),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_145),
.B1(n_148),
.B2(n_109),
.Y(n_155)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_107),
.B1(n_101),
.B2(n_110),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_3),
.C(n_5),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_150),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_122),
.B1(n_107),
.B2(n_109),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_102),
.B1(n_104),
.B2(n_103),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_8),
.Y(n_149)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_106),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_153),
.Y(n_172)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_142),
.B1(n_150),
.B2(n_149),
.C(n_144),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_160),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_165),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_134),
.B1(n_128),
.B2(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_135),
.C(n_131),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_164),
.C(n_137),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_170),
.A2(n_174),
.B1(n_152),
.B2(n_154),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_177),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_155),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_103),
.C(n_138),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_154),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_158),
.C(n_167),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_187),
.C(n_192),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_185),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_160),
.B(n_162),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_152),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_172),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_191),
.B1(n_171),
.B2(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_154),
.B1(n_163),
.B2(n_156),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_147),
.B1(n_116),
.B2(n_123),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_164),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_192),
.C(n_187),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_198),
.C(n_113),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_171),
.C(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_201),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_175),
.B1(n_188),
.B2(n_185),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_179),
.B1(n_164),
.B2(n_139),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_176),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_204),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_194),
.C(n_202),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_206),
.A2(n_196),
.B(n_198),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_115),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_207),
.B(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_211),
.A2(n_206),
.B(n_207),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_112),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_212),
.B(n_204),
.Y(n_215)
);

AOI211xp5_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_112),
.B(n_123),
.C(n_147),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

AOI321xp33_ASAP7_75t_SL g218 ( 
.A1(n_216),
.A2(n_9),
.A3(n_10),
.B1(n_105),
.B2(n_173),
.C(n_210),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_218),
.Y(n_220)
);


endmodule