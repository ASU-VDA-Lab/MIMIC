module real_jpeg_23140_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_0),
.A2(n_26),
.B1(n_39),
.B2(n_43),
.Y(n_83)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g57 ( 
.A(n_4),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_39),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_5),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_46),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_5),
.A2(n_58),
.B(n_103),
.C(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_5),
.A2(n_46),
.B1(n_66),
.B2(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_53),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_55),
.B(n_73),
.C(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_5),
.B(n_24),
.C(n_42),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_5),
.B(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_5),
.B(n_44),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_7),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_7),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_7),
.A2(n_39),
.B1(n_43),
.B2(n_62),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_62),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_34),
.B1(n_39),
.B2(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_34),
.B1(n_61),
.B2(n_67),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_34),
.B1(n_54),
.B2(n_55),
.Y(n_126)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_132),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_130),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_108),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_15),
.B(n_108),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_91),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_79),
.B2(n_80),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_49),
.B2(n_50),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_35),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_35),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_29),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_22),
.A2(n_90),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_23),
.A2(n_24),
.B1(n_41),
.B2(n_42),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_24),
.B(n_196),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_27),
.B(n_33),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_27),
.B(n_89),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_27),
.A2(n_28),
.B(n_89),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_27),
.B(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_28),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_30),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_30),
.B(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_47),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_36),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_45),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_37),
.B(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_37),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_44),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_39),
.A2(n_43),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_39),
.B(n_172),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_43),
.A2(n_46),
.B(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_44),
.B(n_152),
.Y(n_169)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_46),
.A2(n_55),
.B(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_47),
.B(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_69),
.B1(n_70),
.B2(n_78),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_63),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_52),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_68),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_55),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_64),
.Y(n_95)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_119),
.Y(n_118)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B(n_76),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_71),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_71),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_75),
.B(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_77),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_82),
.B(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_84),
.B(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_86),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_90),
.B(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_101),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_106),
.Y(n_157)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_114),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_109),
.A2(n_110),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_230),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_113),
.Y(n_230)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_124),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_117),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_128),
.B(n_212),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_231),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_225),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_163),
.B(n_224),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_153),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_136),
.B(n_153),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.C(n_148),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_137),
.B(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_140),
.C(n_142),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_141),
.B(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_144),
.B(n_148),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_145),
.A2(n_147),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_145),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_147),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_156),
.B(n_157),
.C(n_158),
.Y(n_226)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_219),
.B(n_223),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_207),
.B(n_218),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_186),
.B(n_206),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_167),
.B(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_170),
.B1(n_171),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_180),
.B2(n_185),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_179),
.C(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_193),
.B(n_205),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_188),
.B(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_201),
.B(n_204),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);


endmodule