module fake_jpeg_2165_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_45),
.B(n_46),
.Y(n_110)
);

OR2x2_ASAP7_75t_SL g46 ( 
.A(n_25),
.B(n_0),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_19),
.B(n_2),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_54),
.B(n_71),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_11),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_12),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_78),
.Y(n_88)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_15),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_77),
.Y(n_103)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_34),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_4),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_19),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_82),
.Y(n_94)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_29),
.Y(n_95)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_25),
.C(n_40),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_45),
.B(n_37),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_73),
.C(n_37),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_28),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_28),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_52),
.A2(n_29),
.B1(n_42),
.B2(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_115),
.A2(n_129),
.B1(n_106),
.B2(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_27),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_120),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_30),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_51),
.B(n_30),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_126),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_32),
.B1(n_39),
.B2(n_4),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_106),
.B(n_112),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_62),
.B(n_32),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_48),
.A2(n_5),
.B1(n_39),
.B2(n_53),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_76),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_153),
.Y(n_182)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_131),
.Y(n_169)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_146),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_87),
.B(n_5),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_77),
.B1(n_79),
.B2(n_44),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_160),
.B1(n_164),
.B2(n_85),
.Y(n_171)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_88),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_150),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_97),
.A2(n_5),
.B1(n_118),
.B2(n_91),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_110),
.A2(n_97),
.B(n_89),
.C(n_129),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_92),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_113),
.Y(n_180)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_162),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_91),
.B1(n_86),
.B2(n_122),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_98),
.B(n_90),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_155),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_122),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_124),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_108),
.B(n_119),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_165),
.B(n_162),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_101),
.C(n_113),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_85),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_131),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_168),
.B(n_188),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_101),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_157),
.B(n_149),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_133),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_192),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_135),
.B(n_140),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_151),
.Y(n_202)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_145),
.B(n_161),
.C(n_130),
.D(n_153),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_196),
.A2(n_167),
.B(n_185),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_182),
.A2(n_145),
.B1(n_158),
.B2(n_142),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_199),
.B1(n_204),
.B2(n_198),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_170),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_147),
.B1(n_154),
.B2(n_139),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_200),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_202),
.B(n_203),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_143),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_132),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_141),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_187),
.B(n_180),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_162),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_134),
.Y(n_208)
);

NOR2x1_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_167),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_212),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_168),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_211),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_173),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_187),
.B(n_169),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_197),
.B(n_210),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_209),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_223),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_174),
.Y(n_223)
);

NOR4xp25_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_170),
.C(n_185),
.D(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_174),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_227),
.Y(n_234)
);

AO221x1_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_199),
.B1(n_213),
.B2(n_205),
.C(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_236),
.B1(n_237),
.B2(n_240),
.Y(n_241)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_194),
.B(n_207),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_194),
.B(n_201),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_221),
.C(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_237),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_SL g244 ( 
.A(n_230),
.B(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_249),
.C(n_238),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_233),
.A2(n_228),
.B1(n_216),
.B2(n_222),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_246),
.B1(n_236),
.B2(n_229),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_218),
.B1(n_219),
.B2(n_208),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_213),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_247),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_255),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_241),
.B(n_244),
.Y(n_259)
);

AOI31xp33_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_254),
.A3(n_243),
.B(n_242),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_256),
.B(n_175),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_183),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_183),
.C(n_175),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_251),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_191),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_259),
.A2(n_261),
.B(n_184),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

AOI21x1_ASAP7_75t_L g262 ( 
.A1(n_257),
.A2(n_255),
.B(n_176),
.Y(n_262)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_262),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_265),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_186),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_191),
.C(n_186),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_269),
.A2(n_270),
.B(n_176),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_176),
.Y(n_272)
);


endmodule