module real_jpeg_21385_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_0),
.A2(n_65),
.B1(n_66),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_0),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_0),
.A2(n_41),
.B1(n_48),
.B2(n_92),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_92),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_92),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_1),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_1),
.B(n_71),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_1),
.A2(n_16),
.B(n_33),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_132),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_188),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_1),
.B(n_87),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g218 ( 
.A1(n_1),
.A2(n_48),
.B(n_219),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_2),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_41),
.B1(n_48),
.B2(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_67),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_47),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_4),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_4),
.A2(n_41),
.B1(n_48),
.B2(n_134),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_134),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_134),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_5),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_5),
.A2(n_41),
.B1(n_48),
.B2(n_114),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_114),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_114),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_6),
.A2(n_41),
.B1(n_48),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_50),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_50),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_79)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_13),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_13),
.A2(n_41),
.B1(n_48),
.B2(n_74),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_74),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_74),
.Y(n_163)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_14),
.A2(n_30),
.A3(n_48),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_16),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_95),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_22),
.B(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_76),
.B2(n_94),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_52),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_39),
.B(n_51),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_26),
.B(n_39),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_27),
.A2(n_32),
.B1(n_35),
.B2(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_27),
.A2(n_32),
.B1(n_59),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_27),
.A2(n_32),
.B1(n_82),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_27),
.A2(n_32),
.B1(n_107),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_27),
.A2(n_32),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_27),
.A2(n_32),
.B1(n_184),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_27),
.A2(n_32),
.B1(n_204),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_27),
.A2(n_32),
.B1(n_125),
.B2(n_222),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_29),
.B(n_42),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_30),
.A2(n_31),
.B(n_132),
.C(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_32),
.B(n_132),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_34),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_39)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_40),
.A2(n_44),
.B1(n_85),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_40),
.A2(n_44),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_40),
.A2(n_44),
.B1(n_110),
.B2(n_129),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_40),
.A2(n_44),
.B1(n_158),
.B2(n_218),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_42),
.Y(n_43)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_48),
.B1(n_69),
.B2(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_41),
.A2(n_70),
.B1(n_131),
.B2(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_41),
.B(n_132),
.Y(n_215)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_48),
.B(n_69),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_60),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_61),
.B1(n_62),
.B2(n_75),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_58),
.B1(n_75),
.B2(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B(n_57),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_57),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_55),
.A2(n_56),
.B1(n_79),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_55),
.A2(n_105),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_55),
.A2(n_56),
.B1(n_146),
.B2(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_55),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_55),
.A2(n_147),
.B1(n_174),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_55),
.A2(n_56),
.B1(n_176),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_55),
.A2(n_56),
.B1(n_163),
.B2(n_206),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_56),
.B(n_132),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_58),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_69),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g131 ( 
.A(n_66),
.B(n_132),
.CON(n_131),
.SN(n_131)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_68),
.A2(n_71),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_76),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.C(n_88),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_78),
.B(n_81),
.Y(n_254)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_88),
.B1(n_89),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_86),
.A2(n_87),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_90),
.A2(n_93),
.B1(n_113),
.B2(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_102),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_100),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_102),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_111),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_103),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_260),
.B(n_265),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_164),
.B(n_247),
.C(n_259),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_149),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_119),
.B(n_149),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_135),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_121),
.B(n_122),
.C(n_135),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_130),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_133),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_137),
.B(n_141),
.C(n_142),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_140),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_172),
.B1(n_173),
.B2(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_154),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_150),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_161),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_156),
.B(n_232),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_160),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_246),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_241),
.B(n_245),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_227),
.B(n_240),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_208),
.B(n_226),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_196),
.B(n_207),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_185),
.B(n_195),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_177),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_181),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_190),
.B(n_194),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_189),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_198),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_210),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_216),
.B1(n_224),
.B2(n_225),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_211),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_220),
.B1(n_221),
.B2(n_223),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_223),
.C(n_224),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_229),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_237),
.C(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_236),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_237),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_249),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_258),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_256),
.C(n_258),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);


endmodule