module fake_jpeg_11733_n_440 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_5),
.B(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_48),
.B(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_50),
.Y(n_133)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_53),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_15),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_54),
.B(n_92),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_58),
.B(n_68),
.Y(n_129)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_14),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_73),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_24),
.B(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_85),
.Y(n_112)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_12),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_91),
.Y(n_110)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_12),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_24),
.B1(n_28),
.B2(n_18),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_101),
.A2(n_141),
.B1(n_28),
.B2(n_36),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_21),
.B1(n_44),
.B2(n_41),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_102),
.A2(n_22),
.B1(n_55),
.B2(n_50),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_54),
.A2(n_29),
.B1(n_37),
.B2(n_41),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_103),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_37),
.B(n_17),
.C(n_18),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_119),
.B(n_120),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_65),
.B(n_27),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_53),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_140),
.Y(n_162)
);

HAxp5_ASAP7_75t_SL g124 ( 
.A(n_66),
.B(n_31),
.CON(n_124),
.SN(n_124)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_25),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_26),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_135),
.B(n_139),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_60),
.A2(n_18),
.B(n_17),
.C(n_36),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_19),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_56),
.A2(n_17),
.B1(n_28),
.B2(n_36),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_86),
.B(n_44),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_26),
.Y(n_171)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_145),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_62),
.B1(n_76),
.B2(n_72),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_146),
.A2(n_178),
.B1(n_189),
.B2(n_7),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_83),
.B1(n_79),
.B2(n_47),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_147),
.A2(n_179),
.B1(n_182),
.B2(n_131),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_148),
.Y(n_228)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_149),
.Y(n_227)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_78),
.C(n_67),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_152),
.B(n_191),
.C(n_131),
.Y(n_213)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_157),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_158),
.B(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_60),
.B1(n_34),
.B2(n_21),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_109),
.Y(n_163)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_34),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_166),
.B(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_110),
.B(n_31),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_180),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_176),
.Y(n_198)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_108),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_22),
.B1(n_25),
.B2(n_126),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_96),
.A2(n_90),
.B1(n_88),
.B2(n_45),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_113),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_181),
.A2(n_186),
.B1(n_194),
.B2(n_115),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_101),
.A2(n_45),
.B1(n_1),
.B2(n_2),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_119),
.B(n_0),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_190),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_184),
.B(n_188),
.Y(n_197)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_187),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_99),
.A2(n_45),
.B1(n_4),
.B2(n_5),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_94),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_6),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_141),
.B(n_118),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_132),
.B(n_6),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_193),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_144),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_195),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_115),
.B1(n_144),
.B2(n_117),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_196),
.A2(n_200),
.B1(n_209),
.B2(n_216),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_190),
.A2(n_117),
.B1(n_136),
.B2(n_127),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_169),
.B(n_136),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_220),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_127),
.B1(n_105),
.B2(n_137),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_105),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_230),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_213),
.B(n_222),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_152),
.B(n_106),
.C(n_133),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_133),
.B1(n_137),
.B2(n_10),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_7),
.C(n_9),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_160),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_148),
.B1(n_157),
.B2(n_194),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_173),
.A2(n_162),
.B(n_163),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_205),
.B(n_198),
.Y(n_245)
);

O2A1O1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_226)
);

OA21x2_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_198),
.B(n_207),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_168),
.B(n_153),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_154),
.A2(n_145),
.B(n_178),
.C(n_159),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_207),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g234 ( 
.A1(n_147),
.A2(n_187),
.A3(n_188),
.B1(n_180),
.B2(n_156),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_193),
.Y(n_250)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_241),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_211),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_243),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_203),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_206),
.A2(n_189),
.B1(n_150),
.B2(n_165),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_244),
.A2(n_258),
.B1(n_260),
.B2(n_277),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_245),
.B(n_247),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_204),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_246),
.B(n_249),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_248),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_198),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_251),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_212),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_219),
.B(n_174),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_254),
.B(n_256),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_265),
.B1(n_272),
.B2(n_217),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_197),
.B(n_185),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_206),
.A2(n_176),
.B1(n_149),
.B2(n_175),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_259),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_216),
.A2(n_155),
.B1(n_164),
.B2(n_205),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_262),
.A2(n_264),
.B(n_267),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_221),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_273),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_210),
.A2(n_213),
.B1(n_237),
.B2(n_222),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_237),
.A2(n_208),
.B(n_231),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_265),
.B(n_261),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_SL g267 ( 
.A(n_225),
.B(n_226),
.C(n_222),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_222),
.A2(n_220),
.B1(n_234),
.B2(n_227),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_268),
.A2(n_264),
.B(n_239),
.Y(n_295)
);

AOI22x1_ASAP7_75t_L g270 ( 
.A1(n_238),
.A2(n_236),
.B1(n_199),
.B2(n_232),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_255),
.B(n_271),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_229),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_275),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_227),
.B1(n_202),
.B2(n_217),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_201),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_274),
.B(n_277),
.Y(n_299)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_257),
.Y(n_298)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_233),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_270),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_278),
.B(n_283),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_262),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_279),
.B(n_302),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_310),
.B1(n_276),
.B2(n_248),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_218),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_305),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_223),
.B(n_202),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_287),
.A2(n_303),
.B(n_283),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_218),
.B1(n_253),
.B2(n_260),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_288),
.A2(n_290),
.B(n_295),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_261),
.C(n_240),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_289),
.B(n_300),
.C(n_290),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_244),
.A2(n_258),
.B1(n_263),
.B2(n_269),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_291),
.A2(n_278),
.B1(n_294),
.B2(n_286),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_272),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_297),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_239),
.Y(n_297)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_252),
.B(n_245),
.C(n_247),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_275),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_268),
.A2(n_251),
.B(n_247),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_242),
.B(n_241),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_308),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_264),
.Y(n_308)
);

AO22x1_ASAP7_75t_SL g312 ( 
.A1(n_279),
.A2(n_270),
.B1(n_267),
.B2(n_273),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_327),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_313),
.A2(n_335),
.B1(n_288),
.B2(n_291),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_300),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_322),
.C(n_333),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_319),
.Y(n_363)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_320),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_296),
.Y(n_358)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_300),
.B(n_289),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_325),
.B(n_296),
.Y(n_360)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_309),
.Y(n_326)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_304),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_329),
.Y(n_356)
);

HB1xp67_ASAP7_75t_SL g331 ( 
.A(n_285),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_331),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_284),
.B(n_281),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_332),
.B(n_337),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_283),
.C(n_287),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_286),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_336),
.Y(n_351)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_284),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_302),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_285),
.A2(n_281),
.B(n_308),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_339),
.A2(n_292),
.B(n_307),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_292),
.C(n_307),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_299),
.C(n_301),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_342),
.A2(n_323),
.B(n_318),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_330),
.A2(n_282),
.B1(n_310),
.B2(n_288),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_345),
.A2(n_359),
.B1(n_313),
.B2(n_318),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_346),
.A2(n_363),
.B1(n_344),
.B2(n_349),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_358),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_317),
.B(n_299),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_352),
.C(n_354),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_322),
.C(n_333),
.Y(n_352)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_353),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_340),
.B(n_296),
.C(n_305),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_330),
.A2(n_310),
.B1(n_306),
.B2(n_311),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_343),
.C(n_352),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_334),
.B(n_306),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_316),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_328),
.Y(n_364)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_339),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_370),
.C(n_375),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_367),
.A2(n_377),
.B(n_341),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_353),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_368),
.B(n_379),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_327),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_346),
.A2(n_330),
.B1(n_320),
.B2(n_324),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_372),
.A2(n_376),
.B1(n_359),
.B2(n_345),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_372),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_374),
.B(n_378),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_314),
.C(n_315),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_341),
.A2(n_314),
.B(n_315),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_316),
.C(n_312),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_312),
.C(n_338),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_381),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_347),
.B(n_336),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_382),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_326),
.Y(n_384)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_384),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_387),
.A2(n_373),
.B1(n_382),
.B2(n_351),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_379),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_388),
.B(n_392),
.C(n_396),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_354),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_393),
.Y(n_401)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_394),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_358),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_397),
.A2(n_356),
.B1(n_355),
.B2(n_357),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_367),
.A2(n_362),
.B(n_380),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_398),
.B(n_378),
.Y(n_407)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_376),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_357),
.Y(n_410)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_402),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_385),
.A2(n_377),
.B1(n_371),
.B2(n_310),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_408),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_410),
.Y(n_414)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_386),
.Y(n_409)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_409),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_400),
.A2(n_374),
.B(n_329),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_411),
.B(n_412),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_395),
.B(n_298),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_390),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_421),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_396),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_416),
.B(n_417),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_398),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_406),
.B(n_391),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_388),
.C(n_392),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_422),
.B(n_389),
.C(n_410),
.Y(n_427)
);

XOR2x2_ASAP7_75t_L g424 ( 
.A(n_417),
.B(n_405),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_424),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_422),
.B(n_389),
.C(n_397),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_427),
.C(n_416),
.Y(n_430)
);

AOI21xp33_ASAP7_75t_L g426 ( 
.A1(n_419),
.A2(n_405),
.B(n_399),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_426),
.A2(n_415),
.B(n_403),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_401),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_420),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_430),
.A2(n_432),
.B(n_433),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_431),
.A2(n_429),
.B(n_425),
.Y(n_435)
);

AOI321xp33_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_418),
.A3(n_424),
.B1(n_431),
.B2(n_423),
.C(n_408),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_436),
.A2(n_418),
.B1(n_434),
.B2(n_321),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_296),
.C(n_280),
.Y(n_438)
);

NOR2x1_ASAP7_75t_SL g439 ( 
.A(n_438),
.B(n_280),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_280),
.Y(n_440)
);


endmodule