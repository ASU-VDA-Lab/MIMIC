module fake_jpeg_19724_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_40),
.B(n_10),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_16),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_20),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_53),
.B(n_55),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_34),
.B1(n_20),
.B2(n_33),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_54),
.A2(n_98),
.B1(n_28),
.B2(n_8),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_65),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_61),
.A2(n_69),
.B1(n_76),
.B2(n_85),
.Y(n_115)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_71),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_19),
.C(n_31),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_19),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_18),
.B1(n_36),
.B2(n_24),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_17),
.B1(n_36),
.B2(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_36),
.B1(n_35),
.B2(n_25),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_17),
.B1(n_38),
.B2(n_24),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_26),
.B1(n_38),
.B2(n_33),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_46),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_27),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_83),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_27),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_29),
.B1(n_35),
.B2(n_25),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_35),
.B1(n_25),
.B2(n_28),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_88),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_40),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_31),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_92),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_46),
.B(n_31),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_32),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_46),
.A2(n_34),
.B1(n_32),
.B2(n_37),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_9),
.B1(n_11),
.B2(n_10),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_31),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_100),
.Y(n_131)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_9),
.B1(n_12),
.B2(n_11),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_46),
.A2(n_19),
.B(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_R g111 ( 
.A(n_99),
.B(n_0),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_46),
.B(n_19),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_91),
.B(n_74),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_113),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_66),
.A2(n_32),
.B1(n_28),
.B2(n_19),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_32),
.B1(n_28),
.B2(n_37),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_37),
.Y(n_109)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_111),
.B(n_112),
.CI(n_130),
.CON(n_157),
.SN(n_157)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_64),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_122),
.B1(n_127),
.B2(n_129),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_121),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_54),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_128),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_59),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_98),
.A2(n_8),
.B1(n_12),
.B2(n_7),
.Y(n_129)
);

BUFx24_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

NAND2x1_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_65),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_136),
.A2(n_150),
.B(n_134),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_106),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_140),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_55),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_153),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_83),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_67),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_101),
.C(n_116),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_93),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_145),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_109),
.B(n_53),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_53),
.B1(n_75),
.B2(n_73),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_148),
.A2(n_114),
.B1(n_58),
.B2(n_70),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_117),
.B(n_56),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_88),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_154),
.B(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_92),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_97),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_62),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_163),
.Y(n_199)
);

AO21x2_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_84),
.B(n_60),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_72),
.B1(n_58),
.B2(n_116),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_108),
.B(n_57),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_62),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_164),
.B(n_165),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_125),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_167),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_127),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_118),
.B(n_70),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_197),
.B1(n_162),
.B2(n_155),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_176),
.B(n_191),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_183),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_105),
.B1(n_101),
.B2(n_104),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_178),
.A2(n_179),
.B1(n_184),
.B2(n_143),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_144),
.B1(n_163),
.B2(n_145),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_181),
.A2(n_157),
.B1(n_165),
.B2(n_149),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_164),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_101),
.B1(n_111),
.B2(n_57),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_193),
.C(n_137),
.Y(n_208)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_190),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_128),
.B(n_120),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_195),
.B(n_201),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_147),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_110),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_116),
.C(n_59),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_122),
.C(n_113),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_196),
.B(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_151),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_198),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_110),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_136),
.A2(n_107),
.B(n_132),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_140),
.B(n_81),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_168),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_178),
.A2(n_148),
.B1(n_162),
.B2(n_142),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_204),
.A2(n_206),
.B1(n_210),
.B2(n_228),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_229),
.B1(n_199),
.B2(n_192),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_194),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_209),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_146),
.B1(n_138),
.B2(n_137),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_216),
.B(n_227),
.Y(n_232)
);

HB1xp67_ASAP7_75t_SL g213 ( 
.A(n_201),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_203),
.B(n_175),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_174),
.B(n_175),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_219),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_162),
.B(n_156),
.Y(n_216)
);

AOI221xp5_ASAP7_75t_L g217 ( 
.A1(n_182),
.A2(n_157),
.B1(n_139),
.B2(n_158),
.C(n_153),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_157),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_166),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_221),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_174),
.B(n_146),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_59),
.C(n_162),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_193),
.C(n_188),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_162),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_225),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_152),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_176),
.A2(n_172),
.B(n_170),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_184),
.A2(n_72),
.B1(n_60),
.B2(n_63),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_107),
.B1(n_132),
.B2(n_12),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_173),
.B(n_59),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_230),
.Y(n_241)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_243),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_244),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_222),
.C(n_206),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_238),
.C(n_249),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_247),
.B(n_212),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_202),
.C(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_240),
.Y(n_273)
);

XOR2x2_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_218),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_192),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_204),
.B1(n_228),
.B2(n_223),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_203),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_202),
.C(n_196),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_202),
.C(n_190),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_254),
.C(n_209),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_187),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_211),
.Y(n_259)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_218),
.B(n_195),
.CI(n_177),
.CON(n_253),
.SN(n_253)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_227),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_261),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_258),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_247),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_216),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_242),
.A3(n_232),
.B1(n_248),
.B2(n_252),
.C1(n_215),
.C2(n_237),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_235),
.Y(n_276)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_243),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_267),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_238),
.C(n_249),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_232),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_220),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_270),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_246),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_271),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_225),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_280),
.C(n_287),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_276),
.B(n_283),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_250),
.C(n_244),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_253),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_253),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_288),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_273),
.Y(n_286)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_246),
.C(n_231),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_214),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_289),
.A2(n_189),
.B1(n_226),
.B2(n_207),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_268),
.C(n_266),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_294),
.C(n_302),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_260),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_299),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_272),
.B(n_273),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_277),
.B(n_211),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_260),
.C(n_270),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_282),
.B(n_226),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_278),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_301),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_255),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_284),
.A2(n_257),
.B1(n_205),
.B2(n_264),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_217),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_305),
.Y(n_314)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_307),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_275),
.C(n_274),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_231),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_299),
.A2(n_286),
.B(n_241),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_241),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_318),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_312),
.A2(n_295),
.B(n_290),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_319),
.B(n_230),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_294),
.C(n_291),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_292),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_230),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_310),
.C(n_319),
.Y(n_324)
);

NAND2xp33_ASAP7_75t_SL g321 ( 
.A(n_314),
.B(n_230),
.Y(n_321)
);

O2A1O1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_321),
.A2(n_316),
.B(n_207),
.C(n_194),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_307),
.B1(n_311),
.B2(n_229),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_325),
.B(n_198),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_313),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_327),
.C(n_328),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_322),
.C(n_324),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_323),
.Y(n_331)
);


endmodule