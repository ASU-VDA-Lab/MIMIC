module real_jpeg_32914_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g175 ( 
.A(n_0),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_0),
.Y(n_179)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_0),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_0),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_507),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_1),
.B(n_508),
.Y(n_507)
);

AO22x1_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_2),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_109),
.B1(n_117),
.B2(n_120),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_2),
.A2(n_109),
.B1(n_163),
.B2(n_167),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_2),
.A2(n_109),
.B1(n_290),
.B2(n_292),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_3),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_5),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_6),
.A2(n_62),
.B1(n_66),
.B2(n_72),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_6),
.A2(n_72),
.B1(n_191),
.B2(n_196),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_6),
.A2(n_72),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_6),
.A2(n_72),
.B1(n_283),
.B2(n_285),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_7),
.Y(n_508)
);

OAI22x1_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

AO22x1_ASAP7_75t_L g184 ( 
.A1(n_8),
.A2(n_56),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

AOI22x1_ASAP7_75t_SL g214 ( 
.A1(n_8),
.A2(n_56),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_8),
.B(n_369),
.Y(n_368)
);

OAI32xp33_ASAP7_75t_L g390 ( 
.A1(n_8),
.A2(n_391),
.A3(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_8),
.B(n_155),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_11),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_11),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_11),
.A2(n_246),
.B1(n_255),
.B2(n_258),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g350 ( 
.A1(n_11),
.A2(n_246),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_L g411 ( 
.A1(n_11),
.A2(n_246),
.B1(n_412),
.B2(n_414),
.Y(n_411)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_233),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_231),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_202),
.Y(n_17)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_18),
.B(n_202),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_151),
.C(n_170),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_20),
.B(n_151),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_113),
.B2(n_114),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_23),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g209 ( 
.A1(n_23),
.A2(n_206),
.B1(n_210),
.B2(n_220),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_23),
.A2(n_206),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_23),
.B(n_241),
.C(n_252),
.Y(n_309)
);

OA21x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_50),
.B(n_51),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_24),
.B(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_24),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_24),
.B(n_51),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_24),
.B(n_350),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_33),
.B2(n_35),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_32),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_32),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_R g431 ( 
.A(n_39),
.B(n_56),
.Y(n_431)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_46),
.B2(n_49),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_42),
.Y(n_405)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_45),
.Y(n_287)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_50),
.Y(n_160)
);

NAND2x1p5_ASAP7_75t_L g199 ( 
.A(n_50),
.B(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_50),
.B(n_190),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_50),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_51),
.B(n_160),
.Y(n_159)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_55),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_55),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_56),
.A2(n_136),
.B(n_138),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_56),
.B(n_139),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_SL g298 ( 
.A(n_56),
.B(n_126),
.Y(n_298)
);

AOI32xp33_ASAP7_75t_L g362 ( 
.A1(n_56),
.A2(n_363),
.A3(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_56),
.B(n_392),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_56),
.B(n_178),
.Y(n_440)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_59),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_59),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g205 ( 
.A(n_60),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_73),
.B(n_101),
.Y(n_60)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_65),
.Y(n_216)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_71),
.Y(n_274)
);

INVxp33_ASAP7_75t_SL g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2x1_ASAP7_75t_L g157 ( 
.A(n_74),
.B(n_105),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_74),
.B(n_254),
.Y(n_297)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_75),
.A2(n_214),
.B(n_329),
.Y(n_328)
);

NOR2x1_ASAP7_75t_L g359 ( 
.A(n_75),
.B(n_214),
.Y(n_359)
);

AO21x2_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_83),
.B(n_92),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_77),
.Y(n_366)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_83),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_99),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_98),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_101),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_102),
.B(n_359),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_103),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_104),
.Y(n_329)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_108),
.Y(n_263)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_112),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_113),
.A2(n_114),
.B1(n_204),
.B2(n_207),
.Y(n_203)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_114),
.B(n_205),
.C(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_134),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_115),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_125),
.Y(n_115)
);

NAND2x1p5_ASAP7_75t_L g230 ( 
.A(n_116),
.B(n_141),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_118),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_119),
.Y(n_228)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_121),
.Y(n_224)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_123),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_125),
.B(n_135),
.Y(n_477)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OA21x2_ASAP7_75t_SL g221 ( 
.A1(n_126),
.A2(n_222),
.B(n_229),
.Y(n_221)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2x1p5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_127),
.A2(n_135),
.B(n_141),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_127),
.B(n_243),
.Y(n_242)
);

AO22x2_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_133),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_134),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_138),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_141),
.B(n_243),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_148),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_150),
.Y(n_266)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_152),
.A2(n_153),
.B(n_158),
.Y(n_489)
);

NAND2x1_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

AOI21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_155),
.B(n_254),
.Y(n_253)
);

NOR2x1_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2x1p5_ASAP7_75t_L g252 ( 
.A(n_157),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_159),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_161),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_161),
.B(n_349),
.Y(n_348)
);

AO21x1_ASAP7_75t_L g474 ( 
.A1(n_161),
.A2(n_334),
.B(n_335),
.Y(n_474)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_170),
.B(n_504),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_173),
.B(n_200),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_171),
.B(n_491),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_188),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_172),
.A2(n_173),
.B1(n_362),
.B2(n_373),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_172),
.A2(n_173),
.B1(n_188),
.B2(n_472),
.Y(n_471)
);

OAI22xp33_ASAP7_75t_L g491 ( 
.A1(n_172),
.A2(n_173),
.B1(n_201),
.B2(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_SL g384 ( 
.A(n_173),
.B(n_362),
.Y(n_384)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_176),
.B(n_183),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_176),
.A2(n_282),
.B(n_303),
.Y(n_311)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_177),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_177),
.B(n_184),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_177),
.B(n_411),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_179),
.Y(n_305)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_181),
.Y(n_284)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_181),
.Y(n_414)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_182),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_182),
.Y(n_413)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_182),
.Y(n_439)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_184),
.B(n_337),
.Y(n_336)
);

BUFx4f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_188),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_198),
.B(n_199),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_199),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_199),
.B(n_383),
.Y(n_417)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_201),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_221),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_212),
.B(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2x1p5_ASAP7_75t_L g327 ( 
.A(n_230),
.B(n_242),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_499),
.B(n_505),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_458),
.B(n_496),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_343),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_320),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_306),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_239),
.B(n_307),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_259),
.C(n_294),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_240),
.B(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_250),
.Y(n_240)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_244),
.Y(n_267)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_253),
.B(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XOR2x2_ASAP7_75t_L g454 ( 
.A(n_259),
.B(n_295),
.Y(n_454)
);

XNOR2x1_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_276),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_260),
.B(n_276),
.Y(n_315)
);

OAI31xp33_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_264),
.A3(n_267),
.B(n_268),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_272),
.B(n_275),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_282),
.B(n_288),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_288),
.B(n_336),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_288),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_304),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.C(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_296),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_378),
.Y(n_380)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_301),
.Y(n_435)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_303),
.B(n_410),
.Y(n_432)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_314),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_314),
.C(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_310),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_312),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_313),
.B(n_349),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_317),
.C(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

NAND2x1_ASAP7_75t_L g476 ( 
.A(n_318),
.B(n_477),
.Y(n_476)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_341),
.Y(n_320)
);

AO21x1_ASAP7_75t_L g459 ( 
.A1(n_321),
.A2(n_341),
.B(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_321),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_322),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_331),
.B1(n_332),
.B2(n_340),
.Y(n_324)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_325),
.Y(n_464)
);

XOR2x1_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

XOR2x1_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_327),
.B(n_330),
.C(n_468),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_328),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_331),
.B(n_463),
.C(n_465),
.Y(n_462)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2x1_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

AND2x4_ASAP7_75t_SL g409 ( 
.A(n_336),
.B(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_341),
.Y(n_479)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_452),
.B(n_456),
.Y(n_343)
);

OAI21x1_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_385),
.B(n_451),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_374),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_346),
.B(n_374),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_357),
.C(n_360),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2x1_ASAP7_75t_L g449 ( 
.A(n_348),
.B(n_357),
.Y(n_449)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_SL g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_361),
.B(n_449),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_362),
.Y(n_373)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_381),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_375),
.B(n_382),
.C(n_384),
.Y(n_455)
);

OAI22x1_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_379),
.B2(n_380),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_376),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_444),
.B(n_450),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_420),
.B(n_443),
.Y(n_386)
);

NOR2x1_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_408),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_388),
.B(n_408),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_406),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_389),
.A2(n_390),
.B1(n_406),
.B2(n_407),
.Y(n_422)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_398),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_415),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_409),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_415)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_416),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_417),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_417),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_446),
.C(n_447),
.Y(n_445)
);

AOI21x1_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_429),
.B(n_442),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NOR2x1_ASAP7_75t_L g442 ( 
.A(n_422),
.B(n_423),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_435),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

OAI21x1_ASAP7_75t_SL g429 ( 
.A1(n_430),
.A2(n_433),
.B(n_441),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_432),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_432),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_440),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_448),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_445),
.B(n_448),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_453),
.B(n_455),
.Y(n_457)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NAND3xp33_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_461),
.C(n_481),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_466),
.B1(n_479),
.B2(n_480),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_462),
.B(n_466),
.Y(n_498)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_469),
.Y(n_466)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_473),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_471),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g486 ( 
.A(n_473),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

MAJx2_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_494),
.C(n_495),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.Y(n_475)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_478),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_481),
.A2(n_497),
.B(n_498),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_487),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_487),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.C(n_485),
.Y(n_482)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_493),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

INVxp33_ASAP7_75t_L g501 ( 
.A(n_489),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_490),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_501),
.C(n_502),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_503),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_500),
.B(n_503),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);


endmodule