module fake_jpeg_9927_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_43),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_22),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_22),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_50),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_28),
.B(n_18),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_53),
.Y(n_72)
);

CKINVDCx9p33_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_39),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_65),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_22),
.B1(n_20),
.B2(n_25),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_24),
.B1(n_34),
.B2(n_17),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_20),
.B1(n_25),
.B2(n_29),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_71),
.B1(n_25),
.B2(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_21),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_20),
.B1(n_25),
.B2(n_23),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_68),
.B1(n_55),
.B2(n_51),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_75),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_28),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_84),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_48),
.B(n_24),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_70),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_26),
.B1(n_34),
.B2(n_17),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_85),
.B(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_87),
.Y(n_120)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_57),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_95),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_34),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_98),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_50),
.A3(n_55),
.B1(n_49),
.B2(n_69),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_92),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_90),
.B1(n_89),
.B2(n_74),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_76),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_68),
.B1(n_58),
.B2(n_71),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_110),
.B1(n_113),
.B2(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_106),
.B(n_118),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_67),
.C(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_122),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_68),
.B1(n_49),
.B2(n_58),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_108),
.A2(n_116),
.B1(n_121),
.B2(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_82),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_55),
.B1(n_88),
.B2(n_87),
.Y(n_110)
);

NAND2x1p5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_62),
.Y(n_112)
);

OR2x4_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_82),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_47),
.B1(n_54),
.B2(n_59),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_85),
.A2(n_47),
.B1(n_54),
.B2(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_54),
.B1(n_59),
.B2(n_19),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_18),
.B(n_27),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_74),
.C(n_27),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_125),
.B(n_126),
.Y(n_177)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_73),
.B1(n_83),
.B2(n_88),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_135),
.B1(n_138),
.B2(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_134),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_79),
.B1(n_76),
.B2(n_94),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_146),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_91),
.B1(n_54),
.B2(n_59),
.Y(n_138)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_140),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_145),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_57),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_150),
.Y(n_154)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_57),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_57),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_149),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_56),
.B1(n_26),
.B2(n_19),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_98),
.B(n_32),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_152),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_102),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_161),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_127),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_129),
.B1(n_151),
.B2(n_128),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_165),
.B1(n_171),
.B2(n_179),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_102),
.B(n_107),
.C(n_123),
.D(n_108),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_169),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_97),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_121),
.B1(n_113),
.B2(n_106),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_119),
.B1(n_115),
.B2(n_56),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_173),
.B(n_126),
.Y(n_188)
);

CKINVDCx12_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_130),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_178),
.B(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_115),
.B1(n_111),
.B2(n_101),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_140),
.B(n_12),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_12),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_188),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_132),
.B1(n_142),
.B2(n_131),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_187),
.A2(n_205),
.B1(n_208),
.B2(n_200),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_176),
.A2(n_135),
.B1(n_137),
.B2(n_133),
.Y(n_189)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_193),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_155),
.A2(n_153),
.B1(n_160),
.B2(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_195),
.B1(n_200),
.B2(n_206),
.Y(n_214)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_182),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_196),
.A2(n_197),
.B(n_204),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_149),
.B(n_93),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_134),
.B1(n_101),
.B2(n_100),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_156),
.B1(n_208),
.B2(n_203),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_158),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_100),
.B1(n_96),
.B2(n_93),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_96),
.B1(n_26),
.B2(n_27),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_170),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_212),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_228),
.B1(n_217),
.B2(n_196),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_170),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_167),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_226),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_167),
.C(n_177),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_218),
.C(n_223),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_177),
.C(n_168),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_225),
.B1(n_221),
.B2(n_217),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_232),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_168),
.C(n_166),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_166),
.C(n_173),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_227),
.C(n_199),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_178),
.B(n_164),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_173),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_161),
.C(n_163),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_185),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_229)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_229),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_186),
.A2(n_16),
.B1(n_8),
.B2(n_10),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_231),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_222),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_185),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_193),
.Y(n_239)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_218),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_249),
.C(n_212),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_190),
.B1(n_206),
.B2(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_216),
.A2(n_186),
.B1(n_230),
.B2(n_194),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_248),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_204),
.B1(n_202),
.B2(n_183),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_202),
.C(n_2),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_231),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_235),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_11),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_244),
.A2(n_221),
.B(n_211),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_256),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_226),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_209),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_250),
.C(n_246),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_239),
.B(n_223),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_264),
.B(n_11),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_238),
.B1(n_237),
.B2(n_236),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_224),
.B(n_228),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_16),
.B(n_13),
.Y(n_277)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_250),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_271),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_234),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_234),
.B1(n_241),
.B2(n_243),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_276),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_274),
.B(n_277),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_246),
.C(n_252),
.Y(n_276)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_12),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_0),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_257),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_281),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_265),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_289),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_275),
.A2(n_267),
.B1(n_261),
.B2(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_292),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_268),
.B1(n_266),
.B2(n_258),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_288),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_256),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_276),
.A2(n_258),
.B(n_4),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_284),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_296),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_271),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_273),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_3),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_270),
.C(n_4),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_300),
.C(n_3),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_291),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_303),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_293),
.A2(n_290),
.B(n_292),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_307)
);

AOI31xp67_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_3),
.A3(n_5),
.B(n_6),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_301),
.A2(n_299),
.B(n_294),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_302),
.B(n_6),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_309),
.B(n_307),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_5),
.B(n_6),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_5),
.Y(n_313)
);


endmodule