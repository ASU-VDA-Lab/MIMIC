module fake_ariane_3323_n_1104 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1104);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1104;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_885;
wire n_737;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_928;
wire n_839;
wire n_1099;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_1080;
wire n_576;
wire n_843;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_658;
wire n_617;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_741;
wire n_939;
wire n_747;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_1081;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_931;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1027;
wire n_615;
wire n_751;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_1025;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_68),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_105),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_148),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_5),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_106),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_88),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_90),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_155),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_164),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_111),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_100),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_97),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_204),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_146),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_65),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_83),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_124),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_172),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_32),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_64),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_205),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_192),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_200),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_12),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_8),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_154),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_47),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_66),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_109),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_33),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_119),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_134),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_72),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_147),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_196),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_191),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_21),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_149),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_181),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_12),
.Y(n_258)
);

BUFx2_ASAP7_75t_SL g259 ( 
.A(n_117),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_42),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_3),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_184),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_169),
.Y(n_263)
);

INVxp33_ASAP7_75t_R g264 ( 
.A(n_113),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_27),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_67),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_110),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_188),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_152),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_150),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_57),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_20),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_58),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_98),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_145),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_176),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_126),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_186),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_187),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_50),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_79),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_116),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_235),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_218),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_272),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_233),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_228),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_215),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_268),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_215),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_244),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_244),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_244),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_246),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_236),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_245),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_220),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_230),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_266),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_247),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_261),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_265),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_259),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_274),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_275),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_277),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_254),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_252),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_225),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_320),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_237),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_276),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_289),
.B(n_264),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_333),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_284),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_326),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_287),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_291),
.B(n_252),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_289),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_288),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_303),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_322),
.A2(n_283),
.B1(n_282),
.B2(n_281),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_285),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g354 ( 
.A1(n_326),
.A2(n_256),
.B(n_252),
.Y(n_354)
);

AOI22x1_ASAP7_75t_SL g355 ( 
.A1(n_287),
.A2(n_279),
.B1(n_278),
.B2(n_273),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_300),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_292),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_329),
.B(n_214),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_320),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_306),
.B(n_216),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_307),
.B(n_217),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

BUFx12f_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_308),
.B(n_219),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_310),
.B(n_221),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_295),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_285),
.A2(n_271),
.B1(n_270),
.B2(n_269),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_301),
.A2(n_267),
.B1(n_262),
.B2(n_257),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_330),
.B(n_252),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_300),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_294),
.A2(n_232),
.B1(n_253),
.B2(n_249),
.Y(n_375)
);

BUFx12f_ASAP7_75t_L g376 ( 
.A(n_313),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_321),
.A2(n_227),
.B1(n_239),
.B2(n_238),
.Y(n_377)
);

AO22x1_ASAP7_75t_L g378 ( 
.A1(n_302),
.A2(n_234),
.B1(n_229),
.B2(n_226),
.Y(n_378)
);

OAI22x1_ASAP7_75t_L g379 ( 
.A1(n_304),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_327),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_309),
.Y(n_382)
);

OAI21x1_ASAP7_75t_L g383 ( 
.A1(n_328),
.A2(n_256),
.B(n_36),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_311),
.B(n_256),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_293),
.A2(n_256),
.B(n_0),
.Y(n_385)
);

OAI22x1_ASAP7_75t_R g386 ( 
.A1(n_294),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_386)
);

AND2x2_ASAP7_75t_SL g387 ( 
.A(n_314),
.B(n_1),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_351),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_351),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_367),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_319),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_339),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_346),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_334),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_346),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_343),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_335),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_371),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_340),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_R g407 ( 
.A(n_382),
.B(n_290),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_340),
.B(n_331),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_355),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_372),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_377),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_375),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_338),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_342),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_348),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_348),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_334),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_345),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_360),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_380),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_360),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_378),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g428 ( 
.A(n_373),
.B(n_293),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_381),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_R g430 ( 
.A(n_363),
.B(n_312),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_349),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_364),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_364),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_379),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_368),
.B(n_331),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_R g437 ( 
.A(n_369),
.B(n_315),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_379),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_R g439 ( 
.A(n_337),
.B(n_316),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_336),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_373),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_387),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_386),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_387),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_384),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_362),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_339),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_362),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_350),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_352),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_376),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_353),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_R g455 ( 
.A(n_353),
.B(n_318),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_352),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_350),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_353),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_350),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_324),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_434),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_325),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_442),
.A2(n_445),
.B1(n_420),
.B2(n_405),
.Y(n_466)
);

CKINVDCx14_ASAP7_75t_R g467 ( 
.A(n_402),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_390),
.B(n_389),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_400),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_403),
.Y(n_470)
);

INVx5_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

AND2x6_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_296),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_419),
.B(n_296),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_399),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_418),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_406),
.B(n_297),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_428),
.A2(n_385),
.B1(n_297),
.B2(n_298),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_412),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_432),
.B(n_298),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_440),
.B(n_299),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_404),
.B(n_299),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_449),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_448),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_L g486 ( 
.A(n_433),
.B(n_350),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_399),
.B(n_385),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_410),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_417),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_441),
.B(n_332),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_427),
.B(n_356),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_394),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_401),
.B(n_421),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_R g494 ( 
.A(n_391),
.B(n_35),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_436),
.B(n_313),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_437),
.B(n_356),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_395),
.B(n_4),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_399),
.B(n_436),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_457),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_411),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_428),
.B(n_383),
.Y(n_504)
);

INVx8_ASAP7_75t_L g505 ( 
.A(n_428),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_428),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_408),
.Y(n_507)
);

INVx8_ASAP7_75t_L g508 ( 
.A(n_428),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_451),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_450),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_452),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_462),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_407),
.Y(n_515)
);

INVx8_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_415),
.B(n_5),
.Y(n_519)
);

INVx8_ASAP7_75t_L g520 ( 
.A(n_447),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_393),
.Y(n_521)
);

CKINVDCx11_ASAP7_75t_R g522 ( 
.A(n_444),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_437),
.B(n_356),
.Y(n_523)
);

BUFx4f_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_446),
.B(n_383),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_429),
.A2(n_323),
.B1(n_313),
.B2(n_354),
.Y(n_526)
);

AND2x2_ASAP7_75t_SL g527 ( 
.A(n_414),
.B(n_6),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_439),
.B(n_6),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_396),
.B(n_313),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_398),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_413),
.B(n_7),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_443),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_431),
.A2(n_323),
.B1(n_374),
.B2(n_358),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_430),
.B(n_323),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_454),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_458),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_456),
.Y(n_537)
);

NAND3x1_ASAP7_75t_L g538 ( 
.A(n_409),
.B(n_7),
.C(n_9),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_435),
.B(n_9),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_459),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_439),
.B(n_10),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_455),
.B(n_356),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_430),
.B(n_10),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_459),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_438),
.B(n_11),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_455),
.B(n_453),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_460),
.B(n_11),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_527),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_548)
);

AO22x2_ASAP7_75t_L g549 ( 
.A1(n_531),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_464),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_480),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_505),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_489),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_483),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_463),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_499),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_472),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_465),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_470),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_469),
.B(n_450),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_517),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_521),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_530),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_531),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_468),
.Y(n_565)
);

OR2x6_ASAP7_75t_L g566 ( 
.A(n_505),
.B(n_323),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_535),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_493),
.B(n_500),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_537),
.Y(n_569)
);

NAND2x1p5_ASAP7_75t_L g570 ( 
.A(n_471),
.B(n_358),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_475),
.B(n_16),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_471),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_536),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_471),
.B(n_358),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_476),
.B(n_17),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_493),
.B(n_388),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_476),
.B(n_18),
.Y(n_577)
);

NAND2x1p5_ASAP7_75t_L g578 ( 
.A(n_506),
.B(n_358),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_532),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_473),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_503),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_524),
.B(n_374),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_485),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_510),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_497),
.Y(n_585)
);

OAI221xp5_ASAP7_75t_L g586 ( 
.A1(n_488),
.A2(n_388),
.B1(n_374),
.B2(n_21),
.C(n_22),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_511),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_518),
.A2(n_323),
.B1(n_388),
.B2(n_374),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_528),
.A2(n_388),
.B1(n_20),
.B2(n_22),
.Y(n_589)
);

OR2x2_ASAP7_75t_SL g590 ( 
.A(n_519),
.B(n_19),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_467),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_482),
.B(n_19),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_501),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_500),
.B(n_23),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_509),
.Y(n_595)
);

NAND2x1p5_ASAP7_75t_L g596 ( 
.A(n_506),
.B(n_37),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_490),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_524),
.B(n_23),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_544),
.Y(n_600)
);

NAND2x1p5_ASAP7_75t_L g601 ( 
.A(n_476),
.B(n_38),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_492),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_478),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_522),
.Y(n_604)
);

AO22x2_ASAP7_75t_L g605 ( 
.A1(n_488),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_477),
.B(n_24),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_478),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_484),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_515),
.B(n_25),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_529),
.Y(n_610)
);

NAND2x1p5_ASAP7_75t_L g611 ( 
.A(n_512),
.B(n_40),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_529),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_507),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_555),
.B(n_500),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_576),
.A2(n_525),
.B(n_504),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_576),
.A2(n_525),
.B(n_546),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_568),
.A2(n_546),
.B(n_486),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_555),
.B(n_558),
.Y(n_618)
);

OAI21xp33_ASAP7_75t_L g619 ( 
.A1(n_558),
.A2(n_547),
.B(n_541),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_559),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_572),
.B(n_512),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_552),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_572),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_554),
.B(n_466),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_592),
.A2(n_520),
.B1(n_508),
.B2(n_505),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g626 ( 
.A1(n_568),
.A2(n_504),
.B(n_495),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_573),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_554),
.B(n_466),
.Y(n_628)
);

O2A1O1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_586),
.A2(n_481),
.B(n_543),
.C(n_539),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_560),
.B(n_514),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_582),
.A2(n_508),
.B(n_502),
.Y(n_631)
);

INVx11_ASAP7_75t_L g632 ( 
.A(n_604),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_565),
.B(n_513),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_602),
.B(n_513),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_591),
.B(n_586),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_597),
.B(n_565),
.Y(n_636)
);

INVx11_ASAP7_75t_L g637 ( 
.A(n_608),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_566),
.A2(n_508),
.B(n_520),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_571),
.B(n_500),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_613),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_551),
.A2(n_520),
.B1(n_514),
.B2(n_516),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_548),
.A2(n_516),
.B1(n_498),
.B2(n_534),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_603),
.B(n_512),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_L g644 ( 
.A(n_552),
.B(n_474),
.Y(n_644)
);

BUFx4f_ASAP7_75t_L g645 ( 
.A(n_607),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_566),
.A2(n_516),
.B(n_542),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_553),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_566),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_556),
.B(n_534),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_609),
.B(n_545),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_567),
.A2(n_523),
.B(n_496),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_549),
.A2(n_534),
.B1(n_538),
.B2(n_487),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_575),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_570),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_579),
.A2(n_474),
.B(n_479),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_561),
.B(n_562),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_575),
.Y(n_657)
);

OAI21xp33_ASAP7_75t_L g658 ( 
.A1(n_606),
.A2(n_494),
.B(n_491),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_563),
.B(n_533),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_550),
.B(n_533),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_570),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_569),
.A2(n_474),
.B(n_487),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_594),
.A2(n_578),
.B(n_599),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_578),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_594),
.A2(n_526),
.B(n_474),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_600),
.A2(n_487),
.B(n_122),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_549),
.A2(n_487),
.B1(n_27),
.B2(n_28),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_598),
.A2(n_123),
.B(n_212),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_581),
.B(n_26),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_584),
.B(n_28),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_612),
.B(n_29),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_595),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_587),
.B(n_29),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_577),
.B(n_30),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_577),
.B(n_30),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_616),
.A2(n_596),
.B(n_564),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_637),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_627),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_618),
.B(n_549),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_632),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_635),
.B(n_590),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_623),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_619),
.A2(n_589),
.B(n_605),
.C(n_611),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_640),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_624),
.B(n_611),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_629),
.A2(n_564),
.B(n_610),
.C(n_585),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_672),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_620),
.Y(n_688)
);

BUFx8_ASAP7_75t_L g689 ( 
.A(n_636),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_667),
.A2(n_564),
.B1(n_605),
.B2(n_596),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_656),
.B(n_650),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_659),
.B(n_605),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_615),
.A2(n_601),
.B(n_574),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_633),
.B(n_557),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_628),
.B(n_580),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_653),
.Y(n_696)
);

NOR3xp33_ASAP7_75t_L g697 ( 
.A(n_641),
.B(n_593),
.C(n_583),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_657),
.B(n_601),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_647),
.B(n_588),
.Y(n_699)
);

AO32x2_ASAP7_75t_L g700 ( 
.A1(n_625),
.A2(n_31),
.A3(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_630),
.B(n_31),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_642),
.A2(n_34),
.B1(n_41),
.B2(n_43),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_645),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_645),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_644),
.A2(n_44),
.B(n_45),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_626),
.A2(n_46),
.B(n_48),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_662),
.A2(n_49),
.B(n_51),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_654),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_660),
.B(n_52),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_648),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_614),
.B(n_213),
.Y(n_711)
);

NAND3xp33_ASAP7_75t_SL g712 ( 
.A(n_658),
.B(n_53),
.C(n_54),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_652),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_669),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_634),
.B(n_211),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_655),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_671),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_671),
.B(n_210),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_674),
.A2(n_63),
.B1(n_69),
.B2(n_71),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_643),
.B(n_209),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_670),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_665),
.A2(n_651),
.B(n_617),
.C(n_663),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_666),
.A2(n_639),
.B(n_631),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_675),
.B(n_623),
.Y(n_725)
);

BUFx4f_ASAP7_75t_L g726 ( 
.A(n_648),
.Y(n_726)
);

AOI21xp5_ASAP7_75t_L g727 ( 
.A1(n_638),
.A2(n_73),
.B(n_74),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_623),
.B(n_75),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_649),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_621),
.B(n_80),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_SL g731 ( 
.A(n_648),
.B(n_81),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_654),
.B(n_661),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_661),
.B(n_622),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_661),
.B(n_82),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_687),
.Y(n_735)
);

BUFx12f_ASAP7_75t_L g736 ( 
.A(n_677),
.Y(n_736)
);

BUFx12f_ASAP7_75t_L g737 ( 
.A(n_677),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_682),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_684),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_704),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_678),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_688),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_695),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_726),
.Y(n_744)
);

CKINVDCx11_ASAP7_75t_R g745 ( 
.A(n_680),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_726),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_682),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_689),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_708),
.B(n_732),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_692),
.B(n_664),
.Y(n_750)
);

BUFx2_ASAP7_75t_SL g751 ( 
.A(n_680),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_689),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_696),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_721),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_717),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_723),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_703),
.Y(n_757)
);

CKINVDCx16_ASAP7_75t_R g758 ( 
.A(n_681),
.Y(n_758)
);

INVx6_ASAP7_75t_SL g759 ( 
.A(n_731),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_691),
.Y(n_760)
);

INVx5_ASAP7_75t_L g761 ( 
.A(n_708),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_733),
.Y(n_762)
);

BUFx4f_ASAP7_75t_L g763 ( 
.A(n_714),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_725),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_734),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_700),
.B(n_664),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_698),
.B(n_622),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_730),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_728),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_679),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_699),
.Y(n_771)
);

BUFx4_ASAP7_75t_SL g772 ( 
.A(n_700),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_694),
.Y(n_773)
);

NAND2x1p5_ASAP7_75t_L g774 ( 
.A(n_685),
.B(n_646),
.Y(n_774)
);

INVx6_ASAP7_75t_SL g775 ( 
.A(n_731),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_718),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_690),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_710),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_715),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_700),
.B(n_668),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_686),
.Y(n_781)
);

BUFx12f_ASAP7_75t_L g782 ( 
.A(n_701),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_720),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_683),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_709),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_690),
.B(n_208),
.Y(n_786)
);

BUFx12f_ASAP7_75t_L g787 ( 
.A(n_702),
.Y(n_787)
);

CKINVDCx11_ASAP7_75t_R g788 ( 
.A(n_719),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_676),
.B(n_84),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_712),
.Y(n_790)
);

BUFx2_ASAP7_75t_SL g791 ( 
.A(n_719),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_711),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_729),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_705),
.Y(n_794)
);

BUFx2_ASAP7_75t_SL g795 ( 
.A(n_729),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_697),
.B(n_207),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_693),
.B(n_85),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_707),
.Y(n_798)
);

AOI221xp5_ASAP7_75t_L g799 ( 
.A1(n_780),
.A2(n_713),
.B1(n_716),
.B2(n_706),
.C(n_722),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_735),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_786),
.A2(n_727),
.B(n_724),
.Y(n_801)
);

OA21x2_ASAP7_75t_L g802 ( 
.A1(n_781),
.A2(n_86),
.B(n_87),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_768),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_750),
.B(n_753),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_789),
.A2(n_89),
.B(n_91),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_735),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_773),
.B(n_92),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_798),
.A2(n_93),
.B(n_94),
.Y(n_808)
);

INVx2_ASAP7_75t_R g809 ( 
.A(n_772),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_795),
.B(n_95),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_750),
.B(n_96),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_755),
.B(n_99),
.Y(n_812)
);

AO21x2_ASAP7_75t_L g813 ( 
.A1(n_780),
.A2(n_101),
.B(n_102),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_760),
.B(n_103),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_760),
.B(n_777),
.Y(n_815)
);

INVx6_ASAP7_75t_SL g816 ( 
.A(n_749),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_792),
.B(n_104),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_788),
.A2(n_782),
.B1(n_787),
.B2(n_793),
.Y(n_818)
);

OAI22xp33_ASAP7_75t_L g819 ( 
.A1(n_793),
.A2(n_107),
.B1(n_108),
.B2(n_112),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_773),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_788),
.A2(n_782),
.B1(n_787),
.B2(n_784),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_754),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_762),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_756),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_739),
.Y(n_825)
);

OR2x6_ASAP7_75t_L g826 ( 
.A(n_791),
.B(n_114),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_756),
.B(n_115),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_745),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_764),
.B(n_118),
.Y(n_829)
);

BUFx10_ASAP7_75t_L g830 ( 
.A(n_752),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_743),
.Y(n_831)
);

OAI21x1_ASAP7_75t_SL g832 ( 
.A1(n_738),
.A2(n_120),
.B(n_121),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_739),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_770),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_789),
.A2(n_125),
.B(n_127),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_741),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_771),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_762),
.Y(n_838)
);

OA21x2_ASAP7_75t_L g839 ( 
.A1(n_796),
.A2(n_128),
.B(n_129),
.Y(n_839)
);

OAI21x1_ASAP7_75t_L g840 ( 
.A1(n_798),
.A2(n_130),
.B(n_131),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_764),
.B(n_132),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_762),
.B(n_749),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_784),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_763),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_766),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_763),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_846)
);

OAI21x1_ASAP7_75t_L g847 ( 
.A1(n_798),
.A2(n_143),
.B(n_144),
.Y(n_847)
);

BUFx12f_ASAP7_75t_L g848 ( 
.A(n_745),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_736),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_763),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_759),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_765),
.B(n_151),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_776),
.B(n_153),
.Y(n_853)
);

OAI21x1_ASAP7_75t_L g854 ( 
.A1(n_774),
.A2(n_156),
.B(n_157),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_815),
.A2(n_784),
.B1(n_790),
.B2(n_779),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_848),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_809),
.A2(n_775),
.B1(n_759),
.B2(n_790),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_823),
.Y(n_858)
);

AO21x2_ASAP7_75t_L g859 ( 
.A1(n_801),
.A2(n_766),
.B(n_778),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_831),
.Y(n_860)
);

NAND2x1p5_ASAP7_75t_L g861 ( 
.A(n_850),
.B(n_768),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_808),
.A2(n_774),
.B(n_768),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_831),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_836),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_803),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_837),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_803),
.B(n_769),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_833),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_803),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_851),
.Y(n_870)
);

OAI21x1_ASAP7_75t_L g871 ( 
.A1(n_808),
.A2(n_785),
.B(n_797),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_834),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_822),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_838),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_828),
.Y(n_875)
);

OR2x6_ASAP7_75t_L g876 ( 
.A(n_810),
.B(n_790),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_818),
.A2(n_790),
.B1(n_742),
.B2(n_759),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_838),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_804),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_824),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_816),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_806),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_810),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_820),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_842),
.B(n_785),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_840),
.A2(n_785),
.B(n_797),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_810),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_845),
.B(n_776),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_800),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_800),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_845),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_825),
.B(n_769),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_849),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_816),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_849),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_818),
.A2(n_775),
.B1(n_748),
.B2(n_758),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_879),
.B(n_821),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_896),
.A2(n_814),
.B(n_821),
.C(n_817),
.Y(n_898)
);

AND2x2_ASAP7_75t_SL g899 ( 
.A(n_883),
.B(n_809),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_868),
.Y(n_900)
);

OAI22xp33_ASAP7_75t_L g901 ( 
.A1(n_876),
.A2(n_826),
.B1(n_805),
.B2(n_835),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_875),
.B(n_828),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_R g903 ( 
.A(n_875),
.B(n_752),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_860),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_863),
.Y(n_905)
);

AND2x4_ASAP7_75t_SL g906 ( 
.A(n_883),
.B(n_850),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_858),
.B(n_885),
.Y(n_907)
);

NOR3xp33_ASAP7_75t_SL g908 ( 
.A(n_856),
.B(n_814),
.C(n_817),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_865),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_891),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_864),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_866),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_867),
.B(n_748),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_R g914 ( 
.A(n_856),
.B(n_848),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_893),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_874),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_889),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_865),
.B(n_813),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_869),
.B(n_813),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_R g920 ( 
.A(n_895),
.B(n_736),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_868),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_890),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_R g923 ( 
.A(n_883),
.B(n_737),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_907),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_L g925 ( 
.A(n_908),
.B(n_884),
.C(n_892),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_907),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_910),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_910),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_904),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_905),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_909),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_911),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_912),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_909),
.B(n_859),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_917),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_915),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_901),
.A2(n_775),
.B1(n_897),
.B2(n_783),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_900),
.B(n_859),
.Y(n_938)
);

OAI33xp33_ASAP7_75t_L g939 ( 
.A1(n_921),
.A2(n_872),
.A3(n_877),
.B1(n_880),
.B2(n_873),
.B3(n_882),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_916),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_900),
.B(n_867),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_918),
.B(n_867),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_917),
.Y(n_943)
);

NAND4xp25_ASAP7_75t_L g944 ( 
.A(n_898),
.B(n_869),
.C(n_855),
.D(n_799),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_918),
.B(n_919),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_916),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_939),
.Y(n_947)
);

AOI211xp5_ASAP7_75t_L g948 ( 
.A1(n_944),
.A2(n_919),
.B(n_819),
.C(n_887),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_930),
.Y(n_949)
);

OAI221xp5_ASAP7_75t_L g950 ( 
.A1(n_937),
.A2(n_876),
.B1(n_857),
.B2(n_826),
.C(n_887),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_942),
.A2(n_899),
.B(n_876),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_936),
.A2(n_876),
.B1(n_899),
.B2(n_921),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_930),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_924),
.B(n_926),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_946),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_936),
.Y(n_956)
);

OAI211xp5_ASAP7_75t_L g957 ( 
.A1(n_925),
.A2(n_902),
.B(n_920),
.C(n_903),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_934),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_931),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_934),
.Y(n_960)
);

OAI211xp5_ASAP7_75t_L g961 ( 
.A1(n_940),
.A2(n_914),
.B(n_923),
.C(n_915),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_954),
.B(n_927),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_947),
.A2(n_941),
.B(n_826),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_949),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_956),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_953),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_947),
.B(n_932),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_955),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_959),
.Y(n_969)
);

OAI31xp33_ASAP7_75t_SL g970 ( 
.A1(n_961),
.A2(n_945),
.A3(n_913),
.B(n_933),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_958),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_956),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_959),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_955),
.B(n_945),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_972),
.B(n_913),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_972),
.B(n_948),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_967),
.B(n_962),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_962),
.B(n_928),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_965),
.B(n_913),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_970),
.B(n_940),
.Y(n_980)
);

INVxp67_ASAP7_75t_SL g981 ( 
.A(n_963),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_964),
.B(n_929),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_974),
.B(n_957),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_982),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_982),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_975),
.B(n_969),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_983),
.B(n_973),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_978),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_979),
.B(n_974),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_977),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_989),
.B(n_976),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_987),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_990),
.B(n_981),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_987),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_990),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_988),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_990),
.B(n_966),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_984),
.A2(n_980),
.B(n_966),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_985),
.B(n_830),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_L g1000 ( 
.A(n_988),
.B(n_952),
.C(n_971),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_994),
.B(n_986),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_992),
.B(n_986),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_995),
.B(n_968),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_991),
.B(n_968),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_993),
.B(n_968),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_996),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_991),
.B(n_830),
.Y(n_1007)
);

NOR4xp25_ASAP7_75t_L g1008 ( 
.A(n_997),
.B(n_998),
.C(n_999),
.D(n_971),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1001),
.Y(n_1009)
);

NAND4xp25_ASAP7_75t_L g1010 ( 
.A(n_1002),
.B(n_1000),
.C(n_951),
.D(n_740),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_1006),
.A2(n_960),
.B(n_958),
.C(n_844),
.Y(n_1011)
);

NAND3xp33_ASAP7_75t_L g1012 ( 
.A(n_1005),
.B(n_843),
.C(n_960),
.Y(n_1012)
);

AOI322xp5_ASAP7_75t_L g1013 ( 
.A1(n_1008),
.A2(n_887),
.A3(n_843),
.B1(n_853),
.B2(n_812),
.C1(n_938),
.C2(n_935),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1007),
.A2(n_938),
.B1(n_950),
.B2(n_887),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_1004),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_1003),
.A2(n_870),
.B(n_946),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1009),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1015),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_1012),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1011),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1013),
.B(n_946),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1010),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1018),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1017),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_1020),
.B(n_1016),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_1022),
.B(n_830),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1019),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1021),
.B(n_1014),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1021),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1018),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1027),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1023),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_L g1033 ( 
.A(n_1030),
.B(n_740),
.C(n_807),
.Y(n_1033)
);

NAND3xp33_ASAP7_75t_L g1034 ( 
.A(n_1024),
.B(n_1025),
.C(n_1029),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1028),
.B(n_943),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_1028),
.B(n_737),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1026),
.B(n_916),
.Y(n_1037)
);

NOR4xp25_ASAP7_75t_L g1038 ( 
.A(n_1027),
.B(n_829),
.C(n_827),
.D(n_853),
.Y(n_1038)
);

AOI211xp5_ASAP7_75t_L g1039 ( 
.A1(n_1034),
.A2(n_751),
.B(n_746),
.C(n_846),
.Y(n_1039)
);

AND5x1_ASAP7_75t_L g1040 ( 
.A(n_1036),
.B(n_870),
.C(n_906),
.D(n_832),
.E(n_746),
.Y(n_1040)
);

AOI221xp5_ASAP7_75t_L g1041 ( 
.A1(n_1031),
.A2(n_783),
.B1(n_859),
.B2(n_811),
.C(n_887),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_1032),
.A2(n_757),
.B1(n_744),
.B2(n_839),
.Y(n_1042)
);

OAI221xp5_ASAP7_75t_L g1043 ( 
.A1(n_1035),
.A2(n_839),
.B1(n_744),
.B2(n_802),
.C(n_757),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_1039),
.A2(n_1033),
.B1(n_1037),
.B2(n_1038),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1042),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_1040),
.A2(n_839),
.B(n_802),
.C(n_841),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1041),
.A2(n_757),
.B1(n_906),
.B2(n_802),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_1043),
.A2(n_852),
.B(n_747),
.C(n_861),
.Y(n_1048)
);

OAI221xp5_ASAP7_75t_L g1049 ( 
.A1(n_1039),
.A2(n_757),
.B1(n_738),
.B2(n_861),
.C(n_894),
.Y(n_1049)
);

NAND4xp25_ASAP7_75t_SL g1050 ( 
.A(n_1039),
.B(n_738),
.C(n_888),
.D(n_922),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_1041),
.A2(n_765),
.B1(n_749),
.B2(n_852),
.Y(n_1051)
);

INVxp33_ASAP7_75t_L g1052 ( 
.A(n_1042),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_1044),
.B(n_747),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_1045),
.A2(n_852),
.B1(n_747),
.B2(n_765),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_L g1055 ( 
.A(n_1052),
.B(n_761),
.C(n_765),
.Y(n_1055)
);

AOI322xp5_ASAP7_75t_L g1056 ( 
.A1(n_1051),
.A2(n_881),
.A3(n_894),
.B1(n_794),
.B2(n_888),
.C1(n_922),
.C2(n_878),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_1050),
.Y(n_1057)
);

NOR4xp75_ASAP7_75t_L g1058 ( 
.A(n_1049),
.B(n_878),
.C(n_874),
.D(n_160),
.Y(n_1058)
);

OAI211xp5_ASAP7_75t_L g1059 ( 
.A1(n_1048),
.A2(n_840),
.B(n_847),
.C(n_854),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1047),
.Y(n_1060)
);

NOR2x1_ASAP7_75t_L g1061 ( 
.A(n_1046),
.B(n_881),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1060),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_1057),
.Y(n_1063)
);

NAND4xp75_ASAP7_75t_L g1064 ( 
.A(n_1061),
.B(n_158),
.C(n_159),
.D(n_161),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_1053),
.B(n_761),
.C(n_794),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1058),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_1055),
.B(n_854),
.C(n_847),
.Y(n_1067)
);

NOR3x2_ASAP7_75t_L g1068 ( 
.A(n_1059),
.B(n_162),
.C(n_163),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1054),
.Y(n_1069)
);

AOI211xp5_ASAP7_75t_L g1070 ( 
.A1(n_1056),
.A2(n_871),
.B(n_886),
.C(n_862),
.Y(n_1070)
);

AND4x1_ASAP7_75t_L g1071 ( 
.A(n_1061),
.B(n_165),
.C(n_166),
.D(n_167),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_1057),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1060),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_L g1074 ( 
.A(n_1060),
.B(n_886),
.C(n_871),
.Y(n_1074)
);

NOR2xp67_ASAP7_75t_L g1075 ( 
.A(n_1063),
.B(n_168),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_1072),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1062),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_1064),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_1063),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_1073),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_1066),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_1069),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_1071),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1076),
.Y(n_1084)
);

OA22x2_ASAP7_75t_L g1085 ( 
.A1(n_1079),
.A2(n_1068),
.B1(n_1065),
.B2(n_1070),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1080),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_1077),
.B(n_1067),
.C(n_1074),
.Y(n_1087)
);

OAI22x1_ASAP7_75t_L g1088 ( 
.A1(n_1083),
.A2(n_861),
.B1(n_767),
.B2(n_761),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_1082),
.Y(n_1089)
);

CKINVDCx16_ASAP7_75t_R g1090 ( 
.A(n_1089),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_SL g1091 ( 
.A1(n_1084),
.A2(n_1081),
.B1(n_1078),
.B2(n_1075),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1086),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1090),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_1093),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1094),
.A2(n_1092),
.B(n_1091),
.Y(n_1095)
);

NAND5xp2_ASAP7_75t_L g1096 ( 
.A(n_1095),
.B(n_1085),
.C(n_1087),
.D(n_1088),
.E(n_174),
.Y(n_1096)
);

OAI221xp5_ASAP7_75t_SL g1097 ( 
.A1(n_1095),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.C(n_175),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1096),
.A2(n_177),
.B(n_179),
.Y(n_1098)
);

AOI31xp33_ASAP7_75t_L g1099 ( 
.A1(n_1097),
.A2(n_180),
.A3(n_182),
.B(n_183),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1098),
.A2(n_761),
.B1(n_767),
.B2(n_862),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_SL g1101 ( 
.A1(n_1099),
.A2(n_185),
.B1(n_189),
.B2(n_193),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1101),
.A2(n_194),
.B(n_197),
.Y(n_1102)
);

AOI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1102),
.A2(n_1100),
.B1(n_199),
.B2(n_201),
.C(n_202),
.Y(n_1103)
);

AOI211xp5_ASAP7_75t_L g1104 ( 
.A1(n_1103),
.A2(n_198),
.B(n_203),
.C(n_206),
.Y(n_1104)
);


endmodule