module fake_netlist_6_710_n_29 (n_7, n_6, n_4, n_2, n_3, n_5, n_1, n_0, n_9, n_8, n_29);

input n_7;
input n_6;
input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;
input n_9;
input n_8;

output n_29;

wire n_16;
wire n_18;
wire n_10;
wire n_21;
wire n_24;
wire n_15;
wire n_27;
wire n_14;
wire n_22;
wire n_26;
wire n_13;
wire n_11;
wire n_28;
wire n_23;
wire n_17;
wire n_12;
wire n_20;
wire n_19;
wire n_25;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_8),
.B(n_3),
.Y(n_10)
);

AND2x2_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_5),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_L g12 ( 
.A1(n_1),
.A2(n_6),
.B1(n_9),
.B2(n_8),
.Y(n_12)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_9),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_5),
.B(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

OAI21x1_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_16),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_2),
.Y(n_19)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_2),
.B(n_7),
.Y(n_20)
);

OAI211xp5_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_12),
.B(n_15),
.C(n_10),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

AOI221xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_10),
.B1(n_15),
.B2(n_13),
.C(n_11),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_17),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_17),
.B(n_21),
.C(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_24),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_26),
.B1(n_13),
.B2(n_7),
.Y(n_28)
);

AOI222xp33_ASAP7_75t_SL g29 ( 
.A1(n_28),
.A2(n_2),
.B1(n_4),
.B2(n_13),
.C1(n_15),
.C2(n_16),
.Y(n_29)
);


endmodule