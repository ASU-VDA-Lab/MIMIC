module fake_jpeg_31666_n_25 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_25);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_25;

wire n_13;
wire n_21;
wire n_23;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_8),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_9),
.Y(n_13)
);

CKINVDCx9p33_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_13),
.B(n_0),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_13),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_15),
.C(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_20),
.B(n_11),
.Y(n_22)
);

AOI21x1_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_23),
.B(n_21),
.Y(n_24)
);

AOI322xp5_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_1),
.A3(n_2),
.B1(n_5),
.B2(n_6),
.C1(n_10),
.C2(n_22),
.Y(n_25)
);


endmodule