module fake_jpeg_30769_n_49 (n_3, n_2, n_1, n_0, n_4, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

AOI21xp33_ASAP7_75t_L g12 ( 
.A1(n_3),
.A2(n_5),
.B(n_4),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_0),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_16),
.C(n_17),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_8),
.B1(n_7),
.B2(n_9),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_2),
.C(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_19),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_13),
.B(n_10),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_7),
.A2(n_8),
.B1(n_11),
.B2(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_R g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_14),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_17),
.B(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_25),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_36),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_23),
.C(n_20),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_34),
.C(n_15),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_32),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_11),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_26),
.B(n_30),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_45),
.C(n_39),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_47),
.B(n_13),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_14),
.B(n_13),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_14),
.B(n_13),
.Y(n_49)
);


endmodule