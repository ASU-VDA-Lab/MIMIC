module real_jpeg_3760_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_1),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_1),
.B(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_1),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_1),
.B(n_57),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_1),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_1),
.B(n_88),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_1),
.B(n_280),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_2),
.Y(n_106)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_2),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_3),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_3),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_3),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_3),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_3),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_3),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_4),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_4),
.B(n_51),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_4),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_4),
.B(n_446),
.Y(n_445)
);

NAND2x1_ASAP7_75t_SL g461 ( 
.A(n_4),
.B(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_5),
.Y(n_353)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_7),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_7),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_7),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_7),
.B(n_265),
.Y(n_264)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_8),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_8),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_9),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_9),
.B(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_9),
.B(n_364),
.Y(n_363)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_11),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_11),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_11),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_11),
.B(n_190),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_11),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_11),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_11),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_11),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_42),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_12),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_12),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_12),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_12),
.B(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_12),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_12),
.B(n_101),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_12),
.B(n_465),
.Y(n_464)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_13),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_14),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_14),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_14),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_14),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_14),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_14),
.B(n_379),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_15),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_451),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_423),
.B(n_450),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_270),
.B(n_309),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_227),
.B(n_269),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_197),
.B(n_226),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_22),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_152),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_23),
.B(n_152),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_102),
.C(n_138),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_24),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_71),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_25),
.B(n_72),
.C(n_85),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_46),
.C(n_60),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_26),
.B(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_34),
.B2(n_40),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_28),
.A2(n_29),
.B1(n_431),
.B2(n_432),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_28),
.A2(n_29),
.B1(n_73),
.B2(n_74),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_29),
.B(n_34),
.C(n_41),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_29),
.B(n_206),
.C(n_433),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_48),
.Y(n_47)
);

OR2x2_ASAP7_75t_SL g74 ( 
.A(n_30),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_30),
.B(n_279),
.Y(n_278)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_32),
.Y(n_148)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_32),
.Y(n_332)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_33),
.Y(n_195)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_33),
.Y(n_366)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_38),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_38),
.Y(n_162)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_39),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_39),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_39),
.Y(n_447)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_46),
.A2(n_60),
.B1(n_61),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_46),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.C(n_54),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_47),
.A2(n_54),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_47),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_47),
.A2(n_206),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_47),
.A2(n_206),
.B1(n_433),
.B2(n_434),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_47),
.B(n_124),
.C(n_278),
.Y(n_437)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_50),
.B(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_53),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_54),
.Y(n_207)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_58),
.Y(n_219)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_59),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_59),
.Y(n_290)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_59),
.Y(n_337)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_62),
.A2(n_177),
.B1(n_178),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_180),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_62),
.B(n_178),
.C(n_181),
.Y(n_267)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_65),
.Y(n_376)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

BUFx8_ASAP7_75t_L g320 ( 
.A(n_66),
.Y(n_320)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_85),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_74),
.B(n_78),
.C(n_83),
.Y(n_196)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_79),
.B(n_124),
.Y(n_326)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_81),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_85),
.Y(n_477)
);

FAx1_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_93),
.CI(n_98),
.CON(n_85),
.SN(n_85)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_87),
.B(n_91),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_86),
.B(n_93),
.C(n_98),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_99),
.B(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g463 ( 
.A(n_101),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_102),
.B(n_138),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_119),
.C(n_121),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_103),
.A2(n_119),
.B1(n_120),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_108),
.C(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_105),
.B(n_383),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_105),
.B(n_369),
.Y(n_389)
);

INVx8_ASAP7_75t_L g465 ( 
.A(n_106),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_118),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_111),
.A2(n_112),
.B1(n_247),
.B2(n_251),
.Y(n_246)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_112),
.B(n_178),
.C(n_248),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_116),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_117),
.Y(n_325)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_121),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_128),
.C(n_133),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_122),
.A2(n_123),
.B1(n_410),
.B2(n_411),
.Y(n_409)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_124),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_124),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_124),
.A2(n_236),
.B1(n_278),
.B2(n_281),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_124),
.B(n_239),
.C(n_245),
.Y(n_283)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_134),
.Y(n_411)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_131),
.Y(n_356)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_151),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_141),
.C(n_151),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_147),
.C(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_147),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_147),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_153),
.B(n_155),
.C(n_183),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_183),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_174),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_157),
.B(n_158),
.C(n_174),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_159),
.Y(n_234)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_164),
.B(n_169),
.C(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_173),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_181),
.B2(n_182),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_177),
.A2(n_178),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_177),
.A2(n_178),
.B1(n_317),
.B2(n_318),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_178),
.B(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_181),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_181),
.A2(n_182),
.B1(n_445),
.B2(n_448),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_182),
.B(n_443),
.C(n_445),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_184),
.B(n_186),
.C(n_187),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_189),
.B(n_193),
.C(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_191),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_224),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_198),
.B(n_224),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.C(n_221),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_199),
.A2(n_200),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_203),
.B(n_221),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.C(n_220),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_204),
.B(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_208),
.B(n_220),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.C(n_215),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_212),
.B(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_215),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_216),
.B(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_216),
.B(n_386),
.Y(n_385)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_228),
.B(n_270),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_271),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_230),
.B(n_271),
.Y(n_422)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_252),
.CI(n_268),
.CON(n_230),
.SN(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_246),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_233),
.B(n_235),
.C(n_246),
.Y(n_296)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_245),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_241),
.A2(n_245),
.B1(n_471),
.B2(n_472),
.Y(n_470)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_248),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_255),
.C(n_257),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_267),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_264),
.B2(n_266),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_264),
.C(n_267),
.Y(n_299)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_264),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_264),
.A2(n_266),
.B1(n_305),
.B2(n_308),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_266),
.B(n_301),
.C(n_308),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_272),
.B(n_274),
.C(n_294),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_294),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_282),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_275),
.B(n_283),
.C(n_284),
.Y(n_449)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_293),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_286),
.B(n_288),
.C(n_292),
.Y(n_438)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_288),
.Y(n_291)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_295),
.B(n_299),
.C(n_300),
.Y(n_426)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

AO22x1_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_305),
.Y(n_308)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI31xp33_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_419),
.A3(n_420),
.B(n_422),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_413),
.B(n_418),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_400),
.B(n_412),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_358),
.B(n_399),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_344),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_314),
.B(n_344),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_327),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_315),
.B(n_328),
.C(n_341),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_316),
.B(n_322),
.C(n_326),
.Y(n_408)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_341),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.C(n_338),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_329),
.B(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_333),
.A2(n_334),
.B1(n_338),
.B2(n_339),
.Y(n_346)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.C(n_357),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_345),
.B(n_396),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_347),
.A2(n_348),
.B1(n_357),
.B2(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_354),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_349),
.A2(n_350),
.B1(n_354),
.B2(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_357),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_393),
.B(n_398),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_380),
.B(n_392),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_371),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_371),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_370),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_367),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_367),
.C(n_370),
.Y(n_394)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_377),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_372),
.A2(n_373),
.B1(n_377),
.B2(n_378),
.Y(n_390)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_388),
.B(n_391),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_389),
.B(n_390),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_394),
.B(n_395),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_402),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_404),
.B1(n_406),
.B2(n_407),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_408),
.C(n_409),
.Y(n_417)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_417),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_417),
.Y(n_418)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_415),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_425),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_428),
.C(n_439),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_439),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_435),
.B2(n_436),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_437),
.C(n_438),
.Y(n_456)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_433),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_449),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_442),
.C(n_449),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_445),
.Y(n_448)
);

INVx6_ASAP7_75t_SL g446 ( 
.A(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_473),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_454),
.Y(n_474)
);

BUFx24_ASAP7_75t_SL g475 ( 
.A(n_454),
.Y(n_475)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_456),
.CI(n_457),
.CON(n_454),
.SN(n_454)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_468),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_461),
.A2(n_464),
.B1(n_466),
.B2(n_467),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_461),
.Y(n_466)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g467 ( 
.A(n_464),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);


endmodule