module fake_jpeg_7129_n_231 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_7),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_16),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_16),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_27),
.B(n_25),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_59),
.B(n_35),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_29),
.C(n_30),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_45),
.C(n_38),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_16),
.B1(n_15),
.B2(n_32),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_44),
.B1(n_45),
.B2(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_60),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_15),
.B1(n_31),
.B2(n_17),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_15),
.B1(n_31),
.B2(n_17),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_37),
.B(n_18),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_32),
.B1(n_21),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_35),
.B1(n_20),
.B2(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_67),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_34),
.B1(n_40),
.B2(n_54),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_52),
.B(n_42),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_75),
.C(n_21),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_79),
.B1(n_41),
.B2(n_34),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_44),
.B(n_41),
.C(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_77),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_37),
.B(n_19),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_22),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_59),
.B1(n_49),
.B2(n_52),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_85),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_93),
.B(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_86),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_87),
.B(n_22),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_51),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_68),
.B(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_93),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_91),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_66),
.B(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_78),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_87),
.B1(n_94),
.B2(n_51),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_102),
.B(n_109),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_74),
.B(n_69),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_111),
.C(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_47),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_87),
.Y(n_119)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_114),
.C(n_72),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_84),
.A3(n_88),
.B1(n_89),
.B2(n_86),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_107),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_130),
.B1(n_109),
.B2(n_105),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_88),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_111),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_112),
.A2(n_97),
.B1(n_85),
.B2(n_82),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_129),
.B1(n_131),
.B2(n_104),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_97),
.C(n_47),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_133),
.C(n_102),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_87),
.B1(n_29),
.B2(n_50),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_64),
.C(n_77),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_50),
.B1(n_95),
.B2(n_19),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_139),
.C(n_141),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_106),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_148),
.B1(n_20),
.B2(n_72),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_144),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_98),
.C(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_146),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_26),
.B(n_30),
.C(n_29),
.D(n_105),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_143),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_30),
.C(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_71),
.B1(n_24),
.B2(n_20),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_71),
.B1(n_50),
.B2(n_14),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_117),
.C(n_121),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_150),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_71),
.B1(n_22),
.B2(n_24),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_115),
.C(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_154),
.B(n_160),
.Y(n_178)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

INVxp33_ASAP7_75t_SL g176 ( 
.A(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_166),
.C(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_168),
.B(n_135),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_139),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_172),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_164),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_57),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_143),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_181),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_134),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_170),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_18),
.Y(n_190)
);

OAI21x1_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_95),
.B(n_36),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_159),
.B1(n_163),
.B2(n_155),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_197),
.B1(n_180),
.B2(n_182),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_192),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_194),
.C(n_8),
.Y(n_203)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_193),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_1),
.B(n_2),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_1),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_9),
.C(n_12),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_61),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_1),
.Y(n_207)
);

AO221x1_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_61),
.B1(n_14),
.B2(n_3),
.C(n_4),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_173),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_198),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_177),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_9),
.C(n_11),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_179),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_204),
.B(n_202),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_8),
.B(n_11),
.C(n_10),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_205),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_14),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_2),
.Y(n_213)
);

NOR2x1_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_6),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_214),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_6),
.B(n_11),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_216),
.A2(n_217),
.B(n_222),
.C(n_220),
.Y(n_224)
);

AOI211x1_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_206),
.B(n_10),
.C(n_6),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_221),
.C(n_212),
.Y(n_223)
);

AOI21x1_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_2),
.B(n_3),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_12),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_224),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_226),
.B(n_3),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_3),
.Y(n_229)
);

NAND4xp25_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_4),
.C(n_228),
.D(n_208),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_4),
.Y(n_231)
);


endmodule