module real_jpeg_26589_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_4),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_5),
.A2(n_37),
.B1(n_43),
.B2(n_62),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_5),
.A2(n_23),
.B1(n_26),
.B2(n_62),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_64),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_7),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.Y(n_88)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_37),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_53),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_9),
.A2(n_23),
.B1(n_26),
.B2(n_53),
.Y(n_125)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_37),
.B1(n_43),
.B2(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_43),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_12),
.A2(n_42),
.B(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_12),
.B(n_73),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_12),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_12),
.A2(n_23),
.B(n_58),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_12),
.B(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_12),
.A2(n_31),
.B1(n_110),
.B2(n_125),
.Y(n_127)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_91),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_90),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_65),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_18),
.B(n_65),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_45),
.C(n_54),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_19),
.A2(n_20),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_34),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_30),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_22),
.B(n_28),
.Y(n_112)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_23),
.A2(n_26),
.B1(n_58),
.B2(n_59),
.Y(n_60)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_26),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_27),
.A2(n_28),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_31),
.A2(n_110),
.B1(n_117),
.B2(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_31),
.B(n_98),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.A3(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_36),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_40),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_36),
.A2(n_59),
.B(n_98),
.C(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_37),
.A2(n_43),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_45),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_50),
.B1(n_52),
.B2(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_63),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_60),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_56),
.A2(n_60),
.B1(n_61),
.B2(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_60),
.B(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_83),
.B2(n_84),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_133),
.B(n_138),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_113),
.B(n_132),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_96),
.B1(n_100),
.B2(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_108),
.C(n_109),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B(n_112),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_121),
.B(n_131),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_119),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_126),
.B(n_130),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_123),
.B(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_135),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);


endmodule