module fake_jpeg_6613_n_268 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_268);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_268;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_91;
wire n_33;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g81 ( 
.A(n_37),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_41),
.B(n_43),
.Y(n_80)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g90 ( 
.A(n_42),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_7),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_32),
.Y(n_56)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_50),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_19),
.B1(n_15),
.B2(n_29),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_51),
.A2(n_76),
.B1(n_79),
.B2(n_91),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_55),
.B(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_72),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_86),
.Y(n_110)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_39),
.A2(n_27),
.B1(n_30),
.B2(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_32),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_77),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_34),
.A2(n_21),
.B1(n_18),
.B2(n_27),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_34),
.A2(n_28),
.B1(n_31),
.B2(n_17),
.Y(n_79)
);

CKINVDCx6p67_ASAP7_75t_R g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_28),
.C(n_21),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_9),
.B(n_8),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_21),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_44),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_48),
.A2(n_18),
.B1(n_31),
.B2(n_17),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_16),
.B1(n_31),
.B2(n_18),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_37),
.A2(n_31),
.B1(n_16),
.B2(n_8),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_95),
.B1(n_10),
.B2(n_3),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_37),
.A2(n_16),
.B1(n_8),
.B2(n_9),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_38),
.B(n_16),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_97),
.B(n_12),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_38),
.B(n_13),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_99),
.B(n_118),
.Y(n_135)
);

NAND2xp33_ASAP7_75t_SL g105 ( 
.A(n_50),
.B(n_9),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_105),
.B(n_79),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_80),
.B(n_57),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_68),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_83),
.B1(n_54),
.B2(n_75),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_89),
.C(n_85),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_127),
.C(n_134),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_56),
.C(n_68),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_68),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_128),
.B(n_150),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_55),
.Y(n_129)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_61),
.B1(n_65),
.B2(n_82),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_130),
.A2(n_146),
.B1(n_113),
.B2(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_125),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_87),
.Y(n_132)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_55),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_135),
.B(n_139),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_87),
.Y(n_136)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_141),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_102),
.B(n_58),
.Y(n_142)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_144),
.Y(n_178)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_90),
.Y(n_145)
);

XNOR2x2_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_83),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_84),
.B1(n_65),
.B2(n_82),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_74),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_104),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_54),
.B(n_83),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_60),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_152),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_114),
.B1(n_119),
.B2(n_100),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_150),
.B1(n_128),
.B2(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_70),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_90),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_69),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_147),
.A2(n_98),
.B1(n_72),
.B2(n_73),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_160),
.A2(n_169),
.B1(n_180),
.B2(n_189),
.Y(n_202)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_166),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_151),
.B(n_144),
.Y(n_191)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_168),
.A2(n_174),
.B1(n_149),
.B2(n_53),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_SL g192 ( 
.A1(n_170),
.A2(n_138),
.B(n_143),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_124),
.B1(n_119),
.B2(n_81),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_81),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_135),
.C(n_155),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_145),
.A2(n_100),
.B1(n_117),
.B2(n_109),
.Y(n_180)
);

BUFx4f_ASAP7_75t_SL g181 ( 
.A(n_141),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_188),
.Y(n_190)
);

AO22x1_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_69),
.B1(n_93),
.B2(n_71),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_187),
.A2(n_139),
.B(n_133),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_126),
.A2(n_117),
.B1(n_109),
.B2(n_104),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_180),
.CI(n_189),
.CON(n_217),
.SN(n_217)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_192),
.A2(n_175),
.B1(n_159),
.B2(n_187),
.Y(n_215)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_198),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_152),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_148),
.Y(n_196)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_133),
.B(n_127),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_201),
.B(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_164),
.B(n_128),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_204),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_153),
.C(n_158),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_184),
.C(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_206),
.C(n_207),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_140),
.C(n_69),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_53),
.C(n_149),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_182),
.B1(n_160),
.B2(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_211),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_1),
.B(n_3),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_179),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_226),
.B1(n_227),
.B2(n_201),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_174),
.B1(n_176),
.B2(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_213),
.B(n_228),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_216),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_179),
.B1(n_185),
.B2(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_224),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_206),
.C(n_193),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_181),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_223),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_161),
.C(n_183),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_166),
.B1(n_183),
.B2(n_163),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_163),
.B1(n_62),
.B2(n_103),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_228),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_191),
.A3(n_203),
.B1(n_210),
.B2(n_205),
.C1(n_197),
.C2(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_196),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_242),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_212),
.A2(n_209),
.B1(n_195),
.B2(n_198),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_211),
.B(n_194),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_218),
.C(n_222),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_247),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_239),
.A2(n_226),
.B1(n_215),
.B2(n_218),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_237),
.C(n_243),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_219),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_251),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_216),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_232),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_239),
.B1(n_238),
.B2(n_233),
.Y(n_255)
);

AOI211xp5_ASAP7_75t_L g260 ( 
.A1(n_255),
.A2(n_258),
.B(n_225),
.C(n_247),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_214),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_230),
.C(n_225),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_224),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_260),
.B(n_252),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_244),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_254),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_249),
.C(n_245),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_253),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_264),
.B(n_265),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_231),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_262),
.Y(n_268)
);


endmodule