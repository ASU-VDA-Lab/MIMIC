module real_jpeg_23400_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_16;

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_0),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_15)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_0),
.A2(n_18),
.B1(n_33),
.B2(n_38),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_3),
.A2(n_33),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_3),
.A2(n_16),
.B1(n_17),
.B2(n_45),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_17),
.C(n_31),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_4),
.A2(n_26),
.B1(n_50),
.B2(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_4),
.B(n_67),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_6),
.A2(n_16),
.B1(n_17),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_6),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_16),
.B1(n_17),
.B2(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_59),
.Y(n_10)
);

AOI21xp33_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_46),
.B(n_58),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_28),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_13),
.B(n_28),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_15),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_16),
.A2(n_17),
.B1(n_31),
.B2(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_16),
.B(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_23),
.A2(n_51),
.B(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_29),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_33),
.B1(n_38),
.B2(n_41),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_33),
.A2(n_38),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_42),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_43),
.B1(n_44),
.B2(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_42),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_57),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_78),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_63),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_73),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_70),
.B2(n_72),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);


endmodule