module fake_jpeg_5693_n_232 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_232);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_5),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_33),
.Y(n_52)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_36),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_25),
.Y(n_50)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_20),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_20),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_29),
.A2(n_19),
.B1(n_21),
.B2(n_16),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_19),
.B1(n_24),
.B2(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_13),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_40),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_15),
.B1(n_16),
.B2(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_15),
.B1(n_21),
.B2(n_24),
.Y(n_60)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_58),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_60),
.B1(n_38),
.B2(n_27),
.Y(n_85)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_65),
.Y(n_89)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_52),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_24),
.B1(n_19),
.B2(n_27),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_42),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_26),
.B1(n_13),
.B2(n_32),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_44),
.B1(n_26),
.B2(n_43),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_82),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_85),
.B1(n_88),
.B2(n_90),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_50),
.B1(n_37),
.B2(n_34),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_62),
.A2(n_51),
.B1(n_42),
.B2(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_87),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_41),
.B1(n_52),
.B2(n_34),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_71),
.Y(n_97)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_56),
.CI(n_60),
.CON(n_98),
.SN(n_98)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_102),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_109),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_95),
.Y(n_120)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_110),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_54),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_118),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_69),
.B(n_67),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_77),
.B(n_18),
.Y(n_139)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_124),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_86),
.B1(n_79),
.B2(n_91),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_126),
.B1(n_135),
.B2(n_125),
.Y(n_149)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_82),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_139),
.B(n_117),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_97),
.B1(n_63),
.B2(n_76),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_96),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_134),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_99),
.A2(n_76),
.B(n_83),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_65),
.B1(n_70),
.B2(n_77),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_102),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_49),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_98),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_108),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_100),
.B1(n_114),
.B2(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_135),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_157),
.Y(n_175)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_150),
.B(n_155),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_100),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_132),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_118),
.B1(n_112),
.B2(n_109),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_111),
.B(n_66),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_132),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_159),
.A2(n_66),
.B1(n_81),
.B2(n_128),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_120),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_156),
.B1(n_161),
.B2(n_144),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_153),
.A3(n_146),
.B1(n_142),
.B2(n_160),
.C1(n_147),
.C2(n_130),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_22),
.A3(n_25),
.B1(n_8),
.B2(n_9),
.C1(n_4),
.C2(n_6),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_164),
.B(n_162),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_124),
.C(n_140),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_171),
.C(n_22),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_121),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_156),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_185),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_49),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_186),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_115),
.B1(n_49),
.B2(n_37),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_172),
.B1(n_173),
.B2(n_2),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_25),
.B(n_22),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_49),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_189),
.C(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_22),
.C(n_25),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_185),
.A2(n_164),
.B1(n_177),
.B2(n_175),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_6),
.B(n_10),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_187),
.A2(n_166),
.B1(n_174),
.B2(n_8),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_192),
.A2(n_190),
.B(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_209),
.B(n_11),
.Y(n_217)
);

AO221x1_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_204)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_204),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_197),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_207),
.B(n_210),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_194),
.A2(n_8),
.B(n_11),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_199),
.B1(n_201),
.B2(n_196),
.Y(n_212)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_196),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_0),
.C(n_1),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_191),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_217),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_208),
.A3(n_203),
.B1(n_194),
.B2(n_11),
.C1(n_3),
.C2(n_2),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_0),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_0),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_218),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_213),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_224),
.B(n_225),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_211),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_219),
.B(n_2),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_228),
.C(n_1),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_3),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_3),
.Y(n_232)
);


endmodule