module fake_aes_1236_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
wire n_39;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_8), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
BUFx6f_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_2), .B(n_5), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_0), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_13), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
INVx5_ASAP7_75t_L g22 ( .A(n_14), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_19), .Y(n_23) );
AOI22xp5_ASAP7_75t_L g24 ( .A1(n_21), .A2(n_15), .B1(n_16), .B2(n_12), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_20), .B(n_0), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_22), .Y(n_26) );
NOR5xp2_ASAP7_75t_SL g27 ( .A(n_23), .B(n_1), .C(n_2), .D(n_22), .E(n_20), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_24), .Y(n_29) );
NAND2xp5_ASAP7_75t_L g30 ( .A(n_28), .B(n_26), .Y(n_30) );
INVx1_ASAP7_75t_SL g31 ( .A(n_29), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
AOI21xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_29), .B(n_22), .Y(n_34) );
BUFx3_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
AOI332xp33_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_27), .A3(n_22), .B1(n_18), .B2(n_10), .B3(n_7), .C1(n_4), .C2(n_11), .Y(n_36) );
BUFx6f_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
OAI21xp5_ASAP7_75t_L g38 ( .A1(n_34), .A2(n_18), .B(n_36), .Y(n_38) );
CKINVDCx20_ASAP7_75t_R g39 ( .A(n_37), .Y(n_39) );
NAND3xp33_ASAP7_75t_L g40 ( .A(n_39), .B(n_38), .C(n_37), .Y(n_40) );
endmodule