module fake_jpeg_19298_n_343 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_17),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_45),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_20),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_61),
.Y(n_75)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_63),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_39),
.C(n_48),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_34),
.B1(n_25),
.B2(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_67),
.Y(n_81)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_40),
.B1(n_34),
.B2(n_25),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_25),
.B1(n_70),
.B2(n_36),
.Y(n_118)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_73),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_24),
.B1(n_47),
.B2(n_38),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_107)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_89),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_80),
.B(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_85),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_38),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_88),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_93),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_71),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_101),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_47),
.B1(n_31),
.B2(n_36),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_66),
.A2(n_47),
.B1(n_28),
.B2(n_23),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_31),
.B1(n_36),
.B2(n_23),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_44),
.B(n_30),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_89),
.Y(n_119)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_79),
.B(n_69),
.CI(n_61),
.CON(n_108),
.SN(n_108)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_108),
.B(n_114),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_88),
.B1(n_100),
.B2(n_93),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

CKINVDCx6p67_ASAP7_75t_R g157 ( 
.A(n_110),
.Y(n_157)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_44),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_50),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_119),
.B(n_44),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_20),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_31),
.B1(n_23),
.B2(n_28),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_125),
.B1(n_128),
.B2(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_28),
.B1(n_22),
.B2(n_26),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_81),
.A2(n_26),
.B1(n_33),
.B2(n_43),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_81),
.A2(n_43),
.B1(n_41),
.B2(n_68),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_68),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_50),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_138),
.A2(n_153),
.B(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_76),
.Y(n_141)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_90),
.B1(n_82),
.B2(n_102),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_132),
.B1(n_104),
.B2(n_105),
.Y(n_181)
);

BUFx24_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_76),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_152),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_74),
.B1(n_43),
.B2(n_41),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_148),
.A2(n_106),
.B1(n_113),
.B2(n_112),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_74),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_73),
.B(n_1),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_41),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_155),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_117),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_109),
.A2(n_44),
.B(n_50),
.C(n_46),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_37),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_103),
.B(n_37),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_115),
.B(n_127),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_161),
.A2(n_168),
.B(n_32),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_162),
.A2(n_175),
.B1(n_182),
.B2(n_184),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_163),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_119),
.C(n_111),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_171),
.C(n_186),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_137),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_173),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_176),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_111),
.C(n_131),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_133),
.B1(n_132),
.B2(n_122),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_44),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_110),
.B1(n_123),
.B2(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_140),
.B1(n_157),
.B2(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_104),
.B1(n_105),
.B2(n_123),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_142),
.A2(n_130),
.B1(n_33),
.B2(n_37),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_84),
.C(n_46),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_162),
.B1(n_181),
.B2(n_166),
.Y(n_222)
);

AOI32xp33_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_149),
.A3(n_138),
.B1(n_143),
.B2(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_196),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_154),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_205),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_149),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_200),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_158),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_199),
.B(n_201),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_139),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_150),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_139),
.B1(n_150),
.B2(n_145),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_145),
.B1(n_157),
.B2(n_160),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_146),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_206),
.A2(n_218),
.B(n_32),
.Y(n_243)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_170),
.A2(n_164),
.A3(n_187),
.B1(n_176),
.B2(n_183),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_216),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_180),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_212),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_157),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_157),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_84),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_126),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_214),
.B(n_20),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_84),
.C(n_46),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_183),
.C(n_166),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_160),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_179),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_185),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_241),
.B1(n_217),
.B2(n_189),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_233),
.C(n_197),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_215),
.B(n_213),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_195),
.A2(n_21),
.B1(n_35),
.B2(n_19),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_234),
.B1(n_242),
.B2(n_208),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_195),
.A2(n_35),
.B1(n_21),
.B2(n_19),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_20),
.B(n_21),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_35),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_239),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_35),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_27),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_200),
.B(n_21),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_19),
.B1(n_18),
.B2(n_32),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_218),
.B(n_217),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_259),
.B1(n_265),
.B2(n_226),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_247),
.B(n_228),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_234),
.B1(n_232),
.B2(n_242),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_197),
.C(n_206),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_223),
.C(n_235),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_209),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_250),
.B(n_257),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_260),
.B(n_264),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_261),
.Y(n_278)
);

NAND3xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_207),
.C(n_204),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_204),
.B1(n_209),
.B2(n_196),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_227),
.B(n_209),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_18),
.B1(n_19),
.B2(n_2),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_263),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_0),
.B(n_1),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_8),
.B1(n_17),
.B2(n_3),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_SL g266 ( 
.A(n_245),
.B(n_8),
.C(n_13),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_236),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_249),
.B(n_233),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_271),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_226),
.B(n_223),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_267),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_280),
.B1(n_262),
.B2(n_251),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_256),
.B(n_235),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_237),
.B(n_8),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_231),
.Y(n_275)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_285),
.C(n_268),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_279),
.A2(n_246),
.B1(n_252),
.B2(n_251),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_220),
.B1(n_222),
.B2(n_229),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_253),
.A2(n_221),
.B(n_240),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_221),
.C(n_230),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_276),
.C(n_9),
.Y(n_312)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_290),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_264),
.B1(n_255),
.B2(n_254),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_263),
.C(n_260),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_300),
.C(n_0),
.Y(n_314)
);

NOR3xp33_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_263),
.C(n_239),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_279),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_7),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_298),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_281),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_27),
.C(n_7),
.Y(n_300)
);

AOI321xp33_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_7),
.A3(n_12),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_301),
.A2(n_278),
.B(n_272),
.Y(n_304)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_308),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_271),
.C(n_269),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_313),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_276),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_272),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_312),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_288),
.C(n_300),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_0),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_295),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_318),
.B(n_320),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_299),
.B1(n_293),
.B2(n_294),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_293),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_321),
.B(n_323),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_307),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_9),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_312),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_326),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_307),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_314),
.C(n_308),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_331),
.C(n_322),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_328),
.B(n_324),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_9),
.Y(n_331)
);

NAND2xp33_ASAP7_75t_SL g332 ( 
.A(n_329),
.B(n_316),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_332),
.A2(n_334),
.B(n_330),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_333),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_336),
.A2(n_335),
.B(n_328),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_337),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_6),
.B1(n_10),
.B2(n_11),
.Y(n_341)
);

O2A1O1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_10),
.B(n_13),
.C(n_1),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_13),
.Y(n_343)
);


endmodule