module fake_jpeg_2582_n_686 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_686);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_686;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_60),
.B(n_67),
.Y(n_135)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_63),
.Y(n_143)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_64),
.Y(n_171)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_65),
.Y(n_186)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_66),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g214 ( 
.A(n_70),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_20),
.B(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_72),
.B(n_78),
.Y(n_136)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_75),
.Y(n_193)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_76),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_32),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g162 ( 
.A(n_82),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_83),
.Y(n_212)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_104),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_40),
.B(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_86),
.B(n_88),
.Y(n_160)
);

BUFx16f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_0),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_42),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g140 ( 
.A(n_89),
.Y(n_140)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_91),
.Y(n_218)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_43),
.B(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_94),
.B(n_95),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_43),
.B(n_1),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_97),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_98),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_99),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_100),
.Y(n_229)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_101),
.Y(n_217)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_102),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_21),
.B(n_14),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_105),
.Y(n_232)
);

BUFx16f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_106),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_107),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_30),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_108),
.B(n_116),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_112),
.Y(n_219)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_35),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_36),
.Y(n_118)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_118),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_49),
.Y(n_119)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_122),
.B(n_54),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_39),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_124),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_126),
.Y(n_223)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_128),
.Y(n_228)
);

BUFx16f_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_44),
.Y(n_130)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_48),
.Y(n_132)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_146),
.B(n_179),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_70),
.A2(n_58),
.B1(n_22),
.B2(n_51),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_158),
.A2(n_178),
.B1(n_192),
.B2(n_54),
.Y(n_251)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_167),
.Y(n_260)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_172),
.Y(n_264)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_174),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_102),
.B(n_58),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_176),
.B(n_210),
.Y(n_235)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_71),
.Y(n_177)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_177),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_70),
.A2(n_58),
.B1(n_51),
.B2(n_54),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_129),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_88),
.B(n_48),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_183),
.B(n_201),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_87),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_184),
.B(n_199),
.Y(n_283)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_74),
.Y(n_185)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_185),
.Y(n_294)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_91),
.A2(n_53),
.B1(n_30),
.B2(n_56),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_190),
.A2(n_128),
.B1(n_126),
.B2(n_125),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_110),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_196),
.Y(n_295)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_197),
.Y(n_247)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_198),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_109),
.B(n_38),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_99),
.Y(n_200)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_123),
.B(n_38),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_100),
.Y(n_203)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_123),
.B(n_33),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_207),
.B(n_225),
.Y(n_248)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_105),
.Y(n_208)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_124),
.B(n_56),
.Y(n_210)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_115),
.A2(n_30),
.B1(n_53),
.B2(n_52),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_216),
.A2(n_178),
.B1(n_192),
.B2(n_158),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_106),
.A2(n_55),
.B(n_33),
.Y(n_222)
);

OR2x2_ASAP7_75t_SL g289 ( 
.A(n_222),
.B(n_77),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_96),
.B(n_25),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_119),
.Y(n_226)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_226),
.Y(n_316)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_79),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_127),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_111),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_142),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_233),
.Y(n_365)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_234),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_236),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_135),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_237),
.B(n_242),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_136),
.B(n_55),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_238),
.B(n_244),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_239),
.A2(n_297),
.B1(n_303),
.B2(n_314),
.Y(n_350)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_240),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_135),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_136),
.B(n_25),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_175),
.Y(n_245)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_245),
.Y(n_322)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_159),
.Y(n_249)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_148),
.B(n_23),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_250),
.B(n_273),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_251),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_150),
.B(n_23),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_252),
.B(n_254),
.Y(n_335)
);

INVx4_ASAP7_75t_SL g253 ( 
.A(n_140),
.Y(n_253)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_253),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_155),
.B(n_21),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_256),
.Y(n_347)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_257),
.Y(n_359)
);

BUFx8_ASAP7_75t_L g258 ( 
.A(n_182),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_258),
.Y(n_328)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_137),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_259),
.Y(n_360)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_145),
.Y(n_262)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_262),
.Y(n_380)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_141),
.Y(n_263)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_263),
.Y(n_381)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_180),
.Y(n_265)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_265),
.Y(n_324)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_145),
.Y(n_267)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_267),
.Y(n_351)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_269),
.Y(n_367)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_219),
.Y(n_271)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_271),
.Y(n_341)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_143),
.Y(n_272)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_163),
.B(n_160),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_163),
.B(n_53),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_274),
.B(n_276),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_182),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_161),
.B(n_165),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_277),
.B(n_288),
.Y(n_346)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_156),
.Y(n_278)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_278),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_160),
.B(n_54),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_298),
.Y(n_323)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_156),
.Y(n_280)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_280),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_281),
.A2(n_301),
.B1(n_315),
.B2(n_162),
.Y(n_330)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_285),
.Y(n_368)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_143),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_286),
.B(n_287),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_171),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_170),
.B(n_181),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_289),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_195),
.B(n_57),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_292),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_171),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_291),
.B(n_296),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_209),
.B(n_57),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_204),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_293),
.Y(n_379)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_144),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_222),
.A2(n_57),
.B1(n_131),
.B2(n_82),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_211),
.B(n_169),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_204),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_299),
.B(n_300),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_162),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_196),
.A2(n_225),
.B1(n_227),
.B2(n_194),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_133),
.B(n_1),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_309),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_139),
.A2(n_131),
.B1(n_82),
.B2(n_3),
.Y(n_303)
);

INVx3_ASAP7_75t_SL g304 ( 
.A(n_147),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_304),
.B(n_308),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_169),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_305),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g306 ( 
.A(n_134),
.B(n_103),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_157),
.C(n_202),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_199),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_307),
.A2(n_258),
.B(n_265),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_201),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_207),
.B(n_3),
.Y(n_309)
);

BUFx2_ASAP7_75t_SL g311 ( 
.A(n_153),
.Y(n_311)
);

INVx3_ASAP7_75t_SL g312 ( 
.A(n_206),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_217),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_224),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g315 ( 
.A1(n_153),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_193),
.B(n_7),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_317),
.B(n_318),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_138),
.B(n_10),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_149),
.B(n_14),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_319),
.B(n_10),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_330),
.A2(n_336),
.B1(n_352),
.B2(n_354),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_281),
.A2(n_205),
.B1(n_186),
.B2(n_168),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_334),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_301),
.A2(n_191),
.B1(n_154),
.B2(n_212),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_295),
.A2(n_205),
.B1(n_186),
.B2(n_213),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_337),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_279),
.B(n_151),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_338),
.B(n_356),
.C(n_366),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_339),
.B(n_345),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_235),
.A2(n_191),
.B1(n_229),
.B2(n_218),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_342),
.A2(n_294),
.B1(n_284),
.B2(n_275),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_295),
.A2(n_166),
.B1(n_228),
.B2(n_223),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

OA22x2_ASAP7_75t_L g345 ( 
.A1(n_251),
.A2(n_229),
.B1(n_221),
.B2(n_220),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_348),
.B(n_300),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_235),
.A2(n_221),
.B1(n_220),
.B2(n_218),
.Y(n_352)
);

OA21x2_ASAP7_75t_L g353 ( 
.A1(n_289),
.A2(n_214),
.B(n_154),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_353),
.B(n_371),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_239),
.A2(n_212),
.B1(n_214),
.B2(n_166),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_243),
.B(n_11),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_248),
.B(n_12),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_358),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_306),
.B(n_12),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_306),
.B(n_12),
.C(n_13),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_L g370 ( 
.A1(n_305),
.A2(n_14),
.B1(n_304),
.B2(n_312),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_370),
.A2(n_376),
.B1(n_315),
.B2(n_286),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_266),
.B(n_14),
.C(n_316),
.Y(n_371)
);

OA22x2_ASAP7_75t_L g374 ( 
.A1(n_313),
.A2(n_307),
.B1(n_287),
.B2(n_291),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

OAI22xp33_ASAP7_75t_L g376 ( 
.A1(n_262),
.A2(n_267),
.B1(n_285),
.B2(n_269),
.Y(n_376)
);

AOI21xp33_ASAP7_75t_L g397 ( 
.A1(n_377),
.A2(n_259),
.B(n_253),
.Y(n_397)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_382),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_353),
.A2(n_258),
.B(n_283),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_383),
.A2(n_397),
.B(n_377),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_384),
.A2(n_428),
.B1(n_351),
.B2(n_367),
.Y(n_450)
);

AND2x6_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_353),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_385),
.B(n_413),
.Y(n_460)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_386),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_338),
.B(n_264),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_388),
.B(n_400),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_321),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_389),
.B(n_391),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_330),
.A2(n_310),
.B1(n_270),
.B2(n_261),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_390),
.A2(n_402),
.B1(n_416),
.B2(n_343),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_333),
.B(n_255),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_321),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_393),
.B(n_394),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_355),
.B(n_326),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_332),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_396),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_296),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_398),
.B(n_407),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_349),
.B(n_260),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_362),
.A2(n_246),
.B1(n_282),
.B2(n_241),
.Y(n_402)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_403),
.Y(n_443)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

INVx13_ASAP7_75t_L g406 ( 
.A(n_328),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_406),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_346),
.B(n_271),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_408),
.B(n_421),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_327),
.B(n_234),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_410),
.B(n_412),
.Y(n_433)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_380),
.Y(n_411)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_411),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_272),
.Y(n_412)
);

INVx5_ASAP7_75t_L g413 ( 
.A(n_378),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_378),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_415),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_362),
.A2(n_260),
.B1(n_264),
.B2(n_294),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_417),
.B(n_418),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g418 ( 
.A(n_320),
.B(n_240),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_L g419 ( 
.A(n_325),
.B(n_278),
.C(n_247),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_419),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_350),
.A2(n_249),
.B1(n_256),
.B2(n_233),
.Y(n_422)
);

OAI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_422),
.A2(n_426),
.B1(n_331),
.B2(n_409),
.Y(n_445)
);

BUFx8_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_424),
.A2(n_366),
.B1(n_347),
.B2(n_324),
.Y(n_455)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_380),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_427),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_284),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_358),
.A2(n_275),
.B1(n_268),
.B2(n_257),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_369),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_431),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_340),
.B(n_268),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_423),
.A2(n_404),
.B1(n_414),
.B2(n_336),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_432),
.A2(n_435),
.B1(n_453),
.B2(n_456),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_323),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_434),
.B(n_436),
.C(n_444),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_423),
.A2(n_373),
.B1(n_352),
.B2(n_372),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_323),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_445),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_440),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_388),
.B(n_339),
.C(n_372),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_404),
.A2(n_372),
.B1(n_345),
.B2(n_370),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_446),
.A2(n_450),
.B1(n_451),
.B2(n_455),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_383),
.A2(n_369),
.B(n_374),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_449),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_399),
.A2(n_340),
.B1(n_325),
.B2(n_345),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_404),
.A2(n_345),
.B1(n_374),
.B2(n_348),
.Y(n_453)
);

OAI22x1_ASAP7_75t_L g456 ( 
.A1(n_414),
.A2(n_374),
.B1(n_233),
.B2(n_347),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_414),
.B(n_356),
.C(n_361),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_469),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_384),
.A2(n_351),
.B1(n_367),
.B2(n_368),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_463),
.B(n_473),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_390),
.A2(n_376),
.B1(n_329),
.B2(n_371),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_466),
.A2(n_405),
.B1(n_382),
.B2(n_386),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_387),
.B(n_341),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_387),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_364),
.C(n_324),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_418),
.A2(n_329),
.B1(n_359),
.B2(n_322),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_468),
.Y(n_474)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_474),
.Y(n_524)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_458),
.Y(n_475)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_441),
.B(n_410),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_476),
.B(n_495),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_477),
.B(n_467),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_433),
.B(n_400),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_478),
.B(n_487),
.Y(n_521)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_468),
.Y(n_479)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_479),
.Y(n_520)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_480),
.Y(n_526)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_464),
.Y(n_483)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_483),
.Y(n_528)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_485),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_433),
.B(n_447),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_473),
.Y(n_488)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_488),
.Y(n_537)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_438),
.Y(n_490)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_490),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_457),
.B(n_427),
.Y(n_491)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_491),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_492),
.A2(n_497),
.B1(n_501),
.B2(n_435),
.Y(n_530)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_461),
.Y(n_493)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_493),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_452),
.B(n_425),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_417),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_502),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_446),
.A2(n_395),
.B1(n_424),
.B2(n_408),
.Y(n_497)
);

INVx13_ASAP7_75t_L g498 ( 
.A(n_443),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_498),
.Y(n_522)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_438),
.Y(n_499)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_499),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_457),
.B(n_448),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_509),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_449),
.A2(n_395),
.B1(n_424),
.B2(n_420),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_436),
.B(n_413),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_504),
.Y(n_519)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_442),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_454),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_505),
.B(n_506),
.Y(n_525)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_454),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_453),
.B(n_424),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_508),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g509 ( 
.A(n_460),
.B(n_385),
.Y(n_509)
);

INVx13_ASAP7_75t_L g511 ( 
.A(n_443),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_511),
.B(n_512),
.Y(n_532)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_437),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_434),
.B(n_402),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_513),
.B(n_459),
.C(n_444),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_514),
.B(n_481),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_494),
.A2(n_462),
.B1(n_470),
.B2(n_466),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_515),
.A2(n_484),
.B1(n_488),
.B2(n_501),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_486),
.A2(n_440),
.B(n_465),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_518),
.A2(n_536),
.B(n_545),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_527),
.B(n_489),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_507),
.A2(n_456),
.B1(n_432),
.B2(n_470),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_529),
.A2(n_530),
.B1(n_546),
.B2(n_484),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_452),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_533),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_508),
.A2(n_465),
.B(n_469),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_500),
.B(n_448),
.Y(n_538)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_538),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_486),
.B(n_508),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_539),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_491),
.B(n_437),
.Y(n_542)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_542),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_482),
.B(n_463),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_543),
.B(n_544),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_482),
.B(n_439),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_507),
.A2(n_420),
.B(n_409),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_510),
.A2(n_416),
.B1(n_461),
.B2(n_472),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_492),
.B(n_472),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_547),
.B(n_497),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_494),
.A2(n_392),
.B(n_401),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_550),
.A2(n_484),
.B(n_511),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_477),
.B(n_359),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_551),
.B(n_396),
.Y(n_567)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_554),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_555),
.A2(n_570),
.B1(n_573),
.B2(n_546),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_542),
.B(n_493),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_556),
.B(n_557),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_532),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_558),
.B(n_571),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_561),
.A2(n_550),
.B1(n_543),
.B2(n_537),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_538),
.B(n_479),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_562),
.B(n_563),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_541),
.B(n_474),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_565),
.B(n_566),
.C(n_576),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_527),
.B(n_481),
.C(n_489),
.Y(n_566)
);

CKINVDCx14_ASAP7_75t_R g590 ( 
.A(n_567),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_568),
.A2(n_537),
.B1(n_526),
.B2(n_548),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_521),
.B(n_322),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g605 ( 
.A(n_569),
.B(n_575),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_515),
.A2(n_509),
.B1(n_396),
.B2(n_498),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_514),
.B(n_411),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_524),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g586 ( 
.A(n_572),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_544),
.A2(n_365),
.B1(n_406),
.B2(n_381),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_539),
.A2(n_403),
.B(n_247),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_574),
.A2(n_545),
.B(n_568),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_521),
.B(n_381),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_536),
.B(n_280),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_516),
.B(n_245),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_577),
.B(n_580),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_541),
.B(n_263),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_578),
.B(n_579),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_519),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_535),
.B(n_534),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_522),
.B(n_517),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_581),
.B(n_525),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_566),
.B(n_518),
.C(n_523),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_587),
.B(n_596),
.C(n_599),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_557),
.B(n_522),
.Y(n_591)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_591),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_592),
.A2(n_600),
.B1(n_607),
.B2(n_602),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_552),
.A2(n_560),
.B(n_539),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_593),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_555),
.A2(n_530),
.B1(n_534),
.B2(n_529),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_594),
.A2(n_582),
.B1(n_559),
.B2(n_576),
.Y(n_617)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_595),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_565),
.B(n_523),
.C(n_547),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_597),
.A2(n_607),
.B1(n_608),
.B2(n_552),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_558),
.B(n_517),
.C(n_526),
.Y(n_599)
);

OAI21xp33_ASAP7_75t_R g601 ( 
.A1(n_559),
.A2(n_549),
.B(n_540),
.Y(n_601)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_601),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_571),
.B(n_548),
.C(n_520),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_603),
.B(n_563),
.C(n_574),
.Y(n_620)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_604),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_562),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_606),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_570),
.A2(n_540),
.B1(n_549),
.B2(n_528),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_561),
.A2(n_528),
.B1(n_531),
.B2(n_520),
.Y(n_608)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_613),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_593),
.A2(n_560),
.B(n_554),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_615),
.B(n_626),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_591),
.B(n_556),
.Y(n_616)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_616),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_617),
.A2(n_618),
.B1(n_597),
.B2(n_595),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_592),
.A2(n_582),
.B1(n_553),
.B2(n_564),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_604),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_619),
.B(n_621),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_620),
.B(n_627),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_599),
.B(n_579),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_584),
.B(n_553),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_622),
.B(n_603),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_585),
.A2(n_573),
.B1(n_578),
.B2(n_531),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_624),
.A2(n_629),
.B1(n_590),
.B2(n_600),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_588),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_584),
.B(n_524),
.C(n_572),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_628),
.B(n_586),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_588),
.B(n_606),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_622),
.B(n_596),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_630),
.B(n_635),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_SL g631 ( 
.A(n_615),
.B(n_587),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_SL g656 ( 
.A(n_631),
.B(n_609),
.Y(n_656)
);

XOR2xp5_ASAP7_75t_L g635 ( 
.A(n_610),
.B(n_583),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_610),
.B(n_583),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g650 ( 
.A(n_636),
.B(n_643),
.Y(n_650)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_637),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_638),
.B(n_640),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_628),
.B(n_585),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_623),
.B(n_594),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_641),
.B(n_642),
.Y(n_659)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_626),
.B(n_608),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_620),
.B(n_602),
.C(n_589),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g651 ( 
.A(n_644),
.B(n_645),
.Y(n_651)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_618),
.B(n_598),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_SL g660 ( 
.A(n_646),
.B(n_616),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_630),
.B(n_625),
.C(n_617),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_648),
.B(n_652),
.C(n_653),
.Y(n_664)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_635),
.B(n_611),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_634),
.A2(n_614),
.B1(n_612),
.B2(n_632),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_SL g670 ( 
.A(n_656),
.B(n_648),
.Y(n_670)
);

OAI21xp33_ASAP7_75t_L g657 ( 
.A1(n_632),
.A2(n_625),
.B(n_609),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g667 ( 
.A1(n_657),
.A2(n_643),
.B(n_605),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_647),
.A2(n_623),
.B1(n_614),
.B2(n_629),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_661),
.C(n_605),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_660),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_636),
.B(n_589),
.C(n_598),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_655),
.B(n_644),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_662),
.B(n_663),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_651),
.B(n_633),
.Y(n_663)
);

AOI21x1_ASAP7_75t_SL g665 ( 
.A1(n_659),
.A2(n_631),
.B(n_639),
.Y(n_665)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_665),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_667),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_661),
.B(n_586),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_668),
.B(n_649),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_669),
.B(n_670),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_671),
.B(n_673),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_666),
.B(n_654),
.Y(n_673)
);

AOI21x1_ASAP7_75t_L g678 ( 
.A1(n_676),
.A2(n_666),
.B(n_664),
.Y(n_678)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_678),
.Y(n_681)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_672),
.B(n_649),
.C(n_670),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_679),
.B(n_674),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_680),
.B(n_677),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_682),
.B(n_676),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_SL g684 ( 
.A1(n_683),
.A2(n_681),
.B(n_675),
.Y(n_684)
);

XNOR2xp5_ASAP7_75t_L g685 ( 
.A(n_684),
.B(n_656),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_685),
.A2(n_657),
.B(n_650),
.Y(n_686)
);


endmodule