module fake_jpeg_2900_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_56),
.B(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_74),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_54),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_50),
.B1(n_46),
.B2(n_43),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_62),
.B1(n_59),
.B2(n_54),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_51),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_70),
.B1(n_62),
.B2(n_59),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_43),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_42),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_105),
.B1(n_55),
.B2(n_63),
.Y(n_108)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_0),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_83),
.B1(n_81),
.B2(n_85),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_47),
.B1(n_14),
.B2(n_19),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_2),
.B(n_3),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_64),
.B1(n_55),
.B2(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_76),
.B(n_0),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_1),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_114),
.B1(n_123),
.B2(n_5),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_17),
.C(n_39),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_113),
.C(n_95),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_115),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_15),
.C(n_37),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_1),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_13),
.B1(n_32),
.B2(n_30),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_120),
.B(n_21),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_121),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_12),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_127),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_95),
.C(n_22),
.Y(n_128)
);

XOR2x2_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_138),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_137),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_133),
.B(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_6),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_7),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_24),
.B(n_29),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_113),
.CI(n_23),
.CON(n_142),
.SN(n_142)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_134),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_140)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_126),
.C(n_128),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_143),
.B(n_135),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_149),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_133),
.B1(n_125),
.B2(n_130),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_151),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_129),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_150),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_153),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_152),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_145),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_146),
.B1(n_142),
.B2(n_140),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_26),
.B(n_27),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_36),
.Y(n_162)
);


endmodule