module fake_jpeg_6848_n_345 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_47),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_41),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_29),
.Y(n_53)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_53),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_21),
.B1(n_33),
.B2(n_31),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_27),
.B1(n_34),
.B2(n_25),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_63),
.B1(n_72),
.B2(n_27),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_34),
.B1(n_20),
.B2(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_26),
.C(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_32),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_27),
.B1(n_34),
.B2(n_18),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_81),
.B1(n_21),
.B2(n_17),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_87),
.B1(n_66),
.B2(n_23),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_26),
.B1(n_33),
.B2(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_38),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_91),
.Y(n_103)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_92),
.Y(n_106)
);

AND2x4_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_29),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_99),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_18),
.B1(n_17),
.B2(n_23),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_28),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_75),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_51),
.B(n_39),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_17),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_101),
.Y(n_142)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_108),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_39),
.C(n_36),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_110),
.C(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_56),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_78),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_109),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_50),
.A3(n_66),
.B1(n_58),
.B2(n_48),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_28),
.Y(n_111)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_21),
.B1(n_23),
.B2(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_28),
.Y(n_118)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_94),
.Y(n_120)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_130),
.B1(n_86),
.B2(n_92),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_65),
.C(n_67),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_58),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_32),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_88),
.A2(n_69),
.B1(n_60),
.B2(n_71),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_132),
.A2(n_133),
.B1(n_147),
.B2(n_149),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_94),
.B1(n_70),
.B2(n_77),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_145),
.B1(n_151),
.B2(n_156),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_22),
.C(n_32),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_155),
.Y(n_159)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_148),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_73),
.B1(n_76),
.B2(n_82),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_89),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_115),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_77),
.B1(n_76),
.B2(n_97),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_74),
.B(n_77),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_105),
.B1(n_127),
.B2(n_103),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_32),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_154),
.A2(n_118),
.B(n_111),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_106),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_93),
.B1(n_82),
.B2(n_74),
.Y(n_156)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_160),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_149),
.A2(n_110),
.B1(n_113),
.B2(n_104),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_120),
.B(n_109),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_161),
.A2(n_166),
.B(n_174),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_171),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_164),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_107),
.B1(n_102),
.B2(n_124),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_167),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_116),
.B(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_173),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_114),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_107),
.C(n_122),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_172),
.B(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_131),
.B(n_108),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_178),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_137),
.A2(n_119),
.B(n_93),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_177),
.B(n_179),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_32),
.B(n_22),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_24),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_180),
.C(n_183),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_126),
.C(n_64),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_24),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_182),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_24),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_112),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_147),
.B1(n_136),
.B2(n_153),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_186),
.A2(n_207),
.B1(n_210),
.B2(n_22),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_196),
.C(n_183),
.Y(n_213)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_200),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_131),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_166),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_175),
.B(n_169),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_199),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_171),
.B(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_184),
.A2(n_142),
.B1(n_152),
.B2(n_139),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_197),
.A2(n_206),
.B1(n_212),
.B2(n_198),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_150),
.B(n_142),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_209),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_150),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_211),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_154),
.B1(n_139),
.B2(n_149),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_167),
.A2(n_132),
.B1(n_148),
.B2(n_155),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_164),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_177),
.A2(n_154),
.B1(n_140),
.B2(n_135),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_168),
.A2(n_22),
.B1(n_64),
.B2(n_32),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_214),
.C(n_225),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_176),
.C(n_172),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_181),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_226),
.B(n_192),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_180),
.B1(n_182),
.B2(n_161),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_231),
.B1(n_234),
.B2(n_212),
.Y(n_241)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_223),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_237),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_174),
.C(n_170),
.Y(n_225)
);

A2O1A1O1Ixp25_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_112),
.B(n_22),
.C(n_19),
.D(n_24),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_210),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_158),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_95),
.C(n_24),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_233),
.C(n_29),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_195),
.Y(n_230)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_235),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_95),
.C(n_24),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_95),
.B1(n_22),
.B2(n_24),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_19),
.B(n_24),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_236),
.A2(n_200),
.B(n_190),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_186),
.A2(n_19),
.B1(n_29),
.B2(n_2),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_215),
.B(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_218),
.B(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_187),
.B1(n_212),
.B2(n_199),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_246),
.A2(n_260),
.B1(n_19),
.B2(n_1),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_0),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_238),
.A2(n_206),
.B(n_204),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_237),
.Y(n_262)
);

NAND2x1p5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_197),
.Y(n_250)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_227),
.B1(n_19),
.B2(n_2),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_201),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_255),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_225),
.A2(n_192),
.B(n_193),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_257),
.C(n_261),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_19),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_229),
.C(n_228),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_216),
.B1(n_226),
.B2(n_224),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_29),
.C(n_19),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_264),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_273),
.B1(n_281),
.B2(n_259),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_252),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_269),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_9),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_274),
.C(n_278),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_241),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_1),
.C(n_4),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_278),
.C(n_261),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_256),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_244),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_250),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_1),
.C(n_5),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_247),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_285),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_248),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_255),
.C(n_250),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_290),
.C(n_265),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_297),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_265),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_258),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_262),
.B(n_293),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_243),
.C(n_254),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_249),
.B1(n_246),
.B2(n_6),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_277),
.B1(n_8),
.B2(n_9),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_11),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_12),
.Y(n_312)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_298),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_266),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_12),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_292),
.B(n_263),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_300),
.A2(n_306),
.B(n_308),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_305),
.C(n_307),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_281),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_280),
.C(n_264),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_273),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_277),
.B(n_8),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_8),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_311),
.B(n_312),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_282),
.Y(n_314)
);

AOI31xp33_ASAP7_75t_L g329 ( 
.A1(n_314),
.A2(n_13),
.A3(n_15),
.B(n_16),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_286),
.Y(n_315)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_318),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_318),
.B(n_13),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_301),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_10),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_307),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_11),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_321),
.B(n_317),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_325),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_330),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_310),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_328),
.C(n_329),
.Y(n_338)
);

AOI21x1_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_305),
.B(n_11),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_322),
.C(n_323),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_335),
.C(n_15),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_331),
.B(n_313),
.C(n_13),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_SL g336 ( 
.A(n_332),
.B(n_15),
.Y(n_336)
);

OAI21xp33_ASAP7_75t_SL g340 ( 
.A1(n_336),
.A2(n_16),
.B(n_6),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_339),
.B(n_340),
.C(n_338),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_333),
.B(n_337),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_342),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_16),
.Y(n_344)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_344),
.Y(n_345)
);


endmodule