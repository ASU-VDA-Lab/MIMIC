module fake_jpeg_11696_n_181 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_36),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_26),
.Y(n_68)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_11),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_17),
.A2(n_1),
.B1(n_3),
.B2(n_7),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_42),
.B(n_43),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_3),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_7),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_61),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_14),
.B(n_9),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_22),
.A2(n_7),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_49),
.B(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx5_ASAP7_75t_SL g51 ( 
.A(n_23),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_18),
.A2(n_9),
.B1(n_19),
.B2(n_24),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_31),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_26),
.B1(n_27),
.B2(n_19),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_51),
.B1(n_59),
.B2(n_52),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_45),
.Y(n_67)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_46),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_89),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_29),
.B1(n_31),
.B2(n_27),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_88),
.B1(n_84),
.B2(n_91),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_83),
.A2(n_84),
.B1(n_70),
.B2(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_38),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

CKINVDCx10_ASAP7_75t_R g101 ( 
.A(n_67),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_50),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_108),
.B(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_33),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_113),
.Y(n_132)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_82),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_39),
.B1(n_96),
.B2(n_82),
.Y(n_113)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_78),
.B1(n_71),
.B2(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_75),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_119),
.B(n_120),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_71),
.A2(n_86),
.B1(n_92),
.B2(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_119),
.B1(n_118),
.B2(n_116),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_66),
.B(n_91),
.C(n_94),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_135),
.B(n_99),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_129),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_79),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_77),
.B(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_132),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_143),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_109),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_142),
.C(n_137),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_112),
.C(n_105),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_113),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_126),
.B1(n_124),
.B2(n_133),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_147),
.B(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_121),
.A2(n_103),
.B1(n_115),
.B2(n_100),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_155),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_133),
.B(n_99),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_135),
.C(n_124),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_130),
.C(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

AO21x2_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_145),
.B(n_143),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_159),
.B1(n_163),
.B2(n_155),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_151),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_107),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_144),
.B1(n_142),
.B2(n_147),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_130),
.C(n_128),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_157),
.A2(n_153),
.B1(n_150),
.B2(n_148),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_120),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_161),
.B1(n_110),
.B2(n_128),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_152),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_166),
.B(n_167),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_168),
.A2(n_114),
.B(n_102),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_171),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_172),
.A2(n_166),
.B(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_86),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_168),
.C(n_102),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_102),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_178),
.A2(n_175),
.B(n_76),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_179),
.Y(n_181)
);


endmodule