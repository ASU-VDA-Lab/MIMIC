module fake_aes_8194_n_753 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_753);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_753;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_725;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_40), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_18), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_47), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_55), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_71), .Y(n_86) );
INVx1_ASAP7_75t_SL g87 ( .A(n_9), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_80), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_5), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_43), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_33), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_68), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_11), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_11), .Y(n_94) );
INVxp67_ASAP7_75t_SL g95 ( .A(n_81), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_65), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_16), .Y(n_97) );
XOR2x2_ASAP7_75t_L g98 ( .A(n_9), .B(n_30), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_73), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_2), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_34), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_37), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_17), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_56), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_78), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_72), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_75), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_79), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_27), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_28), .Y(n_111) );
NOR2xp67_ASAP7_75t_L g112 ( .A(n_31), .B(n_48), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_64), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_25), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_35), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_46), .Y(n_116) );
NOR2xp67_ASAP7_75t_L g117 ( .A(n_53), .B(n_6), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_32), .Y(n_118) );
CKINVDCx14_ASAP7_75t_R g119 ( .A(n_39), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_5), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_4), .Y(n_121) );
CKINVDCx14_ASAP7_75t_R g122 ( .A(n_29), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_63), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_54), .Y(n_124) );
INVxp33_ASAP7_75t_L g125 ( .A(n_57), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_10), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_10), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_76), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_19), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_36), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_67), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_105), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_94), .B(n_0), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_97), .B(n_0), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_125), .B(n_1), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_93), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_94), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_108), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_93), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_125), .B(n_100), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_121), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_108), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_119), .B(n_1), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_100), .B(n_2), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_89), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_119), .B(n_3), .Y(n_147) );
XNOR2xp5_ASAP7_75t_L g148 ( .A(n_98), .B(n_3), .Y(n_148) );
NOR2xp33_ASAP7_75t_SL g149 ( .A(n_115), .B(n_42), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
INVxp67_ASAP7_75t_L g151 ( .A(n_103), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_120), .B(n_4), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_108), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_82), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_82), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_114), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_86), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_122), .B(n_6), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_85), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_121), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_83), .B(n_44), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_88), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_83), .B(n_7), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_90), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_91), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_126), .B(n_7), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_92), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_99), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_122), .B(n_8), .Y(n_170) );
OAI22x1_ASAP7_75t_L g171 ( .A1(n_98), .A2(n_8), .B1(n_12), .B2(n_13), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_127), .B(n_12), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_102), .Y(n_173) );
INVxp67_ASAP7_75t_L g174 ( .A(n_87), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_117), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_104), .B(n_13), .Y(n_176) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_174), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_158), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_143), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_141), .B(n_131), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_162), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_162), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_160), .B(n_131), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_137), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_151), .B(n_84), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_133), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_146), .B(n_84), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_133), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_133), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_155), .B(n_101), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_160), .B(n_101), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_154), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_164), .B(n_130), .Y(n_200) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_140), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_163), .B(n_96), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_162), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_167), .A2(n_114), .B1(n_118), .B2(n_95), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_135), .B(n_14), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_144), .B(n_107), .Y(n_206) );
OAI221xp5_ASAP7_75t_L g207 ( .A1(n_155), .A2(n_129), .B1(n_128), .B2(n_124), .C(n_123), .Y(n_207) );
AND2x6_ASAP7_75t_L g208 ( .A(n_164), .B(n_111), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_133), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_134), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_163), .B(n_116), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_150), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_134), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_166), .B(n_113), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
OR2x6_ASAP7_75t_L g216 ( .A(n_171), .B(n_118), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_156), .B(n_110), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_132), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_134), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_166), .B(n_109), .Y(n_222) );
NOR2xp33_ASAP7_75t_SL g223 ( .A(n_149), .B(n_112), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_164), .Y(n_224) );
BUFx10_ASAP7_75t_L g225 ( .A(n_164), .Y(n_225) );
NAND2xp33_ASAP7_75t_L g226 ( .A(n_162), .B(n_106), .Y(n_226) );
AO22x2_ASAP7_75t_L g227 ( .A1(n_167), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_156), .Y(n_229) );
INVxp67_ASAP7_75t_SL g230 ( .A(n_144), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_147), .B(n_159), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_167), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_165), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
INVxp67_ASAP7_75t_SL g236 ( .A(n_159), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_170), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_170), .B(n_15), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_165), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_138), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_168), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_168), .B(n_51), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_168), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_169), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_169), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_181), .B(n_186), .Y(n_246) );
NOR2x1_ASAP7_75t_L g247 ( .A(n_189), .B(n_145), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_177), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_240), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_180), .B(n_136), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_225), .Y(n_251) );
INVx3_ASAP7_75t_L g252 ( .A(n_225), .Y(n_252) );
BUFx8_ASAP7_75t_L g253 ( .A(n_191), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_185), .B(n_172), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_197), .B(n_172), .Y(n_255) );
NAND3xp33_ASAP7_75t_SL g256 ( .A(n_219), .B(n_157), .C(n_142), .Y(n_256) );
NOR2x1p5_ASAP7_75t_L g257 ( .A(n_191), .B(n_148), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_208), .A2(n_173), .B1(n_169), .B2(n_162), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_240), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_234), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_204), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_233), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_230), .B(n_236), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_182), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_234), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_237), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_225), .Y(n_267) );
OR2x6_ASAP7_75t_L g268 ( .A(n_216), .B(n_171), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_235), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_190), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_240), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_182), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_196), .B(n_152), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_212), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_226), .A2(n_173), .B(n_175), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_238), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_235), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_188), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_202), .B(n_173), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_179), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_179), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_239), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_206), .B(n_138), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_201), .B(n_148), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_239), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_241), .Y(n_286) );
INVx5_ASAP7_75t_L g287 ( .A(n_208), .Y(n_287) );
NOR2xp33_ASAP7_75t_R g288 ( .A(n_226), .B(n_161), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_212), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_241), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_206), .B(n_138), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_229), .B(n_138), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_181), .B(n_176), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_243), .Y(n_294) );
AND2x6_ASAP7_75t_SL g295 ( .A(n_216), .B(n_17), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_190), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_231), .A2(n_153), .B1(n_139), .B2(n_134), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_203), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_229), .B(n_153), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_200), .B(n_153), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_181), .B(n_139), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_200), .B(n_153), .Y(n_302) );
INVxp67_ASAP7_75t_L g303 ( .A(n_204), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_186), .B(n_139), .Y(n_304) );
OR2x2_ASAP7_75t_SL g305 ( .A(n_216), .B(n_139), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_193), .A2(n_153), .B(n_139), .C(n_22), .Y(n_306) );
INVx2_ASAP7_75t_SL g307 ( .A(n_200), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_205), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_190), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_193), .B(n_20), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_208), .B(n_21), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_194), .B(n_23), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_243), .Y(n_313) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_186), .B(n_24), .Y(n_314) );
NOR2x1p5_ASAP7_75t_L g315 ( .A(n_205), .B(n_26), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_216), .B(n_38), .Y(n_316) );
NOR3xp33_ASAP7_75t_SL g317 ( .A(n_207), .B(n_45), .C(n_49), .Y(n_317) );
INVx2_ASAP7_75t_SL g318 ( .A(n_238), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_211), .B(n_50), .Y(n_319) );
INVx5_ASAP7_75t_L g320 ( .A(n_287), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_251), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_270), .Y(n_322) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_279), .A2(n_228), .B(n_232), .C(n_224), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_279), .A2(n_228), .B(n_232), .C(n_224), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_251), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_252), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_276), .A2(n_194), .B1(n_209), .B2(n_228), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_248), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_301), .A2(n_203), .B(n_220), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_270), .Y(n_330) );
OR2x6_ASAP7_75t_L g331 ( .A(n_268), .B(n_227), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_248), .B(n_227), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_308), .B(n_208), .Y(n_333) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_273), .A2(n_209), .B(n_222), .C(n_245), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_296), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_276), .A2(n_209), .B1(n_227), .B2(n_245), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_287), .B(n_220), .Y(n_337) );
INVx2_ASAP7_75t_SL g338 ( .A(n_253), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_253), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_283), .A2(n_214), .B(n_244), .C(n_178), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_296), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_309), .Y(n_342) );
NAND2xp33_ASAP7_75t_L g343 ( .A(n_287), .B(n_208), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_278), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_266), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_266), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_303), .A2(n_227), .B1(n_244), .B2(n_215), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_252), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_256), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_262), .B(n_215), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_309), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_274), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_267), .Y(n_353) );
AND3x1_ASAP7_75t_SL g354 ( .A(n_257), .B(n_223), .C(n_184), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_287), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_305), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_292), .Y(n_357) );
OAI21x1_ASAP7_75t_L g358 ( .A1(n_301), .A2(n_242), .B(n_218), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_264), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_304), .A2(n_178), .B(n_184), .Y(n_360) );
OR2x6_ASAP7_75t_L g361 ( .A(n_268), .B(n_187), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_291), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_288), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_316), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_288), .Y(n_365) );
OAI22xp5_ASAP7_75t_SL g366 ( .A1(n_268), .A2(n_187), .B1(n_208), .B2(n_199), .Y(n_366) );
BUFx12f_ASAP7_75t_L g367 ( .A(n_295), .Y(n_367) );
OR2x6_ASAP7_75t_L g368 ( .A(n_307), .B(n_208), .Y(n_368) );
BUFx8_ASAP7_75t_L g369 ( .A(n_284), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_263), .B(n_52), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_260), .Y(n_371) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_254), .A2(n_199), .B(n_198), .C(n_195), .Y(n_372) );
INVx6_ASAP7_75t_L g373 ( .A(n_315), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_264), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_265), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_261), .A2(n_198), .B1(n_192), .B2(n_195), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_320), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_361), .B(n_267), .Y(n_378) );
AO21x2_ASAP7_75t_L g379 ( .A1(n_336), .A2(n_306), .B(n_317), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_328), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_361), .B(n_318), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_345), .B(n_346), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_372), .A2(n_304), .B(n_275), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_352), .Y(n_384) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_347), .B(n_317), .C(n_306), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_344), .B(n_258), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_371), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_336), .A2(n_314), .B(n_311), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_331), .A2(n_258), .B1(n_313), .B2(n_286), .Y(n_389) );
AO21x2_ASAP7_75t_L g390 ( .A1(n_347), .A2(n_314), .B(n_312), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_320), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_375), .Y(n_392) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_339), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_334), .A2(n_255), .B(n_250), .C(n_293), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_357), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_362), .A2(n_250), .B1(n_273), .B2(n_282), .C(n_269), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_327), .A2(n_294), .B1(n_285), .B2(n_290), .C(n_277), .Y(n_397) );
OAI21x1_ASAP7_75t_L g398 ( .A1(n_372), .A2(n_299), .B(n_312), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_358), .A2(n_310), .B(n_319), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_345), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_346), .Y(n_401) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_343), .B(n_310), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_331), .A2(n_289), .B1(n_297), .B2(n_302), .Y(n_403) );
OAI21x1_ASAP7_75t_L g404 ( .A1(n_340), .A2(n_300), .B(n_246), .Y(n_404) );
AO21x2_ASAP7_75t_L g405 ( .A1(n_323), .A2(n_293), .B(n_259), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_350), .B(n_247), .Y(n_406) );
OAI21x1_ASAP7_75t_SL g407 ( .A1(n_340), .A2(n_249), .B(n_271), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_359), .Y(n_408) );
OAI21x1_ASAP7_75t_L g409 ( .A1(n_360), .A2(n_246), .B(n_281), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_361), .B(n_298), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_327), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_396), .A2(n_332), .B1(n_349), .B2(n_338), .C(n_324), .Y(n_412) );
O2A1O1Ixp33_ASAP7_75t_L g413 ( .A1(n_400), .A2(n_331), .B(n_333), .C(n_364), .Y(n_413) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_377), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_402), .A2(n_370), .B(n_368), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g416 ( .A1(n_394), .A2(n_333), .B(n_376), .C(n_353), .Y(n_416) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_396), .A2(n_353), .B(n_360), .C(n_326), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_395), .A2(n_397), .B1(n_411), .B2(n_380), .C(n_387), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_395), .B(n_322), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_402), .A2(n_368), .B(n_329), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_384), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_389), .A2(n_373), .B1(n_363), .B2(n_366), .Y(n_422) );
AOI211xp5_ASAP7_75t_L g423 ( .A1(n_389), .A2(n_356), .B(n_365), .C(n_354), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_384), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_387), .B(n_368), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_382), .B(n_369), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_397), .A2(n_373), .B1(n_321), .B2(n_325), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_411), .A2(n_373), .B1(n_367), .B2(n_369), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_385), .A2(n_321), .B1(n_325), .B2(n_348), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_402), .A2(n_329), .B(n_341), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_377), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
OA21x2_ASAP7_75t_L g434 ( .A1(n_398), .A2(n_351), .B(n_342), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_409), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_409), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_392), .Y(n_437) );
OAI21x1_ASAP7_75t_L g438 ( .A1(n_399), .A2(n_326), .B(n_348), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_377), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_401), .Y(n_440) );
NAND2x1_ASAP7_75t_L g441 ( .A(n_407), .B(n_374), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_412), .A2(n_381), .B1(n_385), .B2(n_406), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_437), .B(n_392), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_437), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_435), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g447 ( .A1(n_422), .A2(n_406), .B1(n_403), .B2(n_386), .C(n_383), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_421), .Y(n_448) );
OR2x6_ASAP7_75t_L g449 ( .A(n_415), .B(n_407), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_418), .B(n_390), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_435), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_433), .B(n_405), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_441), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_433), .B(n_405), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_436), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_414), .Y(n_456) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_436), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_440), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_421), .Y(n_459) );
INVxp67_ASAP7_75t_SL g460 ( .A(n_424), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_424), .B(n_381), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_431), .B(n_390), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_431), .B(n_390), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_434), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_441), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_439), .B(n_381), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_419), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_434), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_414), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_434), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_419), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_438), .Y(n_473) );
AOI21x1_ASAP7_75t_L g474 ( .A1(n_430), .A2(n_398), .B(n_388), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_426), .B(n_393), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_438), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_414), .B(n_381), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_444), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_444), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_469), .B(n_432), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_477), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_458), .Y(n_483) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_450), .A2(n_399), .B(n_388), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_460), .B(n_425), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_464), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_467), .B(n_423), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_442), .B(n_423), .C(n_428), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_460), .B(n_425), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_469), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_464), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_477), .Y(n_492) );
AOI322xp5_ASAP7_75t_L g493 ( .A1(n_467), .A2(n_439), .A3(n_378), .B1(n_417), .B2(n_416), .C1(n_432), .C2(n_410), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_448), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_448), .B(n_432), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_459), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_452), .B(n_427), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_459), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_464), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_447), .A2(n_427), .B(n_429), .Y(n_500) );
INVx2_ASAP7_75t_SL g501 ( .A(n_469), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_468), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_468), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_452), .B(n_390), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_468), .Y(n_505) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_450), .A2(n_399), .B(n_388), .Y(n_506) );
BUFx2_ASAP7_75t_SL g507 ( .A(n_446), .Y(n_507) );
AOI21xp33_ASAP7_75t_L g508 ( .A1(n_447), .A2(n_413), .B(n_429), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_475), .B(n_403), .C(n_378), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_454), .B(n_405), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_465), .B(n_420), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_454), .B(n_405), .Y(n_512) );
AOI31xp33_ASAP7_75t_L g513 ( .A1(n_472), .A2(n_378), .A3(n_410), .B(n_383), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_472), .B(n_379), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_453), .B(n_391), .C(n_410), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_461), .B(n_379), .Y(n_516) );
INVx1_ASAP7_75t_SL g517 ( .A(n_461), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_466), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_471), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_471), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_466), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_465), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_471), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_443), .B(n_379), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_443), .B(n_379), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_465), .B(n_449), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_478), .B(n_378), .Y(n_527) );
OAI33xp33_ASAP7_75t_L g528 ( .A1(n_462), .A2(n_330), .A3(n_192), .B1(n_183), .B2(n_210), .B3(n_221), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_446), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_446), .B(n_408), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_462), .B(n_410), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_488), .A2(n_449), .B1(n_453), .B2(n_463), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_510), .B(n_463), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_510), .B(n_455), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_512), .B(n_455), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_483), .B(n_446), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_512), .B(n_451), .Y(n_538) );
OAI31xp33_ASAP7_75t_L g539 ( .A1(n_509), .A2(n_476), .A3(n_473), .B(n_391), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_479), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_480), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_526), .B(n_465), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_480), .Y(n_543) );
AOI31xp33_ASAP7_75t_L g544 ( .A1(n_500), .A2(n_476), .A3(n_473), .B(n_457), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_531), .B(n_451), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_490), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_495), .Y(n_547) );
AND2x4_ASAP7_75t_SL g548 ( .A(n_481), .B(n_456), .Y(n_548) );
NAND4xp25_ASAP7_75t_L g549 ( .A(n_487), .B(n_470), .C(n_456), .D(n_391), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_518), .B(n_456), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_516), .B(n_455), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_497), .B(n_445), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_482), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_497), .B(n_445), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_482), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_492), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_516), .B(n_451), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_504), .B(n_445), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_521), .B(n_456), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_526), .B(n_511), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_494), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_517), .B(n_470), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_504), .B(n_457), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_525), .B(n_449), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_486), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_508), .A2(n_449), .B1(n_470), .B2(n_465), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_495), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_514), .B(n_449), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_490), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_525), .B(n_474), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_494), .B(n_470), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_496), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_507), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_496), .B(n_465), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_498), .B(n_474), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_492), .B(n_404), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_486), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_514), .B(n_404), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_498), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_485), .B(n_404), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_485), .B(n_391), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_489), .B(n_408), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_489), .A2(n_408), .B1(n_335), .B2(n_359), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_524), .B(n_183), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_491), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_502), .B(n_374), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_529), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_502), .B(n_505), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_505), .B(n_58), .Y(n_589) );
NOR2x1_ASAP7_75t_SL g590 ( .A(n_515), .B(n_320), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_519), .B(n_59), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_519), .B(n_60), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_520), .B(n_61), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_532), .B(n_493), .C(n_513), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_587), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_553), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_546), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_544), .B(n_526), .Y(n_598) );
NAND2x1p5_ASAP7_75t_L g599 ( .A(n_589), .B(n_481), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_533), .B(n_526), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_547), .B(n_520), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_533), .B(n_491), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_569), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_553), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_555), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_558), .B(n_503), .Y(n_606) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_588), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_555), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_589), .B(n_481), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_567), .B(n_499), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_545), .B(n_499), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_573), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_558), .B(n_523), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_534), .B(n_523), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_537), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_545), .B(n_503), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_556), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_556), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_535), .B(n_501), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_549), .B(n_527), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_540), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_534), .B(n_511), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_539), .B(n_511), .C(n_530), .D(n_210), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_565), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_548), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_536), .B(n_511), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_577), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_536), .B(n_538), .Y(n_629) );
INVx2_ASAP7_75t_SL g630 ( .A(n_548), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_538), .B(n_506), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_591), .B(n_501), .Y(n_632) );
NAND2x1_ASAP7_75t_L g633 ( .A(n_561), .B(n_522), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_563), .B(n_507), .Y(n_634) );
NOR2xp67_ASAP7_75t_SL g635 ( .A(n_591), .B(n_522), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_564), .B(n_530), .Y(n_636) );
INVx3_ASAP7_75t_L g637 ( .A(n_560), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_541), .Y(n_638) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_563), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_564), .B(n_528), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_543), .B(n_522), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_572), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_579), .Y(n_643) );
XNOR2x2_ASAP7_75t_L g644 ( .A(n_550), .B(n_506), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_570), .A2(n_522), .B(n_221), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_571), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_551), .B(n_506), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_559), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_574), .Y(n_649) );
NOR4xp25_ASAP7_75t_L g650 ( .A(n_612), .B(n_566), .C(n_581), .D(n_562), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_629), .B(n_560), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_607), .B(n_570), .Y(n_652) );
AOI222xp33_ASAP7_75t_SL g653 ( .A1(n_597), .A2(n_577), .B1(n_585), .B2(n_568), .C1(n_580), .C2(n_560), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_646), .B(n_551), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_639), .B(n_552), .Y(n_655) );
NOR4xp25_ASAP7_75t_SL g656 ( .A(n_598), .B(n_590), .C(n_592), .D(n_593), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_640), .A2(n_576), .B1(n_557), .B2(n_575), .C(n_568), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_594), .A2(n_580), .B1(n_582), .B2(n_578), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_595), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_601), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_606), .Y(n_661) );
OAI21xp33_ASAP7_75t_L g662 ( .A1(n_640), .A2(n_576), .B(n_557), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_621), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_603), .B(n_578), .C(n_583), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_606), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_629), .Y(n_666) );
OAI32xp33_ASAP7_75t_L g667 ( .A1(n_598), .A2(n_552), .A3(n_554), .B1(n_593), .B2(n_592), .Y(n_667) );
INVx1_ASAP7_75t_SL g668 ( .A(n_611), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_616), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_623), .A2(n_599), .B1(n_609), .B2(n_632), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_648), .B(n_554), .Y(n_671) );
INVxp67_ASAP7_75t_L g672 ( .A(n_620), .Y(n_672) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_632), .A2(n_542), .B(n_582), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_638), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_642), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_643), .Y(n_676) );
OAI322xp33_ASAP7_75t_L g677 ( .A1(n_644), .A2(n_584), .A3(n_585), .B1(n_586), .B2(n_522), .C1(n_590), .C2(n_506), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_631), .B(n_542), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_620), .B(n_542), .C(n_484), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_596), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_625), .A2(n_484), .B1(n_374), .B2(n_359), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g682 ( .A1(n_599), .A2(n_484), .B1(n_355), .B2(n_320), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_604), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_625), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_605), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_637), .A2(n_484), .B1(n_217), .B2(n_213), .Y(n_686) );
INVxp67_ASAP7_75t_L g687 ( .A(n_615), .Y(n_687) );
INVx1_ASAP7_75t_SL g688 ( .A(n_630), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_660), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_672), .A2(n_644), .B1(n_600), .B2(n_637), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_672), .B(n_619), .C(n_645), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_660), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_652), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_663), .Y(n_694) );
OAI21x1_ASAP7_75t_SL g695 ( .A1(n_673), .A2(n_630), .B(n_610), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_659), .B(n_600), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_653), .Y(n_697) );
INVx2_ASAP7_75t_SL g698 ( .A(n_684), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_657), .B(n_631), .Y(n_699) );
OAI31xp33_ASAP7_75t_L g700 ( .A1(n_670), .A2(n_609), .A3(n_637), .B(n_634), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_674), .Y(n_701) );
INVx2_ASAP7_75t_SL g702 ( .A(n_688), .Y(n_702) );
OAI21xp33_ASAP7_75t_L g703 ( .A1(n_662), .A2(n_658), .B(n_650), .Y(n_703) );
NAND2x1_ASAP7_75t_SL g704 ( .A(n_656), .B(n_647), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g705 ( .A1(n_670), .A2(n_633), .B(n_602), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_651), .B(n_627), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_658), .A2(n_647), .B1(n_636), .B2(n_614), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_675), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_687), .A2(n_622), .B1(n_627), .B2(n_614), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g710 ( .A1(n_679), .A2(n_641), .B(n_649), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_676), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_680), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_668), .B(n_613), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_702), .B(n_666), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_697), .A2(n_687), .B(n_664), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_700), .A2(n_667), .B(n_677), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_697), .A2(n_671), .B1(n_669), .B2(n_678), .Y(n_717) );
AOI32xp33_ASAP7_75t_L g718 ( .A1(n_703), .A2(n_682), .A3(n_655), .B1(n_661), .B2(n_665), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_707), .A2(n_654), .B1(n_685), .B2(n_683), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_695), .A2(n_682), .B(n_641), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_690), .A2(n_608), .B1(n_617), .B2(n_618), .C(n_622), .Y(n_721) );
O2A1O1Ixp5_ASAP7_75t_L g722 ( .A1(n_705), .A2(n_635), .B(n_626), .C(n_628), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_690), .A2(n_613), .B1(n_624), .B2(n_628), .C(n_626), .Y(n_723) );
AOI221x1_ASAP7_75t_L g724 ( .A1(n_710), .A2(n_624), .B1(n_686), .B2(n_681), .C(n_217), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_689), .Y(n_725) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_704), .A2(n_355), .B(n_337), .C(n_217), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_706), .B(n_62), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_689), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_725), .Y(n_729) );
NAND4xp25_ASAP7_75t_L g730 ( .A(n_718), .B(n_691), .C(n_699), .D(n_709), .Y(n_730) );
AOI321xp33_ASAP7_75t_L g731 ( .A1(n_716), .A2(n_691), .A3(n_692), .B1(n_696), .B2(n_693), .C(n_708), .Y(n_731) );
NOR4xp25_ASAP7_75t_L g732 ( .A(n_715), .B(n_698), .C(n_711), .D(n_701), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g733 ( .A1(n_720), .A2(n_694), .B(n_713), .C(n_712), .Y(n_733) );
AND3x1_ASAP7_75t_L g734 ( .A(n_715), .B(n_66), .C(n_69), .Y(n_734) );
AOI221xp5_ASAP7_75t_SL g735 ( .A1(n_721), .A2(n_213), .B1(n_217), .B2(n_77), .C(n_70), .Y(n_735) );
OAI211xp5_ASAP7_75t_L g736 ( .A1(n_717), .A2(n_213), .B(n_217), .C(n_74), .Y(n_736) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_722), .A2(n_280), .B(n_281), .C(n_213), .Y(n_737) );
NAND2x1_ASAP7_75t_L g738 ( .A(n_729), .B(n_728), .Y(n_738) );
AOI21xp5_ASAP7_75t_SL g739 ( .A1(n_733), .A2(n_726), .B(n_724), .Y(n_739) );
NAND3xp33_ASAP7_75t_L g740 ( .A(n_731), .B(n_723), .C(n_719), .Y(n_740) );
NOR2x1_ASAP7_75t_L g741 ( .A(n_733), .B(n_727), .Y(n_741) );
BUFx2_ASAP7_75t_L g742 ( .A(n_734), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_740), .B(n_732), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_738), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_742), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_745), .Y(n_746) );
NAND3xp33_ASAP7_75t_SL g747 ( .A(n_743), .B(n_737), .C(n_736), .Y(n_747) );
INVx3_ASAP7_75t_L g748 ( .A(n_746), .Y(n_748) );
OAI221xp5_ASAP7_75t_L g749 ( .A1(n_747), .A2(n_741), .B1(n_744), .B2(n_739), .C(n_730), .Y(n_749) );
AO22x1_ASAP7_75t_L g750 ( .A1(n_748), .A2(n_714), .B1(n_735), .B2(n_213), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_750), .A2(n_749), .B1(n_280), .B2(n_272), .Y(n_751) );
OA331x2_ASAP7_75t_L g752 ( .A1(n_751), .A2(n_264), .A3(n_272), .B1(n_298), .B2(n_749), .B3(n_748), .C1(n_746), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g753 ( .A1(n_752), .A2(n_264), .B(n_272), .Y(n_753) );
endmodule