module real_aes_3008_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_379;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_0), .A2(n_66), .B1(n_152), .B2(n_155), .Y(n_151) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_1), .A2(n_53), .B1(n_90), .B2(n_91), .Y(n_89) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_2), .B(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g192 ( .A(n_3), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_4), .B(n_222), .Y(n_272) );
INVx1_ASAP7_75t_L g318 ( .A(n_5), .Y(n_318) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_6), .A2(n_21), .B1(n_90), .B2(n_94), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_7), .Y(n_332) );
INVx2_ASAP7_75t_L g221 ( .A(n_8), .Y(n_221) );
INVx1_ASAP7_75t_L g282 ( .A(n_9), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_10), .Y(n_160) );
AOI222xp33_ASAP7_75t_SL g106 ( .A1(n_11), .A2(n_35), .B1(n_49), .B2(n_107), .C1(n_114), .C2(n_117), .Y(n_106) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_12), .A2(n_175), .B1(n_176), .B2(n_179), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_12), .Y(n_175) );
INVx1_ASAP7_75t_L g279 ( .A(n_13), .Y(n_279) );
INVx1_ASAP7_75t_SL g265 ( .A(n_14), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g83 ( .A1(n_15), .A2(n_67), .B1(n_84), .B2(n_103), .Y(n_83) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_16), .B(n_232), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_17), .A2(n_45), .B1(n_177), .B2(n_178), .Y(n_176) );
INVx1_ASAP7_75t_L g178 ( .A(n_17), .Y(n_178) );
AOI33xp33_ASAP7_75t_L g298 ( .A1(n_18), .A2(n_40), .A3(n_212), .B1(n_227), .B2(n_299), .B3(n_300), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_19), .A2(n_27), .B1(n_145), .B2(n_148), .Y(n_144) );
INVx1_ASAP7_75t_L g326 ( .A(n_20), .Y(n_326) );
OAI221xp5_ASAP7_75t_L g184 ( .A1(n_21), .A2(n_53), .B1(n_56), .B2(n_185), .C(n_187), .Y(n_184) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_22), .A2(n_68), .B(n_221), .Y(n_220) );
OR2x2_ASAP7_75t_L g223 ( .A(n_22), .B(n_68), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_23), .B(n_253), .Y(n_262) );
INVx3_ASAP7_75t_L g90 ( .A(n_24), .Y(n_90) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_25), .A2(n_57), .B1(n_135), .B2(n_139), .Y(n_134) );
OAI22xp5_ASAP7_75t_L g79 ( .A1(n_26), .A2(n_80), .B1(n_170), .B2(n_171), .Y(n_79) );
INVx1_ASAP7_75t_L g171 ( .A(n_26), .Y(n_171) );
INVx1_ASAP7_75t_SL g101 ( .A(n_28), .Y(n_101) );
INVx1_ASAP7_75t_L g194 ( .A(n_29), .Y(n_194) );
AND2x2_ASAP7_75t_L g216 ( .A(n_29), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g241 ( .A(n_29), .B(n_192), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_30), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_31), .B(n_253), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_32), .A2(n_209), .B1(n_219), .B2(n_222), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_33), .B(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_34), .B(n_232), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_36), .B(n_243), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_37), .B(n_232), .Y(n_319) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_38), .A2(n_56), .B1(n_90), .B2(n_97), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_39), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_39), .A2(n_80), .B1(n_170), .B2(n_218), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_41), .B(n_232), .Y(n_310) );
INVx1_ASAP7_75t_L g213 ( .A(n_42), .Y(n_213) );
INVx1_ASAP7_75t_L g234 ( .A(n_42), .Y(n_234) );
AND2x2_ASAP7_75t_L g311 ( .A(n_43), .B(n_259), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_44), .A2(n_58), .B1(n_225), .B2(n_253), .C(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g177 ( .A(n_45), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_45), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g102 ( .A(n_46), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_47), .B(n_219), .Y(n_334) );
AOI21xp5_ASAP7_75t_SL g248 ( .A1(n_48), .A2(n_225), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g275 ( .A(n_50), .Y(n_275) );
INVx1_ASAP7_75t_L g309 ( .A(n_51), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_52), .A2(n_225), .B(n_308), .Y(n_307) );
INVxp33_ASAP7_75t_L g189 ( .A(n_53), .Y(n_189) );
INVx1_ASAP7_75t_L g217 ( .A(n_54), .Y(n_217) );
INVx1_ASAP7_75t_L g236 ( .A(n_54), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_55), .B(n_253), .Y(n_301) );
INVxp67_ASAP7_75t_L g188 ( .A(n_56), .Y(n_188) );
AND2x2_ASAP7_75t_L g267 ( .A(n_59), .B(n_246), .Y(n_267) );
INVx1_ASAP7_75t_L g276 ( .A(n_60), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_61), .A2(n_225), .B(n_264), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_62), .A2(n_72), .B1(n_123), .B2(n_129), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_63), .A2(n_225), .B(n_230), .C(n_242), .Y(n_224) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_63), .Y(n_569) );
AND2x2_ASAP7_75t_SL g245 ( .A(n_64), .B(n_246), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_65), .A2(n_225), .B1(n_296), .B2(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g250 ( .A(n_69), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_70), .A2(n_80), .B1(n_170), .B2(n_561), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_70), .Y(n_561) );
AND2x2_ASAP7_75t_L g302 ( .A(n_71), .B(n_246), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_73), .A2(n_324), .B(n_325), .C(n_327), .Y(n_323) );
OAI22xp5_ASAP7_75t_SL g172 ( .A1(n_74), .A2(n_173), .B1(n_174), .B2(n_180), .Y(n_172) );
INVx1_ASAP7_75t_L g180 ( .A(n_74), .Y(n_180) );
BUFx2_ASAP7_75t_SL g186 ( .A(n_75), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_76), .B(n_232), .Y(n_251) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_181), .B1(n_195), .B2(n_552), .C(n_553), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_172), .Y(n_78) );
INVx1_ASAP7_75t_L g170 ( .A(n_80), .Y(n_170) );
NAND5xp2_ASAP7_75t_L g80 ( .A(n_81), .B(n_121), .C(n_143), .D(n_158), .E(n_166), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_106), .Y(n_82) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_95), .Y(n_87) );
AND2x2_ASAP7_75t_L g126 ( .A(n_88), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g137 ( .A(n_88), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_92), .Y(n_88) );
AND2x2_ASAP7_75t_L g105 ( .A(n_89), .B(n_93), .Y(n_105) );
INVx2_ASAP7_75t_L g113 ( .A(n_89), .Y(n_113) );
INVx1_ASAP7_75t_L g91 ( .A(n_90), .Y(n_91) );
INVx2_ASAP7_75t_L g94 ( .A(n_90), .Y(n_94) );
INVx1_ASAP7_75t_L g97 ( .A(n_90), .Y(n_97) );
OAI22x1_ASAP7_75t_L g99 ( .A1(n_90), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_90), .Y(n_100) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_92), .Y(n_133) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g112 ( .A(n_93), .Y(n_112) );
AND2x4_ASAP7_75t_L g116 ( .A(n_93), .B(n_113), .Y(n_116) );
AND2x4_ASAP7_75t_L g115 ( .A(n_95), .B(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g142 ( .A(n_95), .B(n_111), .Y(n_142) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
BUFx2_ASAP7_75t_L g104 ( .A(n_96), .Y(n_104) );
AND2x2_ASAP7_75t_L g110 ( .A(n_96), .B(n_99), .Y(n_110) );
INVx2_ASAP7_75t_L g128 ( .A(n_96), .Y(n_128) );
AND2x4_ASAP7_75t_L g138 ( .A(n_98), .B(n_128), .Y(n_138) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g127 ( .A(n_99), .B(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_99), .Y(n_157) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x4_ASAP7_75t_L g150 ( .A(n_105), .B(n_138), .Y(n_150) );
AND2x2_ASAP7_75t_L g156 ( .A(n_105), .B(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx6_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x4_ASAP7_75t_L g119 ( .A(n_110), .B(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g131 ( .A(n_110), .B(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g147 ( .A(n_111), .B(n_127), .Y(n_147) );
AND2x4_ASAP7_75t_L g165 ( .A(n_111), .B(n_138), .Y(n_165) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVxp67_ASAP7_75t_L g120 ( .A(n_113), .Y(n_120) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g154 ( .A(n_116), .B(n_127), .Y(n_154) );
AND2x4_ASAP7_75t_L g169 ( .A(n_116), .B(n_138), .Y(n_169) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx6_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_134), .Y(n_121) );
BUFx3_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx6f_ASAP7_75t_SL g129 ( .A(n_130), .Y(n_129) );
BUFx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx8_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_151), .Y(n_143) );
INVx1_ASAP7_75t_SL g145 ( .A(n_146), .Y(n_145) );
INVx6_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx12f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVxp67_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
INVx8_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_174), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_176), .Y(n_179) );
INVx1_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
AND3x1_ASAP7_75t_SL g183 ( .A(n_184), .B(n_190), .C(n_193), .Y(n_183) );
INVxp67_ASAP7_75t_L g559 ( .A(n_184), .Y(n_559) );
CKINVDCx8_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g557 ( .A(n_190), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_190), .A2(n_210), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g211 ( .A(n_191), .B(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_SL g564 ( .A(n_191), .B(n_193), .Y(n_564) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g229 ( .A(n_192), .B(n_213), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_193), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2x1p5_ASAP7_75t_L g226 ( .A(n_194), .B(n_227), .Y(n_226) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND4xp75_ASAP7_75t_L g200 ( .A(n_201), .B(n_403), .C(n_469), .D(n_532), .Y(n_200) );
NOR2x1_ASAP7_75t_L g201 ( .A(n_202), .B(n_366), .Y(n_201) );
OR3x1_ASAP7_75t_L g202 ( .A(n_203), .B(n_336), .C(n_363), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_268), .B(n_291), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_254), .Y(n_205) );
AND2x2_ASAP7_75t_L g466 ( .A(n_206), .B(n_436), .Y(n_466) );
INVx1_ASAP7_75t_L g539 ( .A(n_206), .Y(n_539) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_244), .Y(n_206) );
INVx2_ASAP7_75t_L g290 ( .A(n_207), .Y(n_290) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_207), .Y(n_354) );
AND2x2_ASAP7_75t_L g358 ( .A(n_207), .B(n_271), .Y(n_358) );
AND2x4_ASAP7_75t_L g374 ( .A(n_207), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g378 ( .A(n_207), .Y(n_378) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_224), .Y(n_207) );
NOR3xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_214), .C(n_218), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x4_ASAP7_75t_L g253 ( .A(n_211), .B(n_215), .Y(n_253) );
OR2x6_ASAP7_75t_L g239 ( .A(n_212), .B(n_228), .Y(n_239) );
INVxp33_ASAP7_75t_L g299 ( .A(n_212), .Y(n_299) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x4_ASAP7_75t_L g284 ( .A(n_213), .B(n_235), .Y(n_284) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g228 ( .A(n_217), .Y(n_228) );
AND2x6_ASAP7_75t_L g281 ( .A(n_217), .B(n_233), .Y(n_281) );
INVx4_ASAP7_75t_L g246 ( .A(n_219), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_219), .B(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx4f_ASAP7_75t_L g243 ( .A(n_220), .Y(n_243) );
AND2x4_ASAP7_75t_L g222 ( .A(n_221), .B(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_SL g260 ( .A(n_221), .B(n_223), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_222), .A2(n_248), .B(n_252), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_222), .B(n_240), .Y(n_285) );
INVxp67_ASAP7_75t_L g333 ( .A(n_225), .Y(n_333) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_225), .Y(n_552) );
AND2x4_ASAP7_75t_L g225 ( .A(n_226), .B(n_229), .Y(n_225) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_226), .Y(n_567) );
INVx1_ASAP7_75t_L g300 ( .A(n_227), .Y(n_300) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_237), .B(n_240), .Y(n_230) );
INVx1_ASAP7_75t_L g277 ( .A(n_232), .Y(n_277) );
AND2x4_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_239), .A2(n_240), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_239), .A2(n_240), .B(n_265), .C(n_266), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_239), .A2(n_275), .B1(n_276), .B2(n_277), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_239), .A2(n_240), .B(n_309), .C(n_310), .Y(n_308) );
O2A1O1Ixp33_ASAP7_75t_SL g317 ( .A1(n_239), .A2(n_240), .B(n_318), .C(n_319), .Y(n_317) );
INVxp67_ASAP7_75t_L g324 ( .A(n_239), .Y(n_324) );
INVx1_ASAP7_75t_L g296 ( .A(n_240), .Y(n_296) );
INVx5_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_241), .Y(n_327) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_242), .A2(n_294), .B(n_302), .Y(n_293) );
AO21x2_ASAP7_75t_L g342 ( .A1(n_242), .A2(n_294), .B(n_302), .Y(n_342) );
INVx2_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
OA21x2_ASAP7_75t_L g315 ( .A1(n_243), .A2(n_316), .B(n_320), .Y(n_315) );
AND2x2_ASAP7_75t_L g269 ( .A(n_244), .B(n_270), .Y(n_269) );
INVx4_ASAP7_75t_L g355 ( .A(n_244), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_244), .B(n_345), .Y(n_359) );
INVx2_ASAP7_75t_L g373 ( .A(n_244), .Y(n_373) );
AND2x4_ASAP7_75t_L g377 ( .A(n_244), .B(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_244), .Y(n_412) );
OR2x2_ASAP7_75t_L g418 ( .A(n_244), .B(n_257), .Y(n_418) );
NOR2x1_ASAP7_75t_SL g447 ( .A(n_244), .B(n_271), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_244), .B(n_521), .Y(n_549) );
OR2x6_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
INVx3_ASAP7_75t_L g304 ( .A(n_246), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_246), .A2(n_304), .B1(n_323), .B2(n_328), .Y(n_322) );
INVx1_ASAP7_75t_L g335 ( .A(n_253), .Y(n_335) );
AND2x2_ASAP7_75t_L g446 ( .A(n_254), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2x1_ASAP7_75t_L g480 ( .A(n_255), .B(n_270), .Y(n_480) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g287 ( .A(n_257), .Y(n_287) );
INVx2_ASAP7_75t_L g346 ( .A(n_257), .Y(n_346) );
AND2x2_ASAP7_75t_L g369 ( .A(n_257), .B(n_271), .Y(n_369) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_257), .Y(n_396) );
INVx1_ASAP7_75t_L g437 ( .A(n_257), .Y(n_437) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .B(n_267), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_259), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_286), .Y(n_268) );
AND2x2_ASAP7_75t_L g449 ( .A(n_269), .B(n_344), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_270), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g516 ( .A(n_270), .Y(n_516) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx3_ASAP7_75t_L g375 ( .A(n_271), .Y(n_375) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B(n_285), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_277), .B(n_326), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_280), .B1(n_282), .B2(n_283), .Y(n_278) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI211xp5_ASAP7_75t_SL g452 ( .A1(n_286), .A2(n_453), .B(n_457), .C(n_463), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_SL g368 ( .A(n_288), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g499 ( .A(n_288), .Y(n_499) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g421 ( .A(n_290), .B(n_375), .Y(n_421) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_312), .Y(n_291) );
AOI32xp33_ASAP7_75t_L g457 ( .A1(n_292), .A2(n_441), .A3(n_458), .B1(n_459), .B2(n_461), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_303), .Y(n_292) );
INVx2_ASAP7_75t_L g383 ( .A(n_293), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_293), .B(n_315), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_295), .B(n_301), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx3_ASAP7_75t_L g395 ( .A(n_303), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_303), .B(n_321), .Y(n_426) );
AND2x2_ASAP7_75t_L g431 ( .A(n_303), .B(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_303), .Y(n_513) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_311), .Y(n_303) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_304), .A2(n_305), .B(n_311), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OR2x2_ASAP7_75t_L g414 ( .A(n_312), .B(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g365 ( .A(n_313), .B(n_339), .Y(n_365) );
AND2x2_ASAP7_75t_L g514 ( .A(n_313), .B(n_512), .Y(n_514) );
AND2x4_ASAP7_75t_L g313 ( .A(n_314), .B(n_321), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g351 ( .A(n_315), .Y(n_351) );
AND2x4_ASAP7_75t_L g390 ( .A(n_315), .B(n_391), .Y(n_390) );
INVxp67_ASAP7_75t_L g424 ( .A(n_315), .Y(n_424) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_315), .Y(n_432) );
AND2x2_ASAP7_75t_L g441 ( .A(n_315), .B(n_321), .Y(n_441) );
INVx1_ASAP7_75t_L g525 ( .A(n_315), .Y(n_525) );
INVx2_ASAP7_75t_L g362 ( .A(n_321), .Y(n_362) );
INVx1_ASAP7_75t_L g389 ( .A(n_321), .Y(n_389) );
INVx1_ASAP7_75t_L g456 ( .A(n_321), .Y(n_456) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_329), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B1(n_334), .B2(n_335), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI32xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_347), .A3(n_352), .B1(n_356), .B2(n_360), .Y(n_336) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_338), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_343), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_339), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g440 ( .A(n_339), .B(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g465 ( .A(n_339), .Y(n_465) );
AND2x2_ASAP7_75t_L g546 ( .A(n_339), .B(n_388), .Y(n_546) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g361 ( .A(n_341), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g460 ( .A(n_341), .B(n_383), .Y(n_460) );
NOR2xp67_ASAP7_75t_L g482 ( .A(n_341), .B(n_362), .Y(n_482) );
NOR2x1_ASAP7_75t_L g524 ( .A(n_341), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g391 ( .A(n_342), .Y(n_391) );
INVx1_ASAP7_75t_L g415 ( .A(n_342), .Y(n_415) );
AND2x2_ASAP7_75t_L g430 ( .A(n_342), .B(n_362), .Y(n_430) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g458 ( .A(n_344), .B(n_447), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_344), .B(n_377), .Y(n_528) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_345), .Y(n_497) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_346), .Y(n_479) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g380 ( .A(n_349), .B(n_381), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g464 ( .A(n_349), .B(n_465), .Y(n_464) );
NOR2xp67_ASAP7_75t_SL g551 ( .A(n_349), .B(n_489), .Y(n_551) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g408 ( .A(n_351), .B(n_362), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_352), .B(n_418), .Y(n_476) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_353), .B(n_369), .Y(n_442) );
AND2x4_ASAP7_75t_SL g353 ( .A(n_354), .B(n_355), .Y(n_353) );
NOR2x1_ASAP7_75t_L g401 ( .A(n_355), .B(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g507 ( .A(n_355), .B(n_378), .Y(n_507) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_355), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_356), .B(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
OR2x2_ASAP7_75t_L g478 ( .A(n_357), .B(n_479), .Y(n_478) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_357), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g467 ( .A(n_358), .B(n_412), .Y(n_467) );
INVxp33_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g381 ( .A(n_361), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g541 ( .A(n_361), .B(n_423), .Y(n_541) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_384), .Y(n_366) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B(n_379), .Y(n_367) );
AND2x2_ASAP7_75t_L g502 ( .A(n_369), .B(n_377), .Y(n_502) );
NAND2xp33_ASAP7_75t_R g370 ( .A(n_371), .B(n_376), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g544 ( .A(n_373), .Y(n_544) );
INVx4_ASAP7_75t_L g402 ( .A(n_374), .Y(n_402) );
INVx1_ASAP7_75t_L g521 ( .A(n_375), .Y(n_521) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g515 ( .A(n_377), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_SL g519 ( .A(n_377), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_380), .A2(n_445), .B1(n_549), .B2(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g409 ( .A(n_383), .B(n_395), .Y(n_409) );
AND2x2_ASAP7_75t_L g423 ( .A(n_383), .B(n_424), .Y(n_423) );
A2O1A1Ixp33_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_392), .B(n_397), .C(n_400), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g471 ( .A(n_387), .B(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g399 ( .A(n_388), .Y(n_399) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g459 ( .A(n_389), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g468 ( .A(n_389), .B(n_390), .Y(n_468) );
INVx1_ASAP7_75t_L g500 ( .A(n_389), .Y(n_500) );
AND2x4_ASAP7_75t_L g481 ( .A(n_390), .B(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g503 ( .A(n_390), .B(n_394), .Y(n_503) );
AND2x2_ASAP7_75t_L g511 ( .A(n_390), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVx1_ASAP7_75t_L g486 ( .A(n_394), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_394), .B(n_408), .Y(n_488) );
AND2x2_ASAP7_75t_L g491 ( .A(n_394), .B(n_441), .Y(n_491) );
INVx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_395), .B(n_456), .Y(n_505) );
AND2x2_ASAP7_75t_L g433 ( .A(n_396), .B(n_421), .Y(n_433) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g529 ( .A(n_399), .B(n_409), .Y(n_529) );
BUFx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_401), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g413 ( .A(n_402), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_402), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_443), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_427), .Y(n_404) );
OAI222xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_410), .B1(n_414), .B2(n_416), .C1(n_419), .C2(n_422), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_412), .B(n_421), .Y(n_420) );
OR2x6_ASAP7_75t_L g492 ( .A(n_412), .B(n_462), .Y(n_492) );
NAND5xp2_ASAP7_75t_L g495 ( .A(n_412), .B(n_415), .C(n_431), .D(n_496), .E(n_498), .Y(n_495) );
NAND2x1_ASAP7_75t_L g531 ( .A(n_413), .B(n_417), .Y(n_531) );
INVx2_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_418), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_420), .A2(n_511), .B1(n_514), .B2(n_515), .Y(n_510) );
INVx2_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_421), .B(n_437), .Y(n_474) );
INVx3_ASAP7_75t_L g509 ( .A(n_422), .Y(n_509) );
NAND2x1p5_ASAP7_75t_L g422 ( .A(n_423), .B(n_425), .Y(n_422) );
AND2x2_ASAP7_75t_L g454 ( .A(n_423), .B(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
INVx2_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g450 ( .A(n_426), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_428), .B(n_439), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_433), .B(n_434), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g438 ( .A(n_430), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_433), .A2(n_440), .B1(n_441), .B2(n_442), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_SL g520 ( .A(n_437), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_452), .Y(n_443) );
AOI21xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_448), .B(n_450), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g489 ( .A(n_460), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_466), .B1(n_467), .B2(n_468), .Y(n_463) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_493), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .C(n_483), .Y(n_470) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OA21x2_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_477), .B(n_481), .Y(n_475) );
NAND2xp33_ASAP7_75t_SL g477 ( .A(n_478), .B(n_480), .Y(n_477) );
AOI21xp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_490), .B(n_492), .Y(n_483) );
OAI211xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_487), .B(n_488), .C(n_489), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_487), .A2(n_527), .B1(n_529), .B2(n_530), .Y(n_526) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_517), .Y(n_493) );
NAND4xp25_ASAP7_75t_L g494 ( .A(n_495), .B(n_501), .C(n_508), .D(n_510), .Y(n_494) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g506 ( .A(n_497), .B(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g537 ( .A(n_500), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B1(n_504), .B2(n_506), .Y(n_501) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_506), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI21xp5_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_522), .B(n_526), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_519), .Y(n_518) );
INVxp67_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_547), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_537), .B(n_538), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B1(n_542), .B2(n_545), .Y(n_538) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OAI222xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_560), .B2(n_562), .C1(n_565), .C2(n_568), .Y(n_553) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
endmodule