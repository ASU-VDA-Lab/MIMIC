module fake_jpeg_9055_n_234 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_27),
.B1(n_21),
.B2(n_31),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_54),
.B1(n_31),
.B2(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_22),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_45),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_16),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_16),
.C(n_18),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_19),
.C(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_27),
.B1(n_31),
.B2(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_24),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_36),
.B1(n_31),
.B2(n_40),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_75),
.B1(n_41),
.B2(n_25),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_16),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_62),
.Y(n_92)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_32),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_70),
.Y(n_99)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_67),
.A2(n_41),
.B1(n_39),
.B2(n_33),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_38),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_83),
.B(n_23),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_49),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_76),
.Y(n_103)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_77),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_40),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_18),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_24),
.Y(n_106)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_25),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_98),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_90),
.B(n_106),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_105),
.B1(n_75),
.B2(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_17),
.B(n_29),
.C(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_71),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_78),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_130),
.B1(n_86),
.B2(n_87),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_76),
.C(n_68),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_113),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_76),
.C(n_68),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_74),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_119),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_83),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_66),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_125),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_80),
.C(n_64),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_64),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_77),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_96),
.C(n_100),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_59),
.B1(n_61),
.B2(n_72),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_133),
.B1(n_19),
.B2(n_86),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_41),
.B1(n_62),
.B2(n_60),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_25),
.B1(n_19),
.B2(n_23),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_137),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_142),
.B1(n_147),
.B2(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_90),
.B(n_89),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_125),
.B(n_119),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_28),
.B(n_26),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_154),
.B1(n_123),
.B2(n_91),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

AOI22x1_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_150),
.A2(n_127),
.B1(n_129),
.B2(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_109),
.A2(n_93),
.B1(n_101),
.B2(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_167),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_132),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_168),
.C(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_166),
.B1(n_30),
.B2(n_17),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_113),
.B1(n_112),
.B2(n_124),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_174),
.B1(n_157),
.B2(n_151),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_140),
.B1(n_142),
.B2(n_148),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_116),
.B(n_91),
.C(n_30),
.D(n_20),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_107),
.C(n_39),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_39),
.C(n_33),
.Y(n_170)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_32),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_175),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_153),
.A2(n_33),
.B1(n_23),
.B2(n_29),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_30),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_33),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_170),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_165),
.A2(n_144),
.B1(n_134),
.B2(n_143),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_180),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_185),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_138),
.A3(n_152),
.B1(n_145),
.B2(n_143),
.C1(n_139),
.C2(n_26),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_139),
.B1(n_152),
.B2(n_145),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_189),
.B1(n_190),
.B2(n_2),
.Y(n_201)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_1),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_158),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_171),
.A2(n_164),
.B1(n_167),
.B2(n_169),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_190)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_199),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_160),
.C(n_173),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_201),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_176),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_1),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_187),
.C(n_179),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_2),
.C(n_3),
.Y(n_202)
);

AOI31xp33_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_4),
.A3(n_5),
.B(n_6),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_3),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_190),
.B1(n_189),
.B2(n_191),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_205),
.A2(n_196),
.B(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_188),
.C(n_191),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_213),
.C(n_192),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_211),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_9),
.B(n_10),
.Y(n_215)
);

NOR2x1_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_8),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_8),
.C(n_9),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_204),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_192),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_219),
.B(n_213),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_210),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_205),
.B(n_216),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_207),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_226),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.C(n_223),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_222),
.A2(n_198),
.B(n_10),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_227),
.C(n_10),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_230),
.B1(n_11),
.B2(n_12),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_9),
.Y(n_234)
);


endmodule