module fake_ibex_815_n_888 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_888);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_888;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_357;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_798;
wire n_832;
wire n_732;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_636;
wire n_594;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_562;
wire n_506;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_285;
wire n_379;
wire n_247;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_729;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_231;
wire n_298;
wire n_202;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_54),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_17),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_12),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_87),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_19),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_67),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_27),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_45),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_90),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_37),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_120),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_61),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_136),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_105),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_112),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_43),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_75),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_51),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_70),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_72),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_96),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_29),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_116),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_46),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_139),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_68),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_92),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_42),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_38),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_110),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_104),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_83),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_78),
.B(n_155),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_94),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_124),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_16),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_141),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_149),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_7),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_81),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_125),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_41),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_22),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_153),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_95),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_101),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_44),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_39),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_52),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_119),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_77),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_26),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_154),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_97),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_56),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_74),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_133),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_89),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_114),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_62),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_138),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_147),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_47),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_28),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_71),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_69),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_98),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_159),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_135),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_48),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_163),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_148),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_115),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_91),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_29),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_109),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_121),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_25),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_123),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_157),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_57),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_127),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_113),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_122),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_63),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_34),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_14),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_18),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_145),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_107),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_13),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_84),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_53),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_60),
.B(n_79),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_152),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_177),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_76),
.B(n_162),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_196),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_193),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_169),
.B(n_0),
.Y(n_282)
);

BUFx8_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_193),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_214),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_0),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_194),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_185),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_167),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_214),
.B(n_1),
.Y(n_290)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_196),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_167),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_195),
.Y(n_293)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_185),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_1),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_231),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_195),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_185),
.Y(n_298)
);

BUFx8_ASAP7_75t_L g299 ( 
.A(n_168),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_207),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_217),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_185),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_2),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_201),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_207),
.B(n_2),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g307 ( 
.A(n_173),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_211),
.B(n_3),
.Y(n_309)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_174),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_201),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_211),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_217),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_268),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_171),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_174),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_172),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_272),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_166),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_201),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_224),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_213),
.Y(n_322)
);

BUFx8_ASAP7_75t_L g323 ( 
.A(n_224),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g324 ( 
.A1(n_184),
.A2(n_80),
.B(n_161),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_186),
.B(n_5),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_187),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_210),
.B(n_6),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_188),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_187),
.B(n_222),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_190),
.B(n_6),
.Y(n_330)
);

XNOR2x2_ASAP7_75t_L g331 ( 
.A(n_221),
.B(n_8),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_222),
.B(n_8),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_233),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_172),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_233),
.Y(n_335)
);

INVx5_ASAP7_75t_L g336 ( 
.A(n_213),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_213),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_217),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_242),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_246),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_246),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_198),
.B(n_9),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_203),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_250),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_199),
.B(n_10),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_250),
.B(n_11),
.Y(n_347)
);

BUFx12f_ASAP7_75t_L g348 ( 
.A(n_165),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_178),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_200),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_213),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_288),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_278),
.B(n_216),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_280),
.B(n_204),
.Y(n_357)
);

NAND2xp33_ASAP7_75t_SL g358 ( 
.A(n_287),
.B(n_178),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_307),
.B(n_170),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_280),
.B(n_208),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_290),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_291),
.Y(n_364)
);

NAND2xp33_ASAP7_75t_SL g365 ( 
.A(n_287),
.B(n_191),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_290),
.Y(n_366)
);

BUFx10_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_332),
.B(n_215),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_291),
.B(n_259),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_347),
.B(n_218),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_347),
.B(n_219),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_351),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_291),
.B(n_319),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_289),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_323),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_328),
.B(n_223),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_307),
.Y(n_379)
);

CKINVDCx6p67_ASAP7_75t_R g380 ( 
.A(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_292),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g382 ( 
.A(n_323),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_326),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_277),
.B(n_269),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_292),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_329),
.B(n_175),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_293),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_329),
.B(n_310),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_303),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_293),
.Y(n_390)
);

AO21x2_ASAP7_75t_L g391 ( 
.A1(n_279),
.A2(n_226),
.B(n_225),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_350),
.B(n_228),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_304),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_316),
.B(n_179),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_297),
.Y(n_395)
);

NAND3x1_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_240),
.C(n_238),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_300),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_300),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_312),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_316),
.B(n_241),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_SL g401 ( 
.A(n_282),
.B(n_261),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_308),
.B(n_217),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_342),
.B(n_181),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_311),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_320),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_342),
.B(n_182),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_323),
.B(n_283),
.C(n_299),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_320),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_299),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_283),
.B(n_183),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_333),
.B(n_249),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_335),
.B(n_253),
.Y(n_414)
);

BUFx6f_ASAP7_75t_SL g415 ( 
.A(n_314),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_321),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_317),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_317),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_318),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_281),
.B(n_243),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_284),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_285),
.B(n_254),
.Y(n_422)
);

BUFx10_ASAP7_75t_L g423 ( 
.A(n_327),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_296),
.A2(n_243),
.B1(n_257),
.B2(n_266),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_L g425 ( 
.A1(n_344),
.A2(n_243),
.B1(n_273),
.B2(n_260),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_320),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_L g427 ( 
.A(n_338),
.B(n_189),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_301),
.Y(n_428)
);

CKINVDCx6p67_ASAP7_75t_R g429 ( 
.A(n_295),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_L g430 ( 
.A(n_340),
.B(n_276),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_281),
.B(n_262),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_322),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_354),
.B(n_283),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_353),
.B(n_327),
.Y(n_434)
);

OAI22xp33_ASAP7_75t_L g435 ( 
.A1(n_359),
.A2(n_334),
.B1(n_315),
.B2(n_343),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_353),
.B(n_330),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_360),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_362),
.B(n_346),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_384),
.B(n_341),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_180),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_388),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_341),
.Y(n_443)
);

A2O1A1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_372),
.A2(n_345),
.B(n_279),
.C(n_271),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_377),
.B(n_192),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_363),
.B(n_325),
.Y(n_446)
);

AND3x1_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_331),
.C(n_209),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_379),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_393),
.B(n_306),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_357),
.B(n_197),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_382),
.B(n_202),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_361),
.B(n_386),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_313),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_356),
.A2(n_309),
.B1(n_252),
.B2(n_270),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_418),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_402),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_205),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_420),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_356),
.B(n_206),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_366),
.A2(n_309),
.B1(n_243),
.B2(n_313),
.Y(n_461)
);

BUFx6f_ASAP7_75t_SL g462 ( 
.A(n_411),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_367),
.B(n_212),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_421),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_403),
.B(n_220),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_420),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_428),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_380),
.B(n_15),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_369),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_376),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_368),
.B(n_227),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_415),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_358),
.B(n_17),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_381),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_385),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_387),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_371),
.B(n_229),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_371),
.B(n_373),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_370),
.B(n_232),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_373),
.B(n_234),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_397),
.Y(n_483)
);

BUFx6f_ASAP7_75t_SL g484 ( 
.A(n_364),
.Y(n_484)
);

NOR3xp33_ASAP7_75t_L g485 ( 
.A(n_425),
.B(n_247),
.C(n_237),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_396),
.A2(n_251),
.B1(n_248),
.B2(n_236),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_398),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_401),
.A2(n_264),
.B1(n_263),
.B2(n_239),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_425),
.A2(n_274),
.B1(n_244),
.B2(n_245),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_399),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_375),
.B(n_176),
.Y(n_491)
);

NAND2x1p5_ASAP7_75t_L g492 ( 
.A(n_392),
.B(n_324),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_416),
.Y(n_493)
);

AND2x4_ASAP7_75t_SL g494 ( 
.A(n_429),
.B(n_230),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_394),
.B(n_209),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_365),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_431),
.B(n_302),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_378),
.B(n_339),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_413),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_392),
.B(n_339),
.Y(n_500)
);

AOI221xp5_ASAP7_75t_L g501 ( 
.A1(n_422),
.A2(n_235),
.B1(n_230),
.B2(n_322),
.C(n_337),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_431),
.B(n_235),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_391),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_391),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_404),
.B(n_408),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_427),
.B(n_235),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_430),
.B(n_235),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_414),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_400),
.B(n_294),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_444),
.A2(n_424),
.B(n_426),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_453),
.A2(n_439),
.B(n_436),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_448),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_443),
.Y(n_513)
);

A2O1A1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_442),
.A2(n_322),
.B(n_337),
.C(n_294),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_472),
.Y(n_515)
);

A2O1A1Ixp33_ASAP7_75t_L g516 ( 
.A1(n_446),
.A2(n_467),
.B(n_434),
.C(n_495),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_478),
.A2(n_305),
.B1(n_336),
.B2(n_337),
.Y(n_517)
);

AOI33xp33_ASAP7_75t_L g518 ( 
.A1(n_435),
.A2(n_432),
.A3(n_410),
.B1(n_407),
.B2(n_406),
.B3(n_405),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_456),
.B(n_20),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_485),
.A2(n_305),
.B1(n_336),
.B2(n_405),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_440),
.B(n_21),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_470),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_449),
.A2(n_433),
.B1(n_441),
.B2(n_489),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_462),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_464),
.B(n_21),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_465),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_470),
.B(n_22),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_476),
.B(n_23),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_457),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_454),
.B(n_23),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_466),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_508),
.A2(n_374),
.B1(n_355),
.B2(n_389),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_496),
.B(n_24),
.Y(n_534)
);

AND2x6_ASAP7_75t_SL g535 ( 
.A(n_458),
.B(n_24),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_492),
.A2(n_352),
.B(n_355),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_471),
.A2(n_482),
.B(n_477),
.Y(n_537)
);

CKINVDCx10_ASAP7_75t_R g538 ( 
.A(n_462),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_494),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_468),
.B(n_27),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_459),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_473),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_486),
.B(n_30),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_455),
.B(n_31),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_460),
.B(n_31),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_475),
.B(n_32),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_479),
.B(n_32),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_445),
.B(n_33),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_490),
.B(n_33),
.Y(n_549)
);

BUFx12f_ASAP7_75t_L g550 ( 
.A(n_491),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_499),
.Y(n_551)
);

NOR2xp67_ASAP7_75t_L g552 ( 
.A(n_488),
.B(n_34),
.Y(n_552)
);

O2A1O1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_474),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_501),
.B(n_35),
.C(n_36),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_461),
.B(n_49),
.C(n_50),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_497),
.Y(n_556)
);

AO21x1_ASAP7_75t_L g557 ( 
.A1(n_491),
.A2(n_55),
.B(n_58),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_438),
.B(n_59),
.Y(n_558)
);

A2O1A1Ixp33_ASAP7_75t_L g559 ( 
.A1(n_480),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_559)
);

BUFx4f_ASAP7_75t_L g560 ( 
.A(n_438),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_451),
.B(n_73),
.Y(n_561)
);

BUFx12f_ASAP7_75t_L g562 ( 
.A(n_469),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_483),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_484),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_487),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_493),
.Y(n_566)
);

AO32x2_ASAP7_75t_L g567 ( 
.A1(n_447),
.A2(n_82),
.A3(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_450),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_463),
.B(n_102),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_437),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_563),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_511),
.B(n_513),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_529),
.B(n_452),
.Y(n_573)
);

BUFx12f_ASAP7_75t_L g574 ( 
.A(n_524),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_512),
.B(n_498),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_562),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_526),
.B(n_542),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_537),
.A2(n_481),
.B(n_509),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_523),
.A2(n_500),
.B1(n_506),
.B2(n_507),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_538),
.Y(n_580)
);

BUFx10_ASAP7_75t_L g581 ( 
.A(n_531),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_565),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_564),
.B(n_484),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_532),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_550),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_556),
.B(n_530),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_510),
.A2(n_117),
.B(n_118),
.Y(n_587)
);

BUFx8_ASAP7_75t_L g588 ( 
.A(n_515),
.Y(n_588)
);

NOR2x1_ASAP7_75t_SL g589 ( 
.A(n_564),
.B(n_134),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_560),
.Y(n_590)
);

BUFx2_ASAP7_75t_SL g591 ( 
.A(n_524),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_543),
.B(n_140),
.Y(n_592)
);

O2A1O1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_544),
.A2(n_144),
.B(n_150),
.C(n_151),
.Y(n_593)
);

AO32x2_ASAP7_75t_L g594 ( 
.A1(n_517),
.A2(n_568),
.A3(n_567),
.B1(n_518),
.B2(n_551),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_521),
.B(n_540),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_519),
.B(n_545),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_546),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_547),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_522),
.B(n_534),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_549),
.Y(n_600)
);

OAI21xp33_ASAP7_75t_SL g601 ( 
.A1(n_527),
.A2(n_528),
.B(n_525),
.Y(n_601)
);

OAI21x1_ASAP7_75t_SL g602 ( 
.A1(n_557),
.A2(n_569),
.B(n_553),
.Y(n_602)
);

AO21x2_ASAP7_75t_L g603 ( 
.A1(n_514),
.A2(n_559),
.B(n_555),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_552),
.B(n_548),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_570),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g606 ( 
.A1(n_520),
.A2(n_554),
.B(n_555),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_554),
.A2(n_561),
.B(n_533),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_539),
.B(n_541),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_567),
.A2(n_511),
.B(n_516),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_535),
.A2(n_511),
.B(n_516),
.Y(n_610)
);

OA22x2_ASAP7_75t_L g611 ( 
.A1(n_512),
.A2(n_317),
.B1(n_334),
.B2(n_417),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_511),
.A2(n_516),
.B(n_537),
.C(n_505),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_563),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_563),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_512),
.B(n_393),
.Y(n_615)
);

AOI31xp67_ASAP7_75t_L g616 ( 
.A1(n_558),
.A2(n_503),
.A3(n_504),
.B(n_502),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_562),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_563),
.Y(n_618)
);

NAND2x1_ASAP7_75t_L g619 ( 
.A(n_522),
.B(n_470),
.Y(n_619)
);

NOR2xp67_ASAP7_75t_SL g620 ( 
.A(n_512),
.B(n_379),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_511),
.B(n_513),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_511),
.A2(n_516),
.B(n_537),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_511),
.A2(n_516),
.B(n_537),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_511),
.A2(n_516),
.B(n_537),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_511),
.B(n_513),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_511),
.B(n_513),
.Y(n_626)
);

AO31x2_ASAP7_75t_L g627 ( 
.A1(n_536),
.A2(n_444),
.A3(n_557),
.B(n_504),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_512),
.B(n_456),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_563),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_563),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_511),
.A2(n_516),
.B(n_537),
.C(n_505),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_512),
.B(n_393),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_512),
.B(n_448),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_538),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_512),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_512),
.B(n_448),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_513),
.A2(n_529),
.B1(n_516),
.B2(n_511),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_511),
.A2(n_516),
.B(n_537),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_511),
.B(n_513),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_512),
.B(n_456),
.Y(n_640)
);

AO31x2_ASAP7_75t_L g641 ( 
.A1(n_536),
.A2(n_444),
.A3(n_557),
.B(n_504),
.Y(n_641)
);

INVx5_ASAP7_75t_L g642 ( 
.A(n_562),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_511),
.A2(n_516),
.B(n_537),
.Y(n_643)
);

AO31x2_ASAP7_75t_L g644 ( 
.A1(n_536),
.A2(n_444),
.A3(n_557),
.B(n_504),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_511),
.A2(n_516),
.B(n_537),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_566),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_635),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_SL g648 ( 
.A1(n_625),
.A2(n_637),
.B(n_572),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_642),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_SL g650 ( 
.A1(n_583),
.A2(n_642),
.B1(n_581),
.B2(n_611),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_612),
.A2(n_631),
.B(n_622),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_584),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_633),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_642),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_636),
.Y(n_655)
);

AOI221x1_ASAP7_75t_L g656 ( 
.A1(n_623),
.A2(n_645),
.B1(n_643),
.B2(n_638),
.C(n_624),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_610),
.A2(n_615),
.B1(n_632),
.B2(n_597),
.Y(n_657)
);

OAI211xp5_ASAP7_75t_L g658 ( 
.A1(n_604),
.A2(n_601),
.B(n_628),
.C(n_640),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_620),
.B(n_577),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_617),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_637),
.A2(n_639),
.B(n_621),
.C(n_626),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g662 ( 
.A(n_581),
.B(n_583),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_571),
.B(n_582),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_617),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_586),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_617),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_576),
.B(n_605),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_598),
.A2(n_600),
.B1(n_595),
.B2(n_596),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_613),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_601),
.A2(n_614),
.B1(n_630),
.B2(n_629),
.Y(n_670)
);

OA21x2_ASAP7_75t_L g671 ( 
.A1(n_587),
.A2(n_606),
.B(n_578),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_576),
.B(n_575),
.Y(n_672)
);

CKINVDCx6p67_ASAP7_75t_R g673 ( 
.A(n_574),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_618),
.Y(n_674)
);

NAND3xp33_ASAP7_75t_L g675 ( 
.A(n_607),
.B(n_579),
.C(n_593),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_580),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_592),
.A2(n_579),
.B(n_599),
.C(n_573),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_590),
.B(n_646),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_588),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_585),
.B(n_591),
.Y(n_680)
);

AOI211xp5_ASAP7_75t_L g681 ( 
.A1(n_634),
.A2(n_608),
.B(n_588),
.C(n_594),
.Y(n_681)
);

AO31x2_ASAP7_75t_L g682 ( 
.A1(n_594),
.A2(n_616),
.A3(n_627),
.B(n_641),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_619),
.A2(n_594),
.B(n_627),
.Y(n_683)
);

BUFx2_ASAP7_75t_R g684 ( 
.A(n_603),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_SL g685 ( 
.A1(n_641),
.A2(n_334),
.B1(n_317),
.B2(n_635),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_641),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_644),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_644),
.A2(n_611),
.B1(n_610),
.B2(n_485),
.Y(n_688)
);

OAI22x1_ASAP7_75t_L g689 ( 
.A1(n_635),
.A2(n_317),
.B1(n_334),
.B2(n_417),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_609),
.A2(n_631),
.B(n_612),
.Y(n_690)
);

CKINVDCx6p67_ASAP7_75t_R g691 ( 
.A(n_642),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_609),
.A2(n_631),
.B(n_612),
.Y(n_692)
);

NAND2x1p5_ASAP7_75t_L g693 ( 
.A(n_642),
.B(n_560),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_584),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_584),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_580),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_642),
.B(n_513),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_637),
.A2(n_523),
.B1(n_529),
.B2(n_513),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_610),
.A2(n_601),
.B(n_511),
.C(n_545),
.Y(n_699)
);

NOR2xp67_ASAP7_75t_SL g700 ( 
.A(n_642),
.B(n_580),
.Y(n_700)
);

OAI21x1_ASAP7_75t_SL g701 ( 
.A1(n_589),
.A2(n_587),
.B(n_610),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_633),
.B(n_636),
.Y(n_702)
);

AOI21xp33_ASAP7_75t_L g703 ( 
.A1(n_601),
.A2(n_602),
.B(n_637),
.Y(n_703)
);

NOR2x1_ASAP7_75t_SL g704 ( 
.A(n_642),
.B(n_591),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_615),
.B(n_632),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_611),
.A2(n_610),
.B1(n_485),
.B2(n_542),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_612),
.A2(n_631),
.B(n_645),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_584),
.Y(n_708)
);

INVx6_ASAP7_75t_L g709 ( 
.A(n_642),
.Y(n_709)
);

OAI211xp5_ASAP7_75t_L g710 ( 
.A1(n_610),
.A2(n_349),
.B(n_523),
.C(n_552),
.Y(n_710)
);

AO21x1_ASAP7_75t_L g711 ( 
.A1(n_609),
.A2(n_587),
.B(n_622),
.Y(n_711)
);

AOI222xp33_ASAP7_75t_L g712 ( 
.A1(n_586),
.A2(n_435),
.B1(n_344),
.B2(n_358),
.C1(n_542),
.C2(n_315),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_642),
.B(n_456),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_633),
.B(n_317),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_611),
.A2(n_610),
.B1(n_485),
.B2(n_542),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_642),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_635),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_665),
.B(n_698),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_697),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_685),
.A2(n_657),
.B1(n_714),
.B2(n_705),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_685),
.A2(n_715),
.B1(n_706),
.B2(n_712),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_661),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_678),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_710),
.B(n_672),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_693),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_699),
.B(n_670),
.Y(n_726)
);

OA21x2_ASAP7_75t_L g727 ( 
.A1(n_656),
.A2(n_692),
.B(n_690),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_652),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_670),
.B(n_651),
.Y(n_729)
);

HB1xp67_ASAP7_75t_L g730 ( 
.A(n_647),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_702),
.B(n_653),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_694),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_709),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_695),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_717),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_708),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_655),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_651),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_663),
.B(n_668),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_709),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_693),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_668),
.A2(n_677),
.B1(n_710),
.B2(n_650),
.Y(n_742)
);

OA21x2_ASAP7_75t_L g743 ( 
.A1(n_690),
.A2(n_692),
.B(n_707),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_688),
.B(n_674),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_669),
.B(n_687),
.Y(n_745)
);

OR2x6_ASAP7_75t_L g746 ( 
.A(n_648),
.B(n_701),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_649),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_664),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_654),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_686),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_681),
.B(n_703),
.C(n_683),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_682),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_654),
.Y(n_753)
);

BUFx2_ASAP7_75t_SL g754 ( 
.A(n_716),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_711),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_664),
.Y(n_756)
);

BUFx5_ASAP7_75t_L g757 ( 
.A(n_667),
.Y(n_757)
);

INVxp67_ASAP7_75t_SL g758 ( 
.A(n_659),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_691),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_671),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_660),
.Y(n_761)
);

NOR2x1p5_ASAP7_75t_L g762 ( 
.A(n_751),
.B(n_726),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_729),
.B(n_684),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_729),
.B(n_675),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_723),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_750),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_750),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_730),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_729),
.B(n_658),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_726),
.B(n_658),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_754),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_726),
.B(n_704),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_SL g773 ( 
.A1(n_742),
.A2(n_662),
.B1(n_679),
.B2(n_680),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_746),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_738),
.B(n_718),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_752),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_725),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_760),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_757),
.B(n_689),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_718),
.B(n_712),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_739),
.B(n_666),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_745),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_735),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_727),
.B(n_713),
.Y(n_784)
);

AO31x2_ASAP7_75t_L g785 ( 
.A1(n_722),
.A2(n_700),
.A3(n_673),
.B(n_696),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_739),
.B(n_676),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_727),
.B(n_743),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_776),
.Y(n_788)
);

OR2x6_ASAP7_75t_L g789 ( 
.A(n_774),
.B(n_746),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_765),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_768),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_766),
.B(n_745),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_775),
.B(n_764),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_780),
.B(n_728),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_771),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_778),
.Y(n_796)
);

NOR2x1_ASAP7_75t_L g797 ( 
.A(n_779),
.B(n_754),
.Y(n_797)
);

OR2x6_ASAP7_75t_SL g798 ( 
.A(n_780),
.B(n_751),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_787),
.B(n_743),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_769),
.B(n_743),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_769),
.B(n_755),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_766),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_767),
.B(n_731),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_763),
.B(n_755),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_783),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_763),
.B(n_727),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_788),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_793),
.B(n_782),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_791),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_800),
.B(n_806),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_802),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_790),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_796),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_805),
.Y(n_814)
);

AND2x2_ASAP7_75t_SL g815 ( 
.A(n_802),
.B(n_774),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_793),
.B(n_782),
.Y(n_816)
);

OAI22xp33_ASAP7_75t_L g817 ( 
.A1(n_798),
.A2(n_771),
.B1(n_777),
.B2(n_772),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_794),
.B(n_786),
.Y(n_818)
);

NAND2x1_ASAP7_75t_L g819 ( 
.A(n_797),
.B(n_772),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_789),
.B(n_799),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_799),
.B(n_770),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_807),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_811),
.Y(n_823)
);

AOI22x1_ASAP7_75t_L g824 ( 
.A1(n_811),
.A2(n_772),
.B1(n_759),
.B2(n_762),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_819),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_818),
.B(n_801),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_809),
.B(n_801),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_819),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_820),
.B(n_789),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_807),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_817),
.B(n_795),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_813),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_812),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_808),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_820),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_825),
.A2(n_772),
.B(n_773),
.C(n_820),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_835),
.B(n_810),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_831),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_824),
.A2(n_773),
.B(n_786),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_835),
.B(n_810),
.Y(n_840)
);

OAI322xp33_ASAP7_75t_L g841 ( 
.A1(n_833),
.A2(n_816),
.A3(n_792),
.B1(n_803),
.B2(n_814),
.C1(n_821),
.C2(n_724),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_834),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_827),
.B(n_821),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_822),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_822),
.Y(n_845)
);

NAND2x2_ASAP7_75t_L g846 ( 
.A(n_825),
.B(n_762),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_832),
.Y(n_847)
);

AOI21xp33_ASAP7_75t_SL g848 ( 
.A1(n_838),
.A2(n_824),
.B(n_828),
.Y(n_848)
);

OAI221xp5_ASAP7_75t_L g849 ( 
.A1(n_838),
.A2(n_823),
.B1(n_828),
.B2(n_721),
.C(n_826),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_842),
.B(n_841),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_839),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_849),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_850),
.A2(n_851),
.B1(n_836),
.B2(n_846),
.Y(n_853)
);

OAI221xp5_ASAP7_75t_L g854 ( 
.A1(n_848),
.A2(n_836),
.B1(n_846),
.B2(n_720),
.C(n_845),
.Y(n_854)
);

AOI222xp33_ASAP7_75t_L g855 ( 
.A1(n_852),
.A2(n_837),
.B1(n_840),
.B2(n_758),
.C1(n_844),
.C2(n_737),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_853),
.Y(n_856)
);

NAND4xp25_ASAP7_75t_L g857 ( 
.A(n_856),
.B(n_854),
.C(n_725),
.D(n_761),
.Y(n_857)
);

NAND3xp33_ASAP7_75t_L g858 ( 
.A(n_855),
.B(n_747),
.C(n_753),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_857),
.B(n_798),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_858),
.B(n_843),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_859),
.B(n_740),
.C(n_733),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_860),
.Y(n_862)
);

XNOR2x1_ASAP7_75t_L g863 ( 
.A(n_862),
.B(n_731),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_861),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_862),
.Y(n_865)
);

OAI22x1_ASAP7_75t_L g866 ( 
.A1(n_865),
.A2(n_740),
.B1(n_733),
.B2(n_741),
.Y(n_866)
);

AOI221x1_ASAP7_75t_L g867 ( 
.A1(n_864),
.A2(n_741),
.B1(n_749),
.B2(n_736),
.C(n_734),
.Y(n_867)
);

OAI22xp5_ASAP7_75t_SL g868 ( 
.A1(n_864),
.A2(n_815),
.B1(n_741),
.B2(n_829),
.Y(n_868)
);

AOI21x1_ASAP7_75t_L g869 ( 
.A1(n_863),
.A2(n_719),
.B(n_829),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_863),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_870),
.A2(n_795),
.B1(n_829),
.B2(n_815),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_867),
.B(n_785),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_868),
.A2(n_784),
.B1(n_847),
.B2(n_830),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_866),
.B(n_749),
.C(n_748),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_869),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_870),
.B(n_748),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_870),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_877),
.A2(n_781),
.B1(n_803),
.B2(n_792),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_875),
.Y(n_879)
);

OA21x2_ASAP7_75t_L g880 ( 
.A1(n_876),
.A2(n_732),
.B(n_736),
.Y(n_880)
);

AO21x2_ASAP7_75t_L g881 ( 
.A1(n_872),
.A2(n_734),
.B(n_732),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_879),
.A2(n_880),
.B(n_878),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_SL g883 ( 
.A1(n_880),
.A2(n_881),
.B1(n_871),
.B2(n_874),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_879),
.A2(n_873),
.B(n_749),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_882),
.A2(n_756),
.B(n_744),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_883),
.B(n_785),
.Y(n_886)
);

OR2x6_ASAP7_75t_L g887 ( 
.A(n_886),
.B(n_884),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_887),
.A2(n_885),
.B1(n_784),
.B2(n_804),
.Y(n_888)
);


endmodule