module real_jpeg_7423_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_0),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_0),
.B(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_0),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_0),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_0),
.B(n_350),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_0),
.B(n_405),
.Y(n_404)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_1),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_1),
.Y(n_193)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_1),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_1),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_2),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_2),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_2),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_2),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_2),
.B(n_154),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_2),
.B(n_337),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_2),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_2),
.B(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_3),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_3),
.Y(n_364)
);

BUFx5_ASAP7_75t_L g403 ( 
.A(n_3),
.Y(n_403)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_3),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_4),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_4),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_4),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_4),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_4),
.B(n_166),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_4),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_4),
.B(n_479),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_5),
.Y(n_102)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_5),
.Y(n_378)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_5),
.Y(n_480)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_6),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_7),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_7),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_7),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_7),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_7),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_7),
.B(n_350),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_7),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_7),
.B(n_491),
.Y(n_490)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_8),
.Y(n_139)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_8),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_8),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_8),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_9),
.Y(n_537)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_11),
.Y(n_160)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_11),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_12),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_12),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_12),
.B(n_138),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_12),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_12),
.B(n_162),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_12),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_12),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_12),
.B(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_13),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_13),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g358 ( 
.A(n_13),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_13),
.B(n_393),
.Y(n_437)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_15),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_15),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_15),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_15),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_15),
.B(n_117),
.Y(n_286)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_17),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_17),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_17),
.B(n_38),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_17),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_17),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_17),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_17),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_18),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_18),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_18),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_18),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_18),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_18),
.B(n_317),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_19),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_19),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_19),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_19),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_19),
.B(n_138),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_19),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_19),
.B(n_364),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_532),
.B(n_534),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_74),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_24),
.B(n_44),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_26),
.A2(n_27),
.B1(n_37),
.B2(n_57),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_37),
.C(n_41),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_28),
.B(n_382),
.Y(n_381)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_48),
.C(n_52),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_39),
.Y(n_317)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_40),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_70),
.C(n_72),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_45),
.B(n_522),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_58),
.C(n_60),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_46),
.A2(n_47),
.B1(n_518),
.B2(n_519),
.Y(n_517)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_61),
.C(n_66),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_51),
.A2(n_52),
.B1(n_66),
.B2(n_481),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_54),
.Y(n_154)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_56),
.Y(n_168)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_56),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_56),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_58),
.B(n_60),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_61),
.A2(n_62),
.B1(n_483),
.B2(n_484),
.Y(n_482)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_66),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_66),
.A2(n_436),
.B1(n_437),
.B2(n_481),
.Y(n_497)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_67),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_68),
.Y(n_247)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_69),
.Y(n_345)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_69),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_523),
.Y(n_522)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_72),
.Y(n_523)
);

AO21x1_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_451),
.B(n_525),
.Y(n_75)
);

OAI21x1_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_412),
.B(n_450),
.Y(n_76)
);

AOI21x1_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_368),
.B(n_411),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_321),
.B(n_367),
.Y(n_78)
);

AOI21x1_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_279),
.B(n_320),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_198),
.B(n_278),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_183),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_82),
.B(n_183),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_126),
.B2(n_182),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_83),
.B(n_127),
.C(n_163),
.Y(n_319)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_103),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_85),
.B(n_104),
.C(n_125),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_98),
.C(n_101),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_86),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_188)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_91),
.Y(n_205)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_91),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_91),
.Y(n_383)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_97),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_98),
.B(n_101),
.Y(n_197)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_100),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_100),
.Y(n_434)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_100),
.Y(n_471)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_102),
.Y(n_348)
);

INVx3_ASAP7_75t_SL g442 ( 
.A(n_102),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_113),
.B1(n_124),
.B2(n_125),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_112),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_108),
.Y(n_112)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_112),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_112),
.B(n_284),
.C(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_114),
.B(n_119),
.C(n_122),
.Y(n_318)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_163),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_143),
.C(n_155),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_140),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_135),
.C(n_140),
.Y(n_181)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_133),
.Y(n_350)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_139),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_141),
.Y(n_447)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_143),
.A2(n_144),
.B1(n_155),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.C(n_152),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_145),
.A2(n_146),
.B1(n_152),
.B2(n_153),
.Y(n_271)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_147),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_150),
.Y(n_306)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_161),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_157),
.B(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_157),
.B(n_460),
.Y(n_459)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

BUFx8_ASAP7_75t_L g357 ( 
.A(n_160),
.Y(n_357)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_162),
.Y(n_235)
);

XOR2x1_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_179),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_164),
.B(n_180),
.C(n_181),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_165),
.B(n_173),
.C(n_177),
.Y(n_297)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_169)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_172),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_176),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_196),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_184),
.B(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_187),
.B(n_196),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_189),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_190),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_194),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21x1_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_273),
.B(n_277),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_258),
.B(n_272),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_238),
.B(n_257),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_225),
.B(n_237),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_209),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_209),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_219),
.B2(n_220),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_212),
.B(n_216),
.C(n_219),
.Y(n_256)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g335 ( 
.A(n_215),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_224),
.Y(n_242)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_232),
.B(n_236),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_228),
.Y(n_236)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_256),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_256),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_242),
.C(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_253),
.C(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

INVx11_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_248)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_249),
.Y(n_255)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_261),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_268),
.C(n_269),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_319),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_319),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_299),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_283),
.C(n_299),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_296),
.B2(n_298),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_286),
.B(n_289),
.C(n_291),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_302),
.C(n_312),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_312),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_308),
.C(n_309),
.Y(n_352)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_318),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_316),
.C(n_318),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_323),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_324),
.B(n_341),
.C(n_365),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_341),
.B1(n_365),
.B2(n_366),
.Y(n_325)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_329),
.B2(n_340),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_330),
.C(n_331),
.Y(n_370)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_329),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_339),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_333),
.B(n_336),
.C(n_339),
.Y(n_399)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx6_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_341),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_351),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_342),
.B(n_352),
.C(n_353),
.Y(n_397)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_342),
.Y(n_539)
);

FAx1_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_346),
.CI(n_349),
.CON(n_342),
.SN(n_342)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_343),
.B(n_346),
.C(n_349),
.Y(n_408)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_362),
.B2(n_363),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_358),
.B1(n_360),
.B2(n_361),
.Y(n_355)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_356),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_361),
.C(n_362),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_358),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_358),
.A2(n_361),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_361),
.B(n_375),
.C(n_381),
.Y(n_424)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_410),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_369),
.B(n_410),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_370),
.B(n_372),
.C(n_395),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_395),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_384),
.B2(n_394),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_373),
.B(n_385),
.C(n_386),
.Y(n_418)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_379),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_380),
.A2(n_381),
.B1(n_436),
.B2(n_437),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_380),
.B(n_432),
.C(n_436),
.Y(n_498)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_384),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_392),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_388),
.B(n_389),
.C(n_392),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_397),
.B1(n_398),
.B2(n_409),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_399),
.C(n_400),
.Y(n_414)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_398),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_408),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_404),
.B1(n_406),
.B2(n_407),
.Y(n_401)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_402),
.Y(n_406)
);

INVx8_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_404),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_406),
.C(n_422),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_404),
.A2(n_407),
.B1(n_426),
.B2(n_429),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_407),
.B(n_424),
.C(n_429),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_408),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_449),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_413),
.B(n_449),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_414),
.B(n_416),
.C(n_430),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_430),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_417),
.B(n_421),
.C(n_423),
.Y(n_506)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_423),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_426),
.Y(n_429)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_438),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_439),
.C(n_440),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_436),
.B(n_478),
.C(n_481),
.Y(n_477)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_441),
.B(n_445),
.C(n_448),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_446),
.B2(n_448),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_444),
.Y(n_448)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NOR3xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_510),
.C(n_520),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_507),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_454),
.A2(n_529),
.B(n_530),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_500),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_455),
.B(n_500),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_474),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_456),
.B(n_475),
.C(n_495),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.C(n_472),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_457),
.B(n_502),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_458),
.A2(n_472),
.B1(n_473),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_458),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_463),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_464),
.C(n_467),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_467),
.Y(n_463)
);

INVx6_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_495),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_487),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_477),
.A2(n_482),
.B1(n_485),
.B2(n_486),
.Y(n_476)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_477),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_477),
.B(n_486),
.C(n_487),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_497),
.Y(n_496)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_480),
.Y(n_491)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_482),
.Y(n_486)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_492),
.C(n_494),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_492),
.B1(n_493),
.B2(n_494),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_490),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_498),
.C(n_499),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_505),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_499),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_504),
.C(n_506),
.Y(n_500)
);

FAx1_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_504),
.CI(n_506),
.CON(n_508),
.SN(n_508)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_509),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_508),
.B(n_509),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_508),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_511),
.B(n_528),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_512),
.B(n_513),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_516),
.C(n_517),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

A2O1A1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_520),
.A2(n_526),
.B(n_527),
.C(n_531),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_521),
.B(n_524),
.Y(n_531)
);

INVx8_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx13_ASAP7_75t_L g536 ( 
.A(n_533),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_537),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);


endmodule