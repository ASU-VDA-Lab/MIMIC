module fake_jpeg_23946_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_13),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_42),
.B(n_44),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_57),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_27),
.B1(n_25),
.B2(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_54),
.A2(n_60),
.B1(n_75),
.B2(n_81),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_20),
.B1(n_36),
.B2(n_38),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_46),
.B1(n_41),
.B2(n_19),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_63),
.Y(n_105)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_27),
.B1(n_22),
.B2(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_21),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_20),
.B(n_18),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_79),
.C(n_32),
.Y(n_89)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_71),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_10),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_68),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_22),
.B1(n_25),
.B2(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_21),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_23),
.B1(n_28),
.B2(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_35),
.Y(n_82)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_36),
.B1(n_31),
.B2(n_23),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_38),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_31),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_85),
.B(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_0),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_88),
.B(n_26),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_115),
.Y(n_133)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_92),
.Y(n_148)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_98),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_41),
.B(n_33),
.C(n_28),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_96),
.A2(n_29),
.B(n_26),
.Y(n_154)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_110),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_46),
.B1(n_44),
.B2(n_17),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_116),
.B1(n_54),
.B2(n_19),
.Y(n_137)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_73),
.B(n_41),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_53),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_128),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_70),
.B(n_79),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_126),
.A2(n_127),
.B(n_130),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_64),
.B(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_66),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_78),
.B(n_73),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_56),
.B(n_55),
.C(n_84),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_137),
.B1(n_159),
.B2(n_91),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_134),
.B(n_90),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_92),
.B1(n_93),
.B2(n_104),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_41),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_111),
.Y(n_162)
);

XNOR2x1_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_41),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_150),
.C(n_119),
.Y(n_164)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_89),
.A2(n_61),
.A3(n_68),
.B1(n_41),
.B2(n_49),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_128),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_96),
.A2(n_67),
.B1(n_41),
.B2(n_49),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_149),
.A2(n_124),
.B1(n_143),
.B2(n_147),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_68),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_49),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_155),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_49),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_48),
.B1(n_29),
.B2(n_38),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_160),
.A2(n_163),
.B1(n_171),
.B2(n_174),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_161),
.B(n_194),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_162),
.A2(n_176),
.B(n_183),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_110),
.B1(n_123),
.B2(n_100),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_159),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_170),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_167),
.B(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_169),
.B(n_173),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_106),
.B1(n_118),
.B2(n_95),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_130),
.Y(n_175)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_125),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_114),
.B1(n_109),
.B2(n_107),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_182),
.B1(n_191),
.B2(n_192),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_101),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_178),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_122),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_102),
.B1(n_98),
.B2(n_103),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_1),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_131),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_188),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_48),
.C(n_24),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_190),
.C(n_149),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_133),
.B(n_48),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_138),
.B(n_8),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_126),
.B(n_24),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_129),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_24),
.C(n_1),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_140),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_2),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_193),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_154),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_205),
.Y(n_236)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_210),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_171),
.A2(n_136),
.B1(n_144),
.B2(n_124),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_215),
.B1(n_190),
.B2(n_180),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_144),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_216),
.Y(n_229)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_136),
.A3(n_156),
.B1(n_152),
.B2(n_145),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_174),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_213),
.A2(n_219),
.B(n_220),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_187),
.A2(n_143),
.B1(n_157),
.B2(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_146),
.C(n_158),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_222),
.Y(n_230)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_224),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_166),
.B(n_3),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_175),
.A2(n_5),
.B(n_6),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_186),
.C(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

XOR2x2_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_186),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_221),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_232),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_177),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_210),
.C(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_243),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_208),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_168),
.B1(n_162),
.B2(n_176),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_244),
.B1(n_224),
.B2(n_197),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_162),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_241),
.A2(n_214),
.B(n_204),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_226),
.B1(n_248),
.B2(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_197),
.A2(n_176),
.B1(n_192),
.B2(n_170),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_260),
.B(n_264),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_230),
.C(n_231),
.Y(n_269)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_254),
.B(n_258),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_229),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_259),
.A2(n_263),
.B1(n_183),
.B2(n_7),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_262),
.A2(n_241),
.B1(n_195),
.B2(n_212),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_239),
.A2(n_201),
.B1(n_223),
.B2(n_209),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_234),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_200),
.Y(n_265)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_216),
.C(n_205),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_219),
.C(n_183),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_240),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_272),
.C(n_257),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_184),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_230),
.C(n_240),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_282),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_203),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_279),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_242),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_241),
.B1(n_220),
.B2(n_247),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_247),
.B1(n_221),
.B2(n_219),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_283),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_257),
.C(n_249),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_255),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_284),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_294),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_273),
.A2(n_268),
.B(n_265),
.Y(n_292)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_295),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_272),
.C(n_269),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_277),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_250),
.B(n_260),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_297),
.Y(n_303)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_265),
.B(n_259),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_283),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_274),
.B1(n_271),
.B2(n_263),
.Y(n_301)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_292),
.B(n_291),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_308),
.C(n_287),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_306),
.B(n_290),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_279),
.B1(n_285),
.B2(n_278),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_6),
.C(n_7),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_296),
.C(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_288),
.B(n_9),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_10),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_313),
.C(n_316),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_312),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_290),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_318),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_287),
.C(n_291),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_304),
.C(n_307),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_297),
.Y(n_325)
);

A2O1A1O1Ixp25_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_303),
.B(n_297),
.C(n_302),
.D(n_317),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_324),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_326),
.Y(n_327)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_321),
.Y(n_326)
);

AOI21xp33_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_320),
.B(n_322),
.Y(n_329)
);

AOI21xp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_328),
.B(n_12),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_11),
.B(n_12),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_15),
.B(n_16),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_16),
.Y(n_333)
);


endmodule