module real_jpeg_4753_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_1),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_2),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_2),
.A2(n_81),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_2),
.A2(n_81),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_2),
.A2(n_81),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_21),
.B1(n_119),
.B2(n_123),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_38),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_3),
.A2(n_21),
.B1(n_140),
.B2(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_3),
.A2(n_21),
.B1(n_91),
.B2(n_205),
.Y(n_204)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_3),
.A2(n_220),
.B(n_222),
.C(n_228),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_3),
.B(n_102),
.C(n_138),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_3),
.B(n_92),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_3),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_3),
.B(n_106),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_4),
.A2(n_50),
.B1(n_86),
.B2(n_90),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_4),
.A2(n_50),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_4),
.A2(n_50),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_6),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_6),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_6),
.Y(n_279)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_7),
.Y(n_131)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_9),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_9),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_10),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_10),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_208),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_207),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_174),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_16),
.B(n_174),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.C(n_158),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_17),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_52),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_18),
.B(n_53),
.C(n_94),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_47),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B(n_23),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_24),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_21),
.A2(n_223),
.B(n_225),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_23),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_24),
.Y(n_51)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_26),
.B(n_48),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_38),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_38),
.B(n_194),
.Y(n_193)
);

AO22x1_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_45),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g134 ( 
.A(n_39),
.B(n_63),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_93),
.B1(n_94),
.B2(n_124),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_84),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_75),
.Y(n_55)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_56),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_64),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_59),
.Y(n_221)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_60),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_64),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_69),
.B2(n_72),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_68),
.Y(n_227)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_69),
.Y(n_185)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_71),
.Y(n_242)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_76),
.B(n_92),
.Y(n_160)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_83),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_84),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_85),
.B(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_116),
.B(n_117),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_96),
.B(n_118),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_96),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_96),
.B(n_183),
.Y(n_302)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_100),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_106),
.B(n_238),
.Y(n_254)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_112),
.B2(n_114),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_109),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_113),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_116),
.B(n_117),
.Y(n_236)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_125),
.A2(n_126),
.B1(n_158),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_135),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_127),
.B(n_135),
.Y(n_190)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.A3(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_144),
.B(n_147),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_136),
.A2(n_171),
.B(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_146),
.Y(n_288)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_147),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_148),
.A2(n_167),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_148),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx8_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_157),
.Y(n_286)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.C(n_165),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_162),
.B(n_204),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_165),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_166),
.B(n_277),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_167),
.Y(n_258)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_171),
.B(n_260),
.Y(n_291)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_189),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_181),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_182),
.B(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_200),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.Y(n_192)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_243),
.B(n_315),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_211),
.B(n_214),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.C(n_233),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_215),
.B(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_218),
.A2(n_233),
.B1(n_234),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_218),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_230),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_219),
.A2(n_230),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_219),
.Y(n_307)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_230),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_309),
.B(n_314),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_296),
.B(n_308),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_271),
.B(n_295),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_247),
.B(n_255),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_248),
.A2(n_249),
.B1(n_253),
.B2(n_274),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_254),
.B(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_266),
.Y(n_255)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_256),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_268),
.B(n_269),
.C(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_281),
.B(n_294),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_280),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_290),
.B(n_293),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_289),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_299),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_303),
.C(n_305),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_313),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_313),
.Y(n_314)
);


endmodule