module fake_ariane_324_n_2164 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2164);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2164;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_279;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1661;
wire n_1468;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g216 ( 
.A(n_84),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_81),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_82),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_174),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_77),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_16),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_167),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_173),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_166),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_177),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_72),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_175),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_88),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_103),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_160),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_16),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_95),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_170),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_80),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_187),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_113),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_32),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_142),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_114),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_69),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_111),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_20),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_129),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_119),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_76),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_85),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_29),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_74),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_180),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_96),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_91),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_46),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_87),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_69),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_20),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_185),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_30),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_53),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_26),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_46),
.Y(n_264)
);

INVxp33_ASAP7_75t_R g265 ( 
.A(n_26),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_55),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_72),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_188),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_24),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_144),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_78),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_105),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_50),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_106),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_17),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_145),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_162),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_90),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_99),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_183),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_156),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_94),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_133),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_211),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_135),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_11),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_39),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_147),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_38),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_169),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_30),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_65),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_42),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_51),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_40),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_22),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_39),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_13),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_3),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_203),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_112),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_23),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_5),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_75),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_168),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_140),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_18),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_62),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_98),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_92),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_97),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_24),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_40),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_146),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_4),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_35),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_163),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_60),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_190),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_209),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_212),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_120),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_6),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_107),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_213),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_89),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_50),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_206),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_125),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_131),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_172),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_121),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_198),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_71),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_6),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_9),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_34),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_60),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_136),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_12),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_194),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_53),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_110),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_184),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_47),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_15),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_55),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_31),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_137),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_155),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_49),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_148),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_61),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_122),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_83),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_178),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_31),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_61),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_51),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_42),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_118),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_152),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_36),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_150),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_4),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_12),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_38),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_8),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_195),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_9),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_10),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_191),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_201),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_67),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_28),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_33),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_54),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_205),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_65),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_27),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_179),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_70),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_71),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_176),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_109),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_124),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_1),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_197),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_86),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_123),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_23),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_202),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_93),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_153),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_130),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_132),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_34),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_68),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_14),
.Y(n_400)
);

CKINVDCx11_ASAP7_75t_R g401 ( 
.A(n_48),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_127),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_32),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_47),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_186),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_64),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_57),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_116),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_70),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_108),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_104),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_2),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_126),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_161),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_101),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_18),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_2),
.Y(n_417)
);

BUFx10_ASAP7_75t_L g418 ( 
.A(n_199),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_193),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_15),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_157),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_79),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_8),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_21),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_58),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_324),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_275),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_275),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_343),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_343),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_392),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_401),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_392),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_287),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_388),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_278),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_307),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_388),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_278),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_243),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_344),
.Y(n_443)
);

BUFx6f_ASAP7_75t_SL g444 ( 
.A(n_396),
.Y(n_444)
);

BUFx2_ASAP7_75t_SL g445 ( 
.A(n_396),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_246),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_216),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_355),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_368),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_370),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_368),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_243),
.B(n_0),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_373),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_216),
.B(n_0),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_391),
.Y(n_456)
);

BUFx6f_ASAP7_75t_SL g457 ( 
.A(n_396),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_379),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_R g459 ( 
.A(n_220),
.B(n_73),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_379),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_217),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_232),
.B(n_1),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_246),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_251),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_251),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_261),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_419),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_402),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_402),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_261),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_217),
.B(n_3),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_L g473 ( 
.A(n_232),
.B(n_5),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_227),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_262),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_219),
.B(n_7),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_241),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_262),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_276),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_396),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_267),
.B(n_7),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_244),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_418),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_418),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_276),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_290),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_418),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_267),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_219),
.B(n_10),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_290),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_418),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_296),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_233),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_328),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_256),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_258),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_259),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_296),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_233),
.B(n_13),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_303),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_264),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_266),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_269),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_303),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_240),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_274),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_335),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_328),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_328),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_335),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_288),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_300),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_293),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_337),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_240),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_313),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_248),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_295),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_248),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_328),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_297),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_398),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_298),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_328),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_318),
.B(n_14),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_299),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_260),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_304),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_317),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_260),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_308),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_270),
.Y(n_532)
);

NOR2xp67_ASAP7_75t_L g533 ( 
.A(n_292),
.B(n_17),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_270),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_272),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_398),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_309),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_337),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_292),
.B(n_19),
.Y(n_539)
);

NOR2xp67_ASAP7_75t_L g540 ( 
.A(n_294),
.B(n_19),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_445),
.B(n_480),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_439),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_443),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_512),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_494),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_516),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_447),
.B(n_294),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_445),
.B(n_398),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_448),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_494),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_483),
.B(n_332),
.Y(n_552)
);

CKINVDCx8_ASAP7_75t_R g553 ( 
.A(n_449),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_450),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_453),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_456),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_520),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_483),
.B(n_284),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_509),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_509),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_467),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_447),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_436),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_524),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_433),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_484),
.B(n_284),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_529),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_495),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_461),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_SL g572 ( 
.A(n_428),
.B(n_360),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_488),
.B(n_398),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_428),
.B(n_399),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_484),
.B(n_291),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_493),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_493),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_487),
.B(n_291),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_505),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_505),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_522),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_515),
.B(n_238),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_487),
.B(n_306),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_495),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g585 ( 
.A(n_429),
.B(n_265),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_496),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_496),
.Y(n_587)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_536),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_429),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_515),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_444),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_517),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_R g593 ( 
.A(n_491),
.B(n_221),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_517),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_451),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_488),
.B(n_354),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g597 ( 
.A(n_444),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_497),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_519),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_497),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_519),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_527),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_527),
.A2(n_310),
.B(n_306),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_530),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_532),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_532),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_534),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_534),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_535),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_437),
.B(n_354),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_438),
.B(n_265),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_474),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_491),
.B(n_223),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_502),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_535),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_463),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_427),
.B(n_359),
.Y(n_618)
);

OA21x2_ASAP7_75t_L g619 ( 
.A1(n_454),
.A2(n_322),
.B(n_310),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_502),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_464),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_438),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_465),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_466),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_441),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_455),
.B(n_222),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_475),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_441),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_472),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_440),
.B(n_359),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_549),
.B(n_455),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_541),
.B(n_477),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_549),
.B(n_430),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_564),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_582),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_559),
.B(n_458),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_593),
.B(n_458),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_571),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_560),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_571),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_571),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_545),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_571),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

NOR2x1p5_ASAP7_75t_L g645 ( 
.A(n_570),
.B(n_460),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_571),
.Y(n_646)
);

BUFx10_ASAP7_75t_L g647 ( 
.A(n_552),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_547),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_555),
.B(n_468),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_555),
.B(n_468),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_560),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_561),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_576),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_576),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_SL g655 ( 
.A(n_553),
.B(n_469),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_576),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_576),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_576),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_561),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_558),
.B(n_469),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_582),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_558),
.B(n_431),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_565),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_567),
.B(n_444),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_576),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_569),
.Y(n_666)
);

AND2x2_ASAP7_75t_SL g667 ( 
.A(n_597),
.B(n_452),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_565),
.B(n_575),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_561),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_569),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_561),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_569),
.Y(n_672)
);

INVxp33_ASAP7_75t_L g673 ( 
.A(n_585),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_569),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_582),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_546),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_546),
.Y(n_677)
);

NAND2xp33_ASAP7_75t_L g678 ( 
.A(n_582),
.B(n_525),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_544),
.B(n_462),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_609),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_546),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_609),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_609),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_578),
.B(n_432),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_609),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_573),
.B(n_434),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_582),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_577),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_582),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_596),
.B(n_446),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_553),
.B(n_457),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_563),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_573),
.B(n_435),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_563),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_546),
.Y(n_695)
);

XNOR2xp5_ASAP7_75t_L g696 ( 
.A(n_585),
.B(n_503),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_548),
.B(n_478),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_583),
.B(n_503),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_546),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_584),
.B(n_506),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_563),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_546),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_603),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_604),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_591),
.B(n_506),
.Y(n_705)
);

NOR2x1p5_ASAP7_75t_L g706 ( 
.A(n_586),
.B(n_513),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_551),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_591),
.B(n_513),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_604),
.Y(n_709)
);

AND2x2_ASAP7_75t_SL g710 ( 
.A(n_597),
.B(n_471),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_582),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_551),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_591),
.B(n_577),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_591),
.B(n_580),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_614),
.B(n_457),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_548),
.B(n_624),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_587),
.B(n_518),
.Y(n_717)
);

BUFx4f_ASAP7_75t_L g718 ( 
.A(n_619),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_604),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_606),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_551),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_606),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_596),
.B(n_470),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_589),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_606),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_551),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_548),
.B(n_479),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_551),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_551),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_548),
.B(n_507),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_580),
.B(n_518),
.Y(n_731)
);

INVx4_ASAP7_75t_L g732 ( 
.A(n_617),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_590),
.B(n_592),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_590),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_598),
.B(n_521),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_579),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_600),
.B(n_521),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_618),
.B(n_473),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_592),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_594),
.B(n_599),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_613),
.B(n_457),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_594),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_579),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_599),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_601),
.B(n_523),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_601),
.B(n_523),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_608),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_615),
.B(n_620),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_608),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_603),
.Y(n_750)
);

INVx5_ASAP7_75t_L g751 ( 
.A(n_617),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_624),
.B(n_627),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_619),
.A2(n_476),
.B1(n_499),
.B2(n_489),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_602),
.B(n_605),
.Y(n_754)
);

INVx4_ASAP7_75t_SL g755 ( 
.A(n_602),
.Y(n_755)
);

AND2x2_ASAP7_75t_SL g756 ( 
.A(n_619),
.B(n_588),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_605),
.B(n_528),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_626),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_568),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_607),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_610),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_607),
.B(n_528),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_617),
.B(n_537),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_610),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_617),
.B(n_537),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_616),
.B(n_442),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_616),
.B(n_482),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_621),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_627),
.Y(n_769)
);

INVxp33_ASAP7_75t_L g770 ( 
.A(n_612),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_619),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_542),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_621),
.B(n_501),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_623),
.Y(n_774)
);

AND2x6_ASAP7_75t_L g775 ( 
.A(n_623),
.B(n_322),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_618),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_618),
.A2(n_540),
.B1(n_533),
.B2(n_539),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_588),
.B(n_511),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_595),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_618),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_572),
.A2(n_459),
.B1(n_339),
.B2(n_341),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_626),
.B(n_526),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_611),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_629),
.B(n_328),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_611),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_664),
.B(n_531),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_688),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_698),
.B(n_630),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_727),
.B(n_730),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_755),
.Y(n_790)
);

OR2x6_ASAP7_75t_L g791 ( 
.A(n_634),
.B(n_630),
.Y(n_791)
);

BUFx8_ASAP7_75t_L g792 ( 
.A(n_724),
.Y(n_792)
);

NAND2x1_ASAP7_75t_L g793 ( 
.A(n_635),
.B(n_675),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_739),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_668),
.B(n_253),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_753),
.A2(n_314),
.B1(n_319),
.B2(n_316),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_772),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_761),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_761),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_761),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_761),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_636),
.A2(n_336),
.B1(n_347),
.B2(n_346),
.Y(n_802)
);

AND2x2_ASAP7_75t_SL g803 ( 
.A(n_756),
.B(n_678),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_632),
.B(n_254),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_633),
.B(n_745),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_734),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_635),
.B(n_345),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_756),
.A2(n_625),
.B1(n_628),
.B2(n_622),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_635),
.B(n_345),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_734),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_761),
.Y(n_811)
);

INVx8_ASAP7_75t_L g812 ( 
.A(n_775),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_633),
.B(n_273),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_718),
.A2(n_481),
.B(n_356),
.C(n_362),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_639),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_746),
.B(n_408),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_731),
.A2(n_338),
.B(n_377),
.C(n_371),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_757),
.B(n_369),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_651),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_742),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_675),
.B(n_350),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_763),
.B(n_263),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_765),
.B(n_366),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_684),
.B(n_369),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_758),
.B(n_543),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_758),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_631),
.B(n_348),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_768),
.B(n_416),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_631),
.B(n_349),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_642),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_742),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_663),
.B(n_350),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_722),
.Y(n_833)
);

BUFx5_ASAP7_75t_L g834 ( 
.A(n_666),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_663),
.B(n_356),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_752),
.B(n_362),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_752),
.B(n_363),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_670),
.B(n_363),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_741),
.B(n_550),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_762),
.A2(n_760),
.B1(n_744),
.B2(n_708),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_670),
.B(n_365),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_R g842 ( 
.A(n_772),
.B(n_554),
.Y(n_842)
);

NOR3xp33_ASAP7_75t_L g843 ( 
.A(n_700),
.B(n_358),
.C(n_352),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_670),
.B(n_365),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_683),
.B(n_393),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_647),
.B(n_361),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_683),
.B(n_393),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_683),
.B(n_774),
.Y(n_848)
);

INVxp67_ASAP7_75t_L g849 ( 
.A(n_779),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_648),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_744),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_675),
.B(n_422),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_687),
.B(n_422),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_760),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_687),
.B(n_689),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_652),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_649),
.B(n_364),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_774),
.B(n_338),
.Y(n_858)
);

OAI221xp5_ASAP7_75t_L g859 ( 
.A1(n_781),
.A2(n_412),
.B1(n_377),
.B2(n_378),
.C(n_371),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_718),
.A2(n_286),
.B(n_223),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_716),
.B(n_783),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_716),
.B(n_783),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_666),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_732),
.B(n_378),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_L g865 ( 
.A(n_750),
.B(n_367),
.Y(n_865)
);

NAND2xp33_ASAP7_75t_L g866 ( 
.A(n_750),
.B(n_367),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_732),
.B(n_406),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_690),
.B(n_574),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_732),
.B(n_406),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_652),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_647),
.B(n_372),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_672),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_650),
.B(n_375),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_690),
.B(n_574),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_705),
.A2(n_407),
.B1(n_384),
.B2(n_383),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_678),
.A2(n_581),
.B1(n_311),
.B2(n_286),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_724),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_660),
.B(n_376),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_715),
.A2(n_311),
.B1(n_331),
.B2(n_330),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_771),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_686),
.B(n_409),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_647),
.B(n_767),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_686),
.B(n_409),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_693),
.B(n_412),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_693),
.B(n_776),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_L g886 ( 
.A(n_717),
.B(n_737),
.C(n_735),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_723),
.B(n_612),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_672),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_674),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_723),
.B(n_556),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_710),
.A2(n_252),
.B1(n_305),
.B2(n_302),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_723),
.B(n_557),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_773),
.B(n_380),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_776),
.B(n_420),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_674),
.Y(n_895)
);

O2A1O1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_733),
.A2(n_420),
.B(n_514),
.C(n_485),
.Y(n_896)
);

AOI221xp5_ASAP7_75t_L g897 ( 
.A1(n_782),
.A2(n_404),
.B1(n_400),
.B2(n_417),
.C(n_423),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_750),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_659),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_680),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_780),
.B(n_403),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_687),
.B(n_218),
.Y(n_902)
);

O2A1O1Ixp5_ASAP7_75t_L g903 ( 
.A1(n_703),
.A2(n_538),
.B(n_510),
.C(n_504),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_785),
.B(n_486),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_689),
.B(n_218),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_727),
.Y(n_906)
);

NAND3xp33_ASAP7_75t_L g907 ( 
.A(n_748),
.B(n_425),
.C(n_424),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_710),
.A2(n_237),
.B1(n_255),
.B2(n_250),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_659),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_759),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_718),
.A2(n_280),
.B(n_245),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_689),
.B(n_245),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_785),
.B(n_490),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_646),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_730),
.B(n_749),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_730),
.B(n_562),
.Y(n_916)
);

NAND2xp33_ASAP7_75t_L g917 ( 
.A(n_750),
.B(n_367),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_780),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_637),
.B(n_566),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_749),
.B(n_492),
.Y(n_920)
);

NAND2x1_ASAP7_75t_L g921 ( 
.A(n_711),
.B(n_242),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_749),
.B(n_740),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_655),
.B(n_498),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_680),
.A2(n_353),
.B(n_280),
.C(n_390),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_754),
.B(n_500),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_713),
.A2(n_367),
.B1(n_390),
.B2(n_387),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_667),
.B(n_224),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_682),
.B(n_225),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_775),
.A2(n_230),
.B1(n_415),
.B2(n_414),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_775),
.A2(n_421),
.B1(n_238),
.B2(n_334),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_697),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_775),
.A2(n_229),
.B1(n_413),
.B2(n_411),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_682),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_697),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_SL g935 ( 
.A(n_706),
.B(n_367),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_738),
.B(n_21),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_685),
.B(n_226),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_711),
.B(n_312),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_685),
.B(n_228),
.Y(n_939)
);

AO22x1_ASAP7_75t_L g940 ( 
.A1(n_775),
.A2(n_312),
.B1(n_387),
.B2(n_386),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_669),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_679),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_784),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_711),
.B(n_323),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_738),
.B(n_22),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_775),
.A2(n_315),
.B1(n_410),
.B2(n_405),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_825),
.B(n_696),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_840),
.A2(n_714),
.B(n_750),
.Y(n_948)
);

BUFx2_ASAP7_75t_SL g949 ( 
.A(n_830),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_788),
.B(n_667),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_833),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_804),
.A2(n_738),
.B1(n_784),
.B2(n_645),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_789),
.B(n_691),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_882),
.B(n_778),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_882),
.B(n_673),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_910),
.B(n_770),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_880),
.A2(n_848),
.B(n_865),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_880),
.A2(n_641),
.B(n_640),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_806),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_866),
.A2(n_641),
.B(n_640),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_788),
.B(n_662),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_917),
.A2(n_644),
.B(n_643),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_810),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_805),
.B(n_738),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_903),
.A2(n_771),
.B(n_677),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_820),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_910),
.B(n_696),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_877),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_890),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_898),
.A2(n_771),
.B(n_644),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_831),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_816),
.A2(n_751),
.B1(n_638),
.B2(n_692),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_898),
.A2(n_922),
.B(n_855),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_898),
.A2(n_653),
.B(n_643),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_795),
.B(n_769),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_898),
.A2(n_654),
.B(n_653),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_792),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_822),
.A2(n_704),
.B(n_719),
.C(n_720),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_851),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_822),
.B(n_823),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_815),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_789),
.B(n_751),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_823),
.B(n_769),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_855),
.A2(n_656),
.B(n_654),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_892),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_790),
.Y(n_986)
);

CKINVDCx10_ASAP7_75t_R g987 ( 
.A(n_842),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_826),
.B(n_751),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_854),
.A2(n_751),
.B1(n_638),
.B2(n_725),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_797),
.Y(n_990)
);

O2A1O1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_796),
.A2(n_766),
.B(n_701),
.C(n_704),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_857),
.A2(n_679),
.B1(n_638),
.B2(n_751),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_861),
.Y(n_993)
);

INVx5_ASAP7_75t_L g994 ( 
.A(n_812),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_857),
.B(n_736),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_911),
.A2(n_657),
.B(n_656),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_864),
.A2(n_869),
.B(n_867),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_838),
.A2(n_844),
.B(n_841),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_873),
.B(n_736),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_845),
.A2(n_658),
.B(n_657),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_860),
.A2(n_694),
.B(n_692),
.Y(n_1001)
);

NOR2x1p5_ASAP7_75t_L g1002 ( 
.A(n_868),
.B(n_679),
.Y(n_1002)
);

NAND3xp33_ASAP7_75t_L g1003 ( 
.A(n_849),
.B(n_701),
.C(n_694),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_802),
.A2(n_720),
.B(n_709),
.C(n_719),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_873),
.B(n_743),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_847),
.A2(n_658),
.B(n_665),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_878),
.B(n_743),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_862),
.Y(n_1008)
);

AO21x1_ASAP7_75t_L g1009 ( 
.A1(n_818),
.A2(n_709),
.B(n_725),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_849),
.B(n_679),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_SL g1011 ( 
.A(n_850),
.B(n_661),
.Y(n_1011)
);

AOI22x1_ASAP7_75t_L g1012 ( 
.A1(n_863),
.A2(n_665),
.B1(n_764),
.B2(n_747),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_878),
.B(n_747),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_893),
.B(n_931),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_872),
.A2(n_729),
.B(n_726),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_893),
.A2(n_931),
.B(n_827),
.C(n_829),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_790),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_819),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_885),
.B(n_764),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_906),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_888),
.A2(n_729),
.B(n_676),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_803),
.A2(n_906),
.B1(n_915),
.B2(n_787),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_889),
.A2(n_729),
.B(n_676),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_895),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_813),
.B(n_777),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_900),
.A2(n_661),
.B(n_728),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_786),
.B(n_755),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_897),
.B(n_671),
.C(n_646),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_933),
.A2(n_661),
.B(n_726),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_918),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_936),
.A2(n_671),
.B(n_721),
.C(n_712),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_814),
.A2(n_905),
.B(n_902),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_856),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_925),
.B(n_646),
.Y(n_1034)
);

INVx5_ASAP7_75t_L g1035 ( 
.A(n_812),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_928),
.A2(n_728),
.B(n_721),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_870),
.Y(n_1037)
);

BUFx4f_ASAP7_75t_L g1038 ( 
.A(n_791),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_918),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_920),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_850),
.B(n_646),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_937),
.A2(n_712),
.B(n_707),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_936),
.A2(n_707),
.B(n_702),
.C(n_677),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_923),
.B(n_646),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_L g1045 ( 
.A1(n_858),
.A2(n_702),
.B(n_681),
.C(n_323),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_SL g1046 ( 
.A(n_874),
.B(n_887),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_945),
.A2(n_681),
.B(n_353),
.C(n_386),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_939),
.A2(n_699),
.B(n_695),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_902),
.A2(n_912),
.B(n_905),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_934),
.B(n_695),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_901),
.B(n_695),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_914),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_803),
.A2(n_367),
.B1(n_695),
.B2(n_699),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_901),
.B(n_695),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_793),
.A2(n_699),
.B(n_289),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_938),
.A2(n_421),
.B(n_334),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_824),
.B(n_231),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_808),
.B(n_234),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_876),
.B(n_235),
.Y(n_1059)
);

AO21x1_ASAP7_75t_L g1060 ( 
.A1(n_944),
.A2(n_421),
.B(n_334),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_SL g1061 ( 
.A(n_792),
.B(n_839),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_914),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_927),
.B(n_236),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_899),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_945),
.A2(n_238),
.B(n_395),
.C(n_394),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_891),
.B(n_239),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_894),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_812),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_842),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_791),
.B(n_25),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_908),
.B(n_397),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_904),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_944),
.A2(n_389),
.B(n_385),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_879),
.B(n_382),
.C(n_374),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_913),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_794),
.B(n_247),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_791),
.B(n_249),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_914),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_943),
.A2(n_357),
.B(n_351),
.C(n_342),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_SL g1080 ( 
.A(n_942),
.Y(n_1080)
);

AO21x2_ASAP7_75t_L g1081 ( 
.A1(n_832),
.A2(n_242),
.B(n_149),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_807),
.A2(n_340),
.B(n_333),
.Y(n_1082)
);

AOI21x1_ASAP7_75t_L g1083 ( 
.A1(n_807),
.A2(n_242),
.B(n_327),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_809),
.A2(n_329),
.B(n_326),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_809),
.A2(n_325),
.B(n_321),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_821),
.A2(n_320),
.B(n_301),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_821),
.A2(n_285),
.B(n_283),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_828),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_909),
.A2(n_282),
.B(n_281),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_852),
.A2(n_279),
.B(n_277),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_886),
.B(n_271),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_817),
.A2(n_268),
.B(n_257),
.C(n_242),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_852),
.A2(n_242),
.B(n_102),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_941),
.Y(n_1094)
);

CKINVDCx6p67_ASAP7_75t_R g1095 ( 
.A(n_916),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_835),
.B(n_25),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_836),
.B(n_27),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_837),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_881),
.B(n_28),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_853),
.A2(n_242),
.B(n_115),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_935),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_883),
.B(n_29),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_884),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_875),
.B(n_33),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_846),
.B(n_35),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_896),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_853),
.A2(n_128),
.B(n_214),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_834),
.B(n_36),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_834),
.B(n_37),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_921),
.A2(n_798),
.B(n_799),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_843),
.B(n_37),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_800),
.A2(n_134),
.B(n_210),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_801),
.A2(n_41),
.B(n_43),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_914),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_811),
.A2(n_117),
.B(n_208),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_871),
.A2(n_41),
.B(n_43),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_929),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_907),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_843),
.B(n_44),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_924),
.A2(n_44),
.B(n_45),
.Y(n_1120)
);

AOI21x1_ASAP7_75t_L g1121 ( 
.A1(n_926),
.A2(n_138),
.B(n_207),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_834),
.B(n_45),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_859),
.B(n_48),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_940),
.A2(n_49),
.B(n_52),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_834),
.B(n_52),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_980),
.B(n_919),
.Y(n_1126)
);

INVx4_ASAP7_75t_L g1127 ( 
.A(n_994),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1123),
.A2(n_1105),
.B(n_954),
.C(n_1014),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1062),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_959),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1066),
.A2(n_930),
.B(n_932),
.C(n_946),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1068),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_955),
.B(n_834),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_948),
.A2(n_930),
.B(n_834),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_948),
.A2(n_54),
.B(n_56),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_957),
.A2(n_997),
.B(n_958),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_L g1137 ( 
.A(n_1071),
.B(n_56),
.C(n_57),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_963),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_961),
.B(n_58),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_965),
.A2(n_143),
.B(n_204),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_968),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_SL g1142 ( 
.A(n_1104),
.B(n_952),
.C(n_1116),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_997),
.A2(n_59),
.B(n_62),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1072),
.B(n_59),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_957),
.A2(n_63),
.B(n_64),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_958),
.A2(n_978),
.B(n_998),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_990),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_998),
.A2(n_63),
.B(n_66),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_950),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_987),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1075),
.B(n_139),
.Y(n_1151)
);

O2A1O1Ixp5_ASAP7_75t_L g1152 ( 
.A1(n_1009),
.A2(n_1048),
.B(n_972),
.C(n_1122),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1068),
.Y(n_1153)
);

INVxp67_ASAP7_75t_SL g1154 ( 
.A(n_1044),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1036),
.A2(n_141),
.B(n_151),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1103),
.B(n_993),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_1069),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1008),
.B(n_154),
.Y(n_1158)
);

OAI222xp33_ASAP7_75t_L g1159 ( 
.A1(n_947),
.A2(n_159),
.B1(n_164),
.B2(n_165),
.C1(n_171),
.C2(n_182),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1036),
.A2(n_192),
.B(n_196),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_994),
.B(n_215),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1042),
.A2(n_1021),
.B(n_1015),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_995),
.A2(n_1005),
.B(n_999),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1007),
.A2(n_1013),
.B(n_1051),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_994),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1083),
.A2(n_996),
.B(n_1053),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1098),
.A2(n_1016),
.B(n_1102),
.C(n_1099),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1054),
.A2(n_1042),
.B(n_970),
.Y(n_1168)
);

NAND2xp33_ASAP7_75t_SL g1169 ( 
.A(n_964),
.B(n_1118),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1025),
.B(n_1067),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1015),
.A2(n_1023),
.B(n_1021),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_SL g1172 ( 
.A1(n_1108),
.A2(n_1125),
.B(n_1109),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1034),
.A2(n_1023),
.B(n_1006),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_994),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_973),
.A2(n_1056),
.B(n_1012),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1062),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_996),
.A2(n_1006),
.B(n_1000),
.Y(n_1177)
);

AOI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1058),
.A2(n_967),
.B(n_956),
.Y(n_1178)
);

NOR2xp67_ASAP7_75t_L g1179 ( 
.A(n_977),
.B(n_1010),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1035),
.B(n_1002),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1060),
.A2(n_1000),
.B(n_960),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_985),
.B(n_969),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_L g1183 ( 
.A(n_1116),
.B(n_1065),
.C(n_1119),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_981),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_SL g1185 ( 
.A1(n_1097),
.A2(n_1096),
.B(n_1027),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1020),
.B(n_966),
.Y(n_1186)
);

INVx6_ASAP7_75t_SL g1187 ( 
.A(n_949),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1038),
.B(n_1046),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1022),
.A2(n_1043),
.A3(n_1031),
.B(n_1047),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1038),
.B(n_1070),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_960),
.A2(n_962),
.B(n_1045),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_962),
.A2(n_1001),
.B(n_984),
.Y(n_1192)
);

CKINVDCx6p67_ASAP7_75t_R g1193 ( 
.A(n_1080),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_991),
.A2(n_1004),
.B(n_1028),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_971),
.Y(n_1195)
);

O2A1O1Ixp5_ASAP7_75t_L g1196 ( 
.A1(n_1032),
.A2(n_1106),
.B(n_989),
.C(n_1107),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_974),
.A2(n_976),
.B(n_983),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_1035),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1003),
.A2(n_1040),
.B(n_1110),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1095),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1024),
.A2(n_1073),
.B(n_951),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1117),
.B(n_1030),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1049),
.A2(n_1115),
.B(n_1029),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1121),
.A2(n_975),
.B(n_1019),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1026),
.A2(n_1112),
.B(n_1055),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1093),
.A2(n_1100),
.B(n_1052),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_979),
.B(n_1041),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1124),
.A2(n_1113),
.B(n_1091),
.C(n_1111),
.Y(n_1208)
);

AOI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1063),
.A2(n_1077),
.B(n_1074),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1124),
.A2(n_1113),
.B(n_1120),
.C(n_992),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1062),
.B(n_1114),
.Y(n_1211)
);

OR2x2_ASAP7_75t_L g1212 ( 
.A(n_1039),
.B(n_953),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1035),
.A2(n_1050),
.B1(n_1057),
.B2(n_1076),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_988),
.A2(n_1089),
.B(n_1088),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1052),
.A2(n_982),
.B(n_1059),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1018),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1094),
.B(n_1037),
.Y(n_1217)
);

INVx5_ASAP7_75t_L g1218 ( 
.A(n_1035),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_SL g1219 ( 
.A1(n_1120),
.A2(n_1085),
.B(n_1084),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1079),
.A2(n_1086),
.B(n_1085),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1092),
.A2(n_1084),
.B(n_1082),
.C(n_1086),
.Y(n_1221)
);

INVx3_ASAP7_75t_SL g1222 ( 
.A(n_1078),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_L g1223 ( 
.A(n_986),
.B(n_1017),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1033),
.B(n_1064),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1078),
.A2(n_1114),
.B(n_1087),
.Y(n_1225)
);

AND2x2_ASAP7_75t_SL g1226 ( 
.A(n_1061),
.B(n_1011),
.Y(n_1226)
);

NOR2xp67_ASAP7_75t_SL g1227 ( 
.A(n_1078),
.B(n_1114),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1082),
.A2(n_1101),
.B(n_1081),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1081),
.A2(n_986),
.B(n_1017),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1090),
.A2(n_965),
.B(n_1048),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1080),
.A2(n_948),
.B(n_898),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_959),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_994),
.B(n_789),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_980),
.A2(n_948),
.B(n_957),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_980),
.A2(n_948),
.B(n_957),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_948),
.A2(n_898),
.B(n_997),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_948),
.A2(n_898),
.B(n_997),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1022),
.B(n_803),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_965),
.A2(n_1048),
.B(n_1042),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_965),
.A2(n_1048),
.B(n_1042),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1069),
.B(n_772),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1009),
.A2(n_1060),
.A3(n_1022),
.B(n_1043),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_965),
.A2(n_1048),
.B(n_1042),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_981),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1009),
.A2(n_1060),
.A3(n_1022),
.B(n_1043),
.Y(n_1245)
);

AOI21xp33_ASAP7_75t_L g1246 ( 
.A1(n_980),
.A2(n_1071),
.B(n_1066),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_980),
.B(n_805),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_980),
.A2(n_948),
.B(n_957),
.Y(n_1248)
);

OAI21xp33_ASAP7_75t_SL g1249 ( 
.A1(n_980),
.A2(n_1014),
.B(n_803),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_980),
.B(n_805),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_980),
.B(n_805),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_980),
.B(n_805),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_980),
.B(n_805),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_965),
.A2(n_1048),
.B(n_1042),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1062),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_987),
.Y(n_1256)
);

AOI21xp33_ASAP7_75t_L g1257 ( 
.A1(n_980),
.A2(n_1071),
.B(n_1066),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_965),
.A2(n_1048),
.B(n_1042),
.Y(n_1258)
);

BUFx12f_ASAP7_75t_L g1259 ( 
.A(n_977),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_981),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_965),
.A2(n_1048),
.B(n_1042),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_965),
.A2(n_1048),
.B(n_1042),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_981),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_967),
.B(n_758),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_981),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_980),
.B(n_805),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_980),
.A2(n_948),
.B(n_957),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_987),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_965),
.A2(n_1048),
.B(n_1042),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_968),
.Y(n_1270)
);

AND2x2_ASAP7_75t_SL g1271 ( 
.A(n_1038),
.B(n_803),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1022),
.B(n_803),
.Y(n_1272)
);

OAI21xp33_ASAP7_75t_L g1273 ( 
.A1(n_980),
.A2(n_893),
.B(n_584),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1062),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1048),
.A2(n_911),
.B(n_948),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1069),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_980),
.A2(n_948),
.B(n_957),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1009),
.A2(n_1060),
.A3(n_1022),
.B(n_1043),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_948),
.A2(n_898),
.B(n_997),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_965),
.A2(n_1048),
.B(n_1042),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1022),
.B(n_803),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_987),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1123),
.A2(n_803),
.B1(n_980),
.B2(n_756),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_980),
.A2(n_1123),
.B(n_1105),
.C(n_954),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1256),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1147),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1133),
.B(n_1247),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1200),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1276),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1222),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1182),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1186),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1141),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1222),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1264),
.B(n_1202),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_1268),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1202),
.B(n_1250),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1212),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1246),
.A2(n_1257),
.B1(n_1273),
.B2(n_1284),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1133),
.B(n_1251),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1252),
.B(n_1253),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1190),
.B(n_1178),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1180),
.B(n_1233),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1284),
.A2(n_1128),
.B1(n_1283),
.B2(n_1266),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1188),
.B(n_1128),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1180),
.B(n_1233),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1236),
.A2(n_1279),
.B(n_1237),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1216),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1130),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1283),
.A2(n_1139),
.B1(n_1131),
.B2(n_1135),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1129),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1241),
.B(n_1126),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1187),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1138),
.Y(n_1314)
);

AO32x1_ASAP7_75t_L g1315 ( 
.A1(n_1149),
.A2(n_1213),
.A3(n_1232),
.B1(n_1195),
.B2(n_1185),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1157),
.B(n_1271),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1271),
.B(n_1270),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1156),
.B(n_1150),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_1259),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1244),
.Y(n_1320)
);

INVx5_ASAP7_75t_L g1321 ( 
.A(n_1198),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1161),
.B(n_1179),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1129),
.Y(n_1323)
);

OAI22x1_ASAP7_75t_L g1324 ( 
.A1(n_1137),
.A2(n_1183),
.B1(n_1281),
.B2(n_1272),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1260),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1226),
.B(n_1209),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1129),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1234),
.A2(n_1235),
.B(n_1248),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1282),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1263),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1129),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1169),
.A2(n_1226),
.B1(n_1142),
.B2(n_1249),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1236),
.A2(n_1237),
.B(n_1279),
.Y(n_1333)
);

NAND2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1198),
.B(n_1218),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1142),
.A2(n_1281),
.B1(n_1272),
.B2(n_1238),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1193),
.Y(n_1336)
);

INVx5_ASAP7_75t_L g1337 ( 
.A(n_1198),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1170),
.B(n_1207),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1208),
.A2(n_1167),
.B(n_1196),
.C(n_1214),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1176),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1187),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1265),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1176),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1144),
.B(n_1217),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_SL g1345 ( 
.A(n_1159),
.B(n_1218),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1224),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1201),
.B(n_1176),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1136),
.A2(n_1277),
.B(n_1267),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1154),
.B(n_1163),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1127),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1238),
.B(n_1167),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1132),
.B(n_1153),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1143),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1164),
.B(n_1214),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1151),
.B(n_1158),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1176),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1164),
.B(n_1208),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1134),
.A2(n_1146),
.B(n_1172),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1143),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1255),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1199),
.B(n_1223),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1192),
.A2(n_1173),
.B(n_1168),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1161),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1153),
.B(n_1174),
.Y(n_1365)
);

AOI21xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1211),
.A2(n_1220),
.B(n_1219),
.Y(n_1366)
);

INVx4_ASAP7_75t_L g1367 ( 
.A(n_1255),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1255),
.B(n_1274),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1255),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1274),
.Y(n_1370)
);

INVxp67_ASAP7_75t_SL g1371 ( 
.A(n_1227),
.Y(n_1371)
);

BUFx12f_ASAP7_75t_L g1372 ( 
.A(n_1274),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1148),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1165),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1274),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1210),
.A2(n_1194),
.B(n_1196),
.C(n_1148),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1165),
.B(n_1174),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1215),
.B(n_1210),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1211),
.B(n_1159),
.Y(n_1379)
);

AND2x2_ASAP7_75t_SL g1380 ( 
.A(n_1275),
.B(n_1145),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1145),
.A2(n_1221),
.B1(n_1192),
.B2(n_1215),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1177),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1173),
.A2(n_1168),
.B(n_1197),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1175),
.A2(n_1230),
.B(n_1269),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1171),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1189),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1231),
.B(n_1197),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1221),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1231),
.B(n_1242),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1229),
.A2(n_1152),
.B(n_1275),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1242),
.B(n_1278),
.Y(n_1391)
);

NOR2xp67_ASAP7_75t_L g1392 ( 
.A(n_1225),
.B(n_1228),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1152),
.A2(n_1228),
.B(n_1225),
.C(n_1229),
.Y(n_1393)
);

BUFx4f_ASAP7_75t_L g1394 ( 
.A(n_1185),
.Y(n_1394)
);

NOR2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1204),
.B(n_1181),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1245),
.B(n_1278),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1206),
.B(n_1278),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1245),
.B(n_1278),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1155),
.Y(n_1399)
);

CKINVDCx8_ASAP7_75t_R g1400 ( 
.A(n_1245),
.Y(n_1400)
);

CKINVDCx16_ASAP7_75t_R g1401 ( 
.A(n_1160),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1140),
.B(n_1166),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1162),
.A2(n_1191),
.B1(n_1205),
.B2(n_1280),
.Y(n_1403)
);

O2A1O1Ixp5_ASAP7_75t_SL g1404 ( 
.A1(n_1239),
.A2(n_1240),
.B(n_1243),
.C(n_1254),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1258),
.A2(n_1261),
.B1(n_1262),
.B2(n_1203),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1236),
.A2(n_1279),
.B(n_1237),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1133),
.B(n_1247),
.Y(n_1407)
);

BUFx2_ASAP7_75t_R g1408 ( 
.A(n_1256),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1236),
.A2(n_1279),
.B(n_1237),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1147),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1133),
.B(n_1247),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_L g1412 ( 
.A(n_1246),
.B(n_1257),
.C(n_980),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1182),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1236),
.A2(n_1279),
.B(n_1237),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1264),
.B(n_868),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1246),
.B(n_1257),
.Y(n_1416)
);

O2A1O1Ixp5_ASAP7_75t_L g1417 ( 
.A1(n_1135),
.A2(n_1194),
.B(n_1257),
.C(n_1246),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1200),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1147),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1182),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1133),
.B(n_1247),
.Y(n_1421)
);

AO21x1_ASAP7_75t_L g1422 ( 
.A1(n_1246),
.A2(n_980),
.B(n_1257),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1264),
.B(n_868),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1222),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1184),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1186),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_SL g1427 ( 
.A1(n_1220),
.A2(n_882),
.B(n_1277),
.C(n_1235),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1147),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1184),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1133),
.B(n_1247),
.Y(n_1430)
);

INVx6_ASAP7_75t_L g1431 ( 
.A(n_1198),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1186),
.Y(n_1432)
);

NAND2x1p5_ASAP7_75t_L g1433 ( 
.A(n_1198),
.B(n_1218),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1246),
.A2(n_1257),
.B(n_1284),
.C(n_1128),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1186),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1264),
.B(n_868),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1182),
.B(n_947),
.Y(n_1437)
);

INVx5_ASAP7_75t_L g1438 ( 
.A(n_1198),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1182),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1127),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1236),
.A2(n_1279),
.B(n_1237),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1236),
.A2(n_1279),
.B(n_1237),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1186),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1226),
.A2(n_443),
.B1(n_448),
.B2(n_439),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1321),
.Y(n_1445)
);

NAND2x1p5_ASAP7_75t_L g1446 ( 
.A(n_1321),
.B(n_1337),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1309),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1314),
.Y(n_1448)
);

INVx6_ASAP7_75t_L g1449 ( 
.A(n_1290),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1320),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1415),
.B(n_1423),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1325),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1330),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1342),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1292),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1405),
.A2(n_1403),
.B(n_1383),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1290),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1392),
.A2(n_1366),
.B(n_1390),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1426),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1432),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1383),
.A2(n_1363),
.B(n_1333),
.Y(n_1461)
);

INVx4_ASAP7_75t_L g1462 ( 
.A(n_1321),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1435),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1304),
.A2(n_1310),
.B1(n_1345),
.B2(n_1416),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1345),
.A2(n_1304),
.B1(n_1379),
.B2(n_1326),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1310),
.A2(n_1422),
.B1(n_1412),
.B2(n_1444),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1443),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1431),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1436),
.B(n_1295),
.Y(n_1469)
);

AO21x2_ASAP7_75t_L g1470 ( 
.A1(n_1390),
.A2(n_1355),
.B(n_1398),
.Y(n_1470)
);

CKINVDCx6p67_ASAP7_75t_R g1471 ( 
.A(n_1296),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1340),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_1370),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1305),
.A2(n_1299),
.B1(n_1437),
.B2(n_1301),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1356),
.A2(n_1388),
.B1(n_1352),
.B2(n_1302),
.Y(n_1475)
);

INVx1_ASAP7_75t_SL g1476 ( 
.A(n_1318),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_SL g1477 ( 
.A1(n_1312),
.A2(n_1407),
.B1(n_1300),
.B2(n_1287),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1363),
.A2(n_1442),
.B(n_1441),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1404),
.A2(n_1384),
.B(n_1441),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1311),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1308),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1322),
.A2(n_1332),
.B1(n_1411),
.B2(n_1287),
.Y(n_1482)
);

AOI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1405),
.A2(n_1403),
.B(n_1324),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1425),
.Y(n_1484)
);

NAND2x1p5_ASAP7_75t_L g1485 ( 
.A(n_1321),
.B(n_1337),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1337),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1429),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1290),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1300),
.A2(n_1411),
.B1(n_1430),
.B2(n_1407),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1307),
.A2(n_1442),
.B(n_1409),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_SL g1491 ( 
.A(n_1319),
.Y(n_1491)
);

BUFx2_ASAP7_75t_SL g1492 ( 
.A(n_1289),
.Y(n_1492)
);

INVx6_ASAP7_75t_L g1493 ( 
.A(n_1424),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1434),
.A2(n_1430),
.B1(n_1421),
.B2(n_1335),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1355),
.A2(n_1398),
.B(n_1389),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1364),
.B(n_1303),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1298),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1346),
.Y(n_1498)
);

INVx1_ASAP7_75t_SL g1499 ( 
.A(n_1286),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1291),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1328),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1439),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1347),
.Y(n_1503)
);

AO21x1_ASAP7_75t_L g1504 ( 
.A1(n_1349),
.A2(n_1359),
.B(n_1362),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1338),
.A2(n_1344),
.B1(n_1391),
.B2(n_1396),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1413),
.A2(n_1420),
.B1(n_1322),
.B2(n_1386),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1328),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1438),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1349),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1323),
.Y(n_1510)
);

AOI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1322),
.A2(n_1317),
.B1(n_1364),
.B2(n_1316),
.Y(n_1511)
);

NAND2x1p5_ASAP7_75t_L g1512 ( 
.A(n_1438),
.B(n_1413),
.Y(n_1512)
);

AOI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1359),
.A2(n_1402),
.B(n_1387),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1420),
.B(n_1294),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1368),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1378),
.Y(n_1516)
);

AOI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1387),
.A2(n_1348),
.B(n_1381),
.Y(n_1517)
);

AOI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1348),
.A2(n_1381),
.B(n_1360),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1431),
.Y(n_1519)
);

AOI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1354),
.A2(n_1373),
.B(n_1385),
.Y(n_1520)
);

BUFx12f_ASAP7_75t_L g1521 ( 
.A(n_1285),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1368),
.Y(n_1522)
);

INVx1_ASAP7_75t_SL g1523 ( 
.A(n_1419),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1375),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1395),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1294),
.B(n_1410),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1362),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1357),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1424),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1357),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1311),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1406),
.A2(n_1414),
.B(n_1339),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1311),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1428),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1327),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1303),
.B(n_1306),
.Y(n_1536)
);

AOI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1382),
.A2(n_1358),
.B(n_1378),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1358),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1327),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1376),
.A2(n_1371),
.B1(n_1380),
.B2(n_1394),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1438),
.B(n_1306),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1377),
.B(n_1343),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1293),
.B(n_1353),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1288),
.B(n_1418),
.Y(n_1544)
);

AO21x1_ASAP7_75t_L g1545 ( 
.A1(n_1376),
.A2(n_1389),
.B(n_1397),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1313),
.B(n_1353),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1400),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1417),
.A2(n_1397),
.B1(n_1401),
.B2(n_1319),
.Y(n_1548)
);

AOI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1406),
.A2(n_1414),
.B(n_1350),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1336),
.A2(n_1431),
.B1(n_1365),
.B2(n_1341),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1334),
.A2(n_1433),
.B1(n_1374),
.B2(n_1372),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1327),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1331),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1369),
.B(n_1374),
.Y(n_1554)
);

BUFx8_ASAP7_75t_L g1555 ( 
.A(n_1331),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1361),
.B(n_1350),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1361),
.B(n_1367),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1334),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1329),
.A2(n_1440),
.B1(n_1351),
.B2(n_1367),
.Y(n_1559)
);

NAND2x1p5_ASAP7_75t_L g1560 ( 
.A(n_1361),
.B(n_1351),
.Y(n_1560)
);

NOR2x1_ASAP7_75t_SL g1561 ( 
.A(n_1399),
.B(n_1427),
.Y(n_1561)
);

CKINVDCx20_ASAP7_75t_R g1562 ( 
.A(n_1408),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1440),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1315),
.A2(n_1246),
.B1(n_1257),
.B2(n_955),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1315),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1315),
.A2(n_1345),
.B1(n_980),
.B2(n_1299),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1393),
.Y(n_1567)
);

NAND2x1p5_ASAP7_75t_L g1568 ( 
.A(n_1408),
.B(n_1321),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1309),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1309),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1309),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1309),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1345),
.A2(n_980),
.B1(n_1299),
.B2(n_1304),
.Y(n_1573)
);

BUFx2_ASAP7_75t_R g1574 ( 
.A(n_1285),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1309),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1309),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1304),
.A2(n_1257),
.B1(n_1246),
.B2(n_1283),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1309),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1290),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1328),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1290),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1309),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1309),
.Y(n_1583)
);

BUFx12f_ASAP7_75t_L g1584 ( 
.A(n_1285),
.Y(n_1584)
);

BUFx2_ASAP7_75t_SL g1585 ( 
.A(n_1289),
.Y(n_1585)
);

AO21x2_ASAP7_75t_L g1586 ( 
.A1(n_1392),
.A2(n_1228),
.B(n_1366),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1364),
.B(n_1303),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1340),
.Y(n_1588)
);

CKINVDCx11_ASAP7_75t_R g1589 ( 
.A(n_1296),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1309),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1309),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1415),
.B(n_1423),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_SL g1593 ( 
.A1(n_1345),
.A2(n_439),
.B1(n_448),
.B2(n_443),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1364),
.B(n_1303),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1345),
.A2(n_980),
.B1(n_1326),
.B2(n_1297),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1321),
.Y(n_1596)
);

OAI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1479),
.A2(n_1518),
.B(n_1456),
.Y(n_1597)
);

INVx5_ASAP7_75t_L g1598 ( 
.A(n_1508),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1516),
.B(n_1503),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1516),
.B(n_1495),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_R g1601 ( 
.A(n_1589),
.B(n_1521),
.Y(n_1601)
);

AO21x2_ASAP7_75t_L g1602 ( 
.A1(n_1566),
.A2(n_1573),
.B(n_1520),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1447),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1497),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1538),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1500),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1448),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1569),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1457),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1504),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1505),
.B(n_1509),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1567),
.B(n_1501),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1499),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1501),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1507),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1507),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1490),
.A2(n_1549),
.B(n_1517),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1580),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1545),
.A2(n_1483),
.B(n_1513),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1523),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1525),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1580),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1537),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1458),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1572),
.B(n_1575),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1547),
.B(n_1515),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1502),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1527),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1510),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1522),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1528),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1576),
.B(n_1578),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1458),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1589),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1582),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1530),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1586),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1586),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1512),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1470),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1474),
.B(n_1470),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1464),
.B(n_1547),
.Y(n_1643)
);

AOI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1540),
.A2(n_1461),
.B(n_1494),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1583),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1590),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1461),
.A2(n_1478),
.B(n_1532),
.Y(n_1647)
);

OAI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1461),
.A2(n_1478),
.B(n_1532),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1556),
.B(n_1542),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1591),
.Y(n_1650)
);

AO21x2_ASAP7_75t_L g1651 ( 
.A1(n_1566),
.A2(n_1573),
.B(n_1564),
.Y(n_1651)
);

BUFx4f_ASAP7_75t_SL g1652 ( 
.A(n_1521),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1514),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1478),
.A2(n_1532),
.B(n_1548),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1464),
.A2(n_1466),
.B1(n_1577),
.B2(n_1465),
.C(n_1482),
.Y(n_1655)
);

OA21x2_ASAP7_75t_L g1656 ( 
.A1(n_1577),
.A2(n_1548),
.B(n_1454),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1450),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1452),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1453),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1455),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1524),
.A2(n_1460),
.B(n_1467),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1565),
.Y(n_1662)
);

AO21x2_ASAP7_75t_L g1663 ( 
.A1(n_1561),
.A2(n_1459),
.B(n_1463),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1498),
.Y(n_1664)
);

AO21x1_ASAP7_75t_SL g1665 ( 
.A1(n_1466),
.A2(n_1511),
.B(n_1550),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1476),
.B(n_1469),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1481),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1449),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1526),
.Y(n_1669)
);

OAI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1477),
.A2(n_1489),
.B(n_1595),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1484),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1487),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1565),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1526),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1531),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1533),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1535),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1457),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1508),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1539),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1462),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1552),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1553),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1563),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1593),
.A2(n_1475),
.B1(n_1451),
.B2(n_1592),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1555),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1488),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1563),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1480),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1480),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1480),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1506),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1554),
.B(n_1542),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1506),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1542),
.B(n_1557),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1560),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1534),
.B(n_1529),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1568),
.B(n_1543),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1445),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1560),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1445),
.Y(n_1701)
);

CKINVDCx20_ASAP7_75t_R g1702 ( 
.A(n_1562),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1496),
.B(n_1587),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_SL g1704 ( 
.A(n_1472),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1486),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1486),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1596),
.Y(n_1707)
);

OR2x6_ASAP7_75t_L g1708 ( 
.A(n_1568),
.B(n_1446),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1596),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_1562),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1555),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1661),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1661),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1605),
.B(n_1588),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1679),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1632),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1605),
.B(n_1588),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1612),
.B(n_1588),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1612),
.B(n_1588),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1630),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1623),
.B(n_1472),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1661),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1623),
.B(n_1626),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1661),
.Y(n_1724)
);

AO21x2_ASAP7_75t_L g1725 ( 
.A1(n_1624),
.A2(n_1551),
.B(n_1559),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1645),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1633),
.B(n_1599),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1642),
.B(n_1473),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1633),
.B(n_1472),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1642),
.B(n_1473),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1609),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1645),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1646),
.Y(n_1733)
);

AND2x4_ASAP7_75t_SL g1734 ( 
.A(n_1708),
.B(n_1473),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1599),
.B(n_1546),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_R g1736 ( 
.A(n_1635),
.B(n_1471),
.Y(n_1736)
);

OAI211xp5_ASAP7_75t_L g1737 ( 
.A1(n_1670),
.A2(n_1550),
.B(n_1544),
.C(n_1579),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1646),
.B(n_1585),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1653),
.B(n_1492),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1669),
.B(n_1529),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1650),
.Y(n_1741)
);

NOR2xp67_ASAP7_75t_L g1742 ( 
.A(n_1674),
.B(n_1468),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1600),
.B(n_1579),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1604),
.Y(n_1744)
);

NAND3xp33_ASAP7_75t_L g1745 ( 
.A(n_1610),
.B(n_1555),
.C(n_1488),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1631),
.B(n_1581),
.Y(n_1746)
);

OAI31xp33_ASAP7_75t_L g1747 ( 
.A1(n_1655),
.A2(n_1551),
.A3(n_1587),
.B(n_1594),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1614),
.B(n_1471),
.Y(n_1748)
);

INVxp67_ASAP7_75t_L g1749 ( 
.A(n_1606),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1628),
.B(n_1449),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1651),
.A2(n_1491),
.B1(n_1587),
.B2(n_1496),
.C(n_1594),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1673),
.B(n_1594),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1675),
.Y(n_1753)
);

INVx4_ASAP7_75t_L g1754 ( 
.A(n_1681),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1614),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1663),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1615),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1629),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1651),
.A2(n_1491),
.B1(n_1519),
.B2(n_1468),
.C(n_1536),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1615),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1629),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1660),
.B(n_1493),
.Y(n_1762)
);

INVxp67_ASAP7_75t_SL g1763 ( 
.A(n_1610),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1662),
.B(n_1493),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1627),
.B(n_1508),
.Y(n_1765)
);

NOR3xp33_ASAP7_75t_SL g1766 ( 
.A(n_1684),
.B(n_1574),
.C(n_1584),
.Y(n_1766)
);

BUFx2_ASAP7_75t_L g1767 ( 
.A(n_1616),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1657),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1616),
.B(n_1519),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_SL g1770 ( 
.A1(n_1651),
.A2(n_1656),
.B1(n_1602),
.B2(n_1643),
.Y(n_1770)
);

OA21x2_ASAP7_75t_L g1771 ( 
.A1(n_1647),
.A2(n_1485),
.B(n_1558),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1658),
.Y(n_1772)
);

AO21x2_ASAP7_75t_L g1773 ( 
.A1(n_1624),
.A2(n_1541),
.B(n_1584),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1659),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1603),
.B(n_1607),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1663),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1608),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1636),
.B(n_1666),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1621),
.B(n_1693),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1621),
.B(n_1693),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1618),
.B(n_1622),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1667),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1666),
.B(n_1637),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1618),
.B(n_1622),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1716),
.B(n_1663),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1720),
.B(n_1744),
.Y(n_1786)
);

NAND3xp33_ASAP7_75t_L g1787 ( 
.A(n_1770),
.B(n_1688),
.C(n_1684),
.Y(n_1787)
);

AOI211xp5_ASAP7_75t_L g1788 ( 
.A1(n_1737),
.A2(n_1654),
.B(n_1698),
.C(n_1643),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1753),
.B(n_1637),
.Y(n_1789)
);

OAI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1728),
.A2(n_1656),
.B1(n_1611),
.B2(n_1708),
.Y(n_1790)
);

NAND3xp33_ASAP7_75t_L g1791 ( 
.A(n_1756),
.B(n_1688),
.C(n_1682),
.Y(n_1791)
);

OAI21xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1759),
.A2(n_1644),
.B(n_1711),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1749),
.B(n_1676),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1784),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1776),
.B(n_1676),
.C(n_1682),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1718),
.A2(n_1685),
.B1(n_1710),
.B2(n_1702),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1727),
.B(n_1677),
.Y(n_1797)
);

AOI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1763),
.A2(n_1677),
.B1(n_1680),
.B2(n_1692),
.C(n_1694),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_L g1799 ( 
.A(n_1748),
.B(n_1691),
.C(n_1689),
.D(n_1697),
.Y(n_1799)
);

OA211x2_ASAP7_75t_L g1800 ( 
.A1(n_1751),
.A2(n_1704),
.B(n_1601),
.C(n_1665),
.Y(n_1800)
);

OA21x2_ASAP7_75t_L g1801 ( 
.A1(n_1712),
.A2(n_1648),
.B(n_1647),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1727),
.B(n_1723),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1723),
.B(n_1779),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1783),
.B(n_1680),
.Y(n_1804)
);

OAI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1747),
.A2(n_1698),
.B1(n_1656),
.B2(n_1611),
.C(n_1620),
.Y(n_1805)
);

OAI21xp33_ASAP7_75t_L g1806 ( 
.A1(n_1781),
.A2(n_1641),
.B(n_1654),
.Y(n_1806)
);

NAND3xp33_ASAP7_75t_SL g1807 ( 
.A(n_1736),
.B(n_1613),
.C(n_1711),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1725),
.A2(n_1634),
.B(n_1625),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1779),
.B(n_1625),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1728),
.A2(n_1692),
.B1(n_1665),
.B2(n_1656),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1735),
.B(n_1695),
.Y(n_1811)
);

NAND4xp25_ASAP7_75t_L g1812 ( 
.A(n_1748),
.B(n_1689),
.C(n_1691),
.D(n_1686),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1735),
.B(n_1683),
.Y(n_1813)
);

NAND3xp33_ASAP7_75t_L g1814 ( 
.A(n_1730),
.B(n_1634),
.C(n_1709),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1778),
.B(n_1683),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1738),
.B(n_1678),
.Y(n_1816)
);

OAI211xp5_ASAP7_75t_L g1817 ( 
.A1(n_1750),
.A2(n_1686),
.B(n_1701),
.C(n_1709),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1742),
.B(n_1678),
.Y(n_1818)
);

OAI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1766),
.A2(n_1664),
.B1(n_1671),
.B2(n_1672),
.C(n_1696),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1780),
.B(n_1619),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1780),
.B(n_1719),
.Y(n_1821)
);

OA21x2_ASAP7_75t_L g1822 ( 
.A1(n_1713),
.A2(n_1648),
.B(n_1597),
.Y(n_1822)
);

NOR3xp33_ASAP7_75t_SL g1823 ( 
.A(n_1745),
.B(n_1652),
.C(n_1701),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1738),
.B(n_1687),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1740),
.B(n_1687),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1719),
.B(n_1619),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1768),
.B(n_1772),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1714),
.B(n_1619),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1784),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1714),
.B(n_1619),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_SL g1831 ( 
.A1(n_1725),
.A2(n_1704),
.B1(n_1627),
.B2(n_1640),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1717),
.B(n_1641),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1768),
.B(n_1705),
.Y(n_1833)
);

OA21x2_ASAP7_75t_L g1834 ( 
.A1(n_1722),
.A2(n_1724),
.B(n_1617),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1772),
.B(n_1705),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1717),
.B(n_1641),
.Y(n_1836)
);

OAI21xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1734),
.A2(n_1681),
.B(n_1703),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1739),
.B(n_1668),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1721),
.B(n_1638),
.Y(n_1839)
);

NAND3xp33_ASAP7_75t_L g1840 ( 
.A(n_1769),
.B(n_1707),
.C(n_1699),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1774),
.B(n_1707),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1769),
.B(n_1706),
.C(n_1699),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1774),
.B(n_1690),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1777),
.B(n_1690),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1777),
.B(n_1706),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1746),
.B(n_1700),
.Y(n_1846)
);

NOR3xp33_ASAP7_75t_L g1847 ( 
.A(n_1762),
.B(n_1696),
.C(n_1639),
.Y(n_1847)
);

NAND3xp33_ASAP7_75t_L g1848 ( 
.A(n_1755),
.B(n_1760),
.C(n_1757),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1758),
.B(n_1664),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1758),
.B(n_1649),
.Y(n_1850)
);

AND2x2_ASAP7_75t_SL g1851 ( 
.A(n_1734),
.B(n_1703),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1729),
.B(n_1639),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1715),
.B(n_1679),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1820),
.B(n_1803),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1802),
.B(n_1755),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1794),
.B(n_1757),
.Y(n_1856)
);

BUFx3_ASAP7_75t_L g1857 ( 
.A(n_1851),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1794),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1829),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1829),
.B(n_1760),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1826),
.B(n_1752),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1834),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1785),
.B(n_1767),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1834),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1834),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1827),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1801),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1849),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1828),
.B(n_1754),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1801),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1830),
.B(n_1767),
.Y(n_1871)
);

NOR2x1_ASAP7_75t_L g1872 ( 
.A(n_1848),
.B(n_1731),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1801),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1791),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1833),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1807),
.B(n_1739),
.Y(n_1876)
);

NAND2x1p5_ASAP7_75t_SL g1877 ( 
.A(n_1818),
.B(n_1668),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1835),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1786),
.Y(n_1879)
);

AND2x2_ASAP7_75t_SL g1880 ( 
.A(n_1851),
.B(n_1765),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1841),
.B(n_1761),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1809),
.B(n_1741),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_L g1883 ( 
.A(n_1792),
.B(n_1731),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1845),
.B(n_1761),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1821),
.B(n_1839),
.Y(n_1885)
);

NAND2x1_ASAP7_75t_L g1886 ( 
.A(n_1840),
.B(n_1754),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1804),
.B(n_1741),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1797),
.B(n_1775),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1843),
.Y(n_1889)
);

NAND2x1p5_ASAP7_75t_L g1890 ( 
.A(n_1818),
.B(n_1771),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1844),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1813),
.B(n_1743),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1789),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1793),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1822),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1795),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1815),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1825),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1847),
.B(n_1782),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1842),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1822),
.Y(n_1901)
);

INVx4_ASAP7_75t_R g1902 ( 
.A(n_1852),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1896),
.B(n_1850),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1881),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1881),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1896),
.B(n_1874),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1884),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1874),
.B(n_1798),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1900),
.B(n_1811),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1884),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1857),
.B(n_1814),
.Y(n_1911)
);

OR2x6_ASAP7_75t_L g1912 ( 
.A(n_1883),
.B(n_1808),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1866),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1894),
.B(n_1817),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1866),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1900),
.B(n_1846),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1899),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1855),
.B(n_1879),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1857),
.B(n_1773),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1899),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1868),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1875),
.B(n_1726),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1868),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1862),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1854),
.B(n_1852),
.Y(n_1925)
);

OR2x6_ASAP7_75t_L g1926 ( 
.A(n_1883),
.B(n_1890),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1875),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1878),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1876),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1854),
.B(n_1832),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1862),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1878),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1863),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1855),
.B(n_1799),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1887),
.Y(n_1935)
);

OR2x2_ASAP7_75t_L g1936 ( 
.A(n_1879),
.B(n_1816),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1854),
.B(n_1832),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1889),
.B(n_1732),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1889),
.B(n_1733),
.Y(n_1939)
);

NAND4xp25_ASAP7_75t_SL g1940 ( 
.A(n_1872),
.B(n_1788),
.C(n_1810),
.D(n_1805),
.Y(n_1940)
);

NAND4xp75_ASAP7_75t_L g1941 ( 
.A(n_1872),
.B(n_1800),
.C(n_1823),
.D(n_1853),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1863),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1892),
.B(n_1824),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1887),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1891),
.B(n_1782),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1892),
.B(n_1812),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1857),
.B(n_1836),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1888),
.B(n_1836),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1885),
.B(n_1838),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1862),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1885),
.B(n_1837),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1898),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1869),
.B(n_1773),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1885),
.B(n_1764),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1858),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1924),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1922),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1909),
.B(n_1888),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1909),
.B(n_1871),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1924),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1931),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1931),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1917),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1917),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1920),
.B(n_1893),
.Y(n_1965)
);

OAI21xp33_ASAP7_75t_L g1966 ( 
.A1(n_1906),
.A2(n_1871),
.B(n_1860),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1920),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1938),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1939),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1916),
.B(n_1856),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1908),
.B(n_1891),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1951),
.B(n_1861),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1951),
.B(n_1861),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1955),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1952),
.B(n_1880),
.Y(n_1975)
);

O2A1O1Ixp33_ASAP7_75t_SL g1976 ( 
.A1(n_1929),
.A2(n_1886),
.B(n_1877),
.C(n_1860),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1941),
.A2(n_1880),
.B1(n_1787),
.B2(n_1886),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1921),
.Y(n_1978)
);

NOR2xp67_ASAP7_75t_SL g1979 ( 
.A(n_1918),
.B(n_1598),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1903),
.B(n_1882),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1923),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1925),
.B(n_1930),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1935),
.B(n_1856),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1926),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1944),
.B(n_1858),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1925),
.B(n_1861),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1950),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1950),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1930),
.B(n_1937),
.Y(n_1989)
);

INVx2_ASAP7_75t_SL g1990 ( 
.A(n_1926),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1940),
.A2(n_1880),
.B(n_1806),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1948),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1927),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1928),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1932),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1914),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1913),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1912),
.A2(n_1800),
.B1(n_1796),
.B2(n_1790),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1904),
.B(n_1882),
.Y(n_1999)
);

AOI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1912),
.A2(n_1890),
.B(n_1859),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1915),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1933),
.B(n_1859),
.Y(n_2002)
);

INVx1_ASAP7_75t_SL g2003 ( 
.A(n_1936),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1905),
.B(n_1882),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1945),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1912),
.A2(n_1831),
.B1(n_1819),
.B2(n_1897),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1972),
.B(n_1933),
.Y(n_2007)
);

NAND2xp33_ASAP7_75t_SL g2008 ( 
.A(n_1977),
.B(n_1946),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1997),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1956),
.Y(n_2010)
);

BUFx2_ASAP7_75t_L g2011 ( 
.A(n_1974),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_2002),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1958),
.B(n_1907),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_2003),
.B(n_1910),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1970),
.B(n_1942),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1970),
.B(n_1942),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_2002),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1956),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1972),
.B(n_1949),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1960),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1978),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1996),
.B(n_1934),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1981),
.Y(n_2023)
);

INVx1_ASAP7_75t_SL g2024 ( 
.A(n_1965),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1960),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1957),
.B(n_1949),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1973),
.B(n_1947),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1993),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1994),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1995),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2001),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1963),
.B(n_1964),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1961),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1967),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1982),
.B(n_1926),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1973),
.B(n_1947),
.Y(n_2036)
);

BUFx12f_ASAP7_75t_L g2037 ( 
.A(n_1984),
.Y(n_2037)
);

BUFx2_ASAP7_75t_L g2038 ( 
.A(n_1975),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1985),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1985),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1983),
.B(n_1943),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1982),
.B(n_1937),
.Y(n_2042)
);

INVx1_ASAP7_75t_SL g2043 ( 
.A(n_1971),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1989),
.B(n_1911),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1968),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1969),
.Y(n_2046)
);

AOI221xp5_ASAP7_75t_L g2047 ( 
.A1(n_2008),
.A2(n_1991),
.B1(n_1976),
.B2(n_2000),
.C(n_1966),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2011),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_2043),
.B(n_1975),
.Y(n_2049)
);

AOI32xp33_ASAP7_75t_L g2050 ( 
.A1(n_2038),
.A2(n_1911),
.A3(n_1990),
.B1(n_1984),
.B2(n_1919),
.Y(n_2050)
);

OAI21xp33_ASAP7_75t_L g2051 ( 
.A1(n_2022),
.A2(n_2005),
.B(n_1992),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_2041),
.B(n_1992),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_2035),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_2041),
.B(n_2015),
.Y(n_2054)
);

O2A1O1Ixp33_ASAP7_75t_L g2055 ( 
.A1(n_2043),
.A2(n_1976),
.B(n_1912),
.C(n_1926),
.Y(n_2055)
);

OAI32xp33_ASAP7_75t_L g2056 ( 
.A1(n_2015),
.A2(n_1990),
.A3(n_1959),
.B1(n_1980),
.B2(n_1983),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2019),
.B(n_2044),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2011),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2038),
.B(n_1989),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2024),
.B(n_1986),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_2044),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2019),
.B(n_1986),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2028),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2027),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2032),
.Y(n_2065)
);

AOI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2037),
.A2(n_1998),
.B1(n_2006),
.B2(n_1911),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_2027),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_2035),
.A2(n_2004),
.B1(n_1999),
.B2(n_1953),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2032),
.Y(n_2069)
);

AOI221x1_ASAP7_75t_SL g2070 ( 
.A1(n_2012),
.A2(n_1953),
.B1(n_1867),
.B2(n_1873),
.C(n_1870),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2007),
.B(n_2009),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_2035),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2021),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2007),
.B(n_1954),
.Y(n_2074)
);

NOR2xp33_ASAP7_75t_L g2075 ( 
.A(n_2037),
.B(n_1979),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2054),
.Y(n_2076)
);

NOR2xp33_ASAP7_75t_L g2077 ( 
.A(n_2053),
.B(n_2037),
.Y(n_2077)
);

INVxp67_ASAP7_75t_SL g2078 ( 
.A(n_2049),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_2057),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2052),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2064),
.Y(n_2081)
);

NOR2x1_ASAP7_75t_L g2082 ( 
.A(n_2048),
.B(n_2034),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_2061),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2057),
.B(n_2042),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2064),
.B(n_2042),
.Y(n_2085)
);

INVx3_ASAP7_75t_L g2086 ( 
.A(n_2053),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2062),
.B(n_2036),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2061),
.Y(n_2088)
);

INVx1_ASAP7_75t_SL g2089 ( 
.A(n_2059),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2067),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_2053),
.B(n_2016),
.Y(n_2091)
);

AOI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_2047),
.A2(n_2033),
.B1(n_2018),
.B2(n_2025),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2067),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2049),
.B(n_2036),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_2055),
.B(n_2035),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2073),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2058),
.B(n_2012),
.Y(n_2097)
);

AOI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_2056),
.A2(n_2016),
.B(n_2014),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_2078),
.B(n_2072),
.Y(n_2099)
);

AOI211xp5_ASAP7_75t_L g2100 ( 
.A1(n_2098),
.A2(n_2075),
.B(n_2066),
.C(n_2051),
.Y(n_2100)
);

OR3x1_ASAP7_75t_L g2101 ( 
.A(n_2077),
.B(n_2075),
.C(n_2069),
.Y(n_2101)
);

AOI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_2092),
.A2(n_2072),
.B1(n_2060),
.B2(n_2065),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2083),
.Y(n_2103)
);

AOI211xp5_ASAP7_75t_L g2104 ( 
.A1(n_2095),
.A2(n_2091),
.B(n_2076),
.C(n_2089),
.Y(n_2104)
);

O2A1O1Ixp33_ASAP7_75t_SL g2105 ( 
.A1(n_2094),
.A2(n_2071),
.B(n_2063),
.C(n_2072),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2087),
.B(n_2070),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2087),
.B(n_2074),
.Y(n_2107)
);

AOI222xp33_ASAP7_75t_L g2108 ( 
.A1(n_2080),
.A2(n_2076),
.B1(n_2082),
.B2(n_2088),
.C1(n_2096),
.C2(n_2093),
.Y(n_2108)
);

OAI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_2079),
.A2(n_2046),
.B(n_2045),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2079),
.B(n_2026),
.Y(n_2110)
);

AOI221xp5_ASAP7_75t_SL g2111 ( 
.A1(n_2097),
.A2(n_2034),
.B1(n_2046),
.B2(n_2045),
.C(n_2017),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2084),
.B(n_2017),
.Y(n_2112)
);

NOR3xp33_ASAP7_75t_L g2113 ( 
.A(n_2099),
.B(n_2086),
.C(n_2080),
.Y(n_2113)
);

OA22x2_ASAP7_75t_L g2114 ( 
.A1(n_2102),
.A2(n_2088),
.B1(n_2093),
.B2(n_2090),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2107),
.B(n_2086),
.Y(n_2115)
);

NOR2xp67_ASAP7_75t_L g2116 ( 
.A(n_2103),
.B(n_2086),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2110),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2108),
.B(n_2085),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2104),
.B(n_2081),
.Y(n_2119)
);

OA211x2_ASAP7_75t_L g2120 ( 
.A1(n_2106),
.A2(n_2050),
.B(n_2090),
.C(n_2081),
.Y(n_2120)
);

NAND3xp33_ASAP7_75t_L g2121 ( 
.A(n_2100),
.B(n_2105),
.C(n_2111),
.Y(n_2121)
);

AND4x1_ASAP7_75t_L g2122 ( 
.A(n_2109),
.B(n_2096),
.C(n_2039),
.D(n_2040),
.Y(n_2122)
);

OAI211xp5_ASAP7_75t_L g2123 ( 
.A1(n_2111),
.A2(n_2039),
.B(n_2040),
.C(n_2068),
.Y(n_2123)
);

NAND3xp33_ASAP7_75t_L g2124 ( 
.A(n_2121),
.B(n_2112),
.C(n_2023),
.Y(n_2124)
);

NOR2x1_ASAP7_75t_L g2125 ( 
.A(n_2116),
.B(n_2101),
.Y(n_2125)
);

NAND2x1p5_ASAP7_75t_L g2126 ( 
.A(n_2117),
.B(n_2021),
.Y(n_2126)
);

NOR3xp33_ASAP7_75t_SL g2127 ( 
.A(n_2119),
.B(n_2029),
.C(n_2023),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_2115),
.B(n_2029),
.Y(n_2128)
);

INVxp33_ASAP7_75t_L g2129 ( 
.A(n_2113),
.Y(n_2129)
);

NOR2x1_ASAP7_75t_L g2130 ( 
.A(n_2118),
.B(n_2030),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2126),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2130),
.B(n_2122),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2128),
.Y(n_2133)
);

AOI22xp5_ASAP7_75t_L g2134 ( 
.A1(n_2125),
.A2(n_2120),
.B1(n_2114),
.B2(n_2123),
.Y(n_2134)
);

INVxp67_ASAP7_75t_L g2135 ( 
.A(n_2124),
.Y(n_2135)
);

AOI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_2129),
.A2(n_2033),
.B1(n_2010),
.B2(n_2018),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2127),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2126),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2133),
.B(n_2030),
.Y(n_2139)
);

OAI311xp33_ASAP7_75t_L g2140 ( 
.A1(n_2134),
.A2(n_2013),
.A3(n_2031),
.B1(n_2025),
.C1(n_2020),
.Y(n_2140)
);

NAND4xp25_ASAP7_75t_L g2141 ( 
.A(n_2132),
.B(n_2031),
.C(n_2013),
.D(n_2025),
.Y(n_2141)
);

NOR4xp25_ASAP7_75t_L g2142 ( 
.A(n_2135),
.B(n_2033),
.C(n_2020),
.D(n_2018),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2137),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2131),
.Y(n_2144)
);

AOI221xp5_ASAP7_75t_L g2145 ( 
.A1(n_2136),
.A2(n_2020),
.B1(n_2010),
.B2(n_1864),
.C(n_1865),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_2139),
.Y(n_2146)
);

NAND4xp75_ASAP7_75t_L g2147 ( 
.A(n_2144),
.B(n_2138),
.C(n_2010),
.D(n_1962),
.Y(n_2147)
);

INVxp33_ASAP7_75t_SL g2148 ( 
.A(n_2143),
.Y(n_2148)
);

NAND2xp33_ASAP7_75t_L g2149 ( 
.A(n_2140),
.B(n_1961),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2142),
.B(n_1954),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2150),
.Y(n_2151)
);

INVxp67_ASAP7_75t_L g2152 ( 
.A(n_2147),
.Y(n_2152)
);

OR4x2_ASAP7_75t_L g2153 ( 
.A(n_2151),
.B(n_2148),
.C(n_2141),
.D(n_2146),
.Y(n_2153)
);

NAND3xp33_ASAP7_75t_L g2154 ( 
.A(n_2152),
.B(n_2149),
.C(n_2145),
.Y(n_2154)
);

OAI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_2154),
.A2(n_2153),
.B(n_1987),
.Y(n_2155)
);

AOI21xp33_ASAP7_75t_L g2156 ( 
.A1(n_2154),
.A2(n_1987),
.B(n_1962),
.Y(n_2156)
);

AOI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_2155),
.A2(n_1988),
.B(n_1870),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2156),
.Y(n_2158)
);

AO21x1_ASAP7_75t_L g2159 ( 
.A1(n_2158),
.A2(n_2157),
.B(n_1988),
.Y(n_2159)
);

AO21x2_ASAP7_75t_L g2160 ( 
.A1(n_2158),
.A2(n_1877),
.B(n_1870),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_2159),
.B(n_1864),
.Y(n_2161)
);

AOI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_2161),
.A2(n_2160),
.B1(n_1895),
.B2(n_1901),
.Y(n_2162)
);

OAI221xp5_ASAP7_75t_R g2163 ( 
.A1(n_2162),
.A2(n_1877),
.B1(n_1902),
.B2(n_1953),
.C(n_1919),
.Y(n_2163)
);

AOI211xp5_ASAP7_75t_L g2164 ( 
.A1(n_2163),
.A2(n_1919),
.B(n_1865),
.C(n_1864),
.Y(n_2164)
);


endmodule