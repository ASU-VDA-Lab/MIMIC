module fake_jpeg_648_n_78 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_32),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_27),
.B1(n_25),
.B2(n_23),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_37),
.B1(n_32),
.B2(n_25),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_24),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_33),
.B(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_44),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_45),
.B(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_24),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_26),
.C(n_22),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_53),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_59),
.B1(n_54),
.B2(n_57),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_40),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.C(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_35),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_32),
.B1(n_31),
.B2(n_35),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_20),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_52),
.C(n_19),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_49),
.B(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_1),
.Y(n_63)
);

A2O1A1O1Ixp25_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_65),
.B(n_66),
.C(n_5),
.D(n_6),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_67),
.B1(n_2),
.B2(n_3),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_2),
.B(n_3),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

MAJx2_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_18),
.C(n_16),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_71),
.C(n_15),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.A3(n_70),
.B1(n_68),
.B2(n_13),
.C1(n_14),
.C2(n_10),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_7),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_9),
.C(n_10),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_9),
.Y(n_78)
);


endmodule