module fake_jpeg_14681_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_182;
wire n_19;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_266;
wire n_218;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_SL g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_45),
.B(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_7),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_17),
.B(n_6),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_27),
.Y(n_83)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx5_ASAP7_75t_SL g103 ( 
.A(n_53),
.Y(n_103)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_37),
.B1(n_15),
.B2(n_16),
.Y(n_79)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_17),
.B(n_8),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_59),
.B(n_63),
.Y(n_102)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_28),
.B(n_5),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_15),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_26),
.B1(n_35),
.B2(n_38),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_67),
.B1(n_91),
.B2(n_33),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_37),
.B1(n_15),
.B2(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_69),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_32),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_41),
.B1(n_42),
.B2(n_56),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_21),
.C(n_23),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_90),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_39),
.A2(n_29),
.B(n_36),
.C(n_27),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_82),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_100),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_29),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_92),
.B(n_9),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_86),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_23),
.C(n_25),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_37),
.B1(n_36),
.B2(n_20),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_36),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_40),
.A2(n_27),
.B1(n_16),
.B2(n_30),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_18),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_35),
.B1(n_26),
.B2(n_16),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_21),
.B(n_23),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_43),
.B(n_30),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_18),
.Y(n_101)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_51),
.B(n_33),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_105),
.B(n_4),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_18),
.Y(n_107)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_109),
.A2(n_111),
.B1(n_119),
.B2(n_129),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_122),
.Y(n_157)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_25),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_113),
.B(n_116),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_25),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_117),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_10),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_76),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_135),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_67),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_46),
.B(n_62),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_128),
.A2(n_106),
.B(n_111),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_75),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_129)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_66),
.B1(n_74),
.B2(n_79),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_1),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_9),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_75),
.A2(n_13),
.B1(n_14),
.B2(n_3),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_140),
.B1(n_142),
.B2(n_145),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_93),
.B1(n_108),
.B2(n_74),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_144),
.Y(n_171)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_83),
.A2(n_1),
.B1(n_4),
.B2(n_80),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g146 ( 
.A(n_94),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_77),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_4),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_94),
.Y(n_164)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_152),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_90),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_156),
.B(n_174),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_168),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_175),
.B1(n_182),
.B2(n_184),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_161),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_179),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_72),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_125),
.A2(n_77),
.B1(n_73),
.B2(n_81),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_114),
.B(n_73),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_134),
.B(n_145),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_126),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_130),
.A2(n_86),
.B1(n_96),
.B2(n_81),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_125),
.B(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_188),
.B(n_197),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_183),
.A2(n_109),
.B1(n_125),
.B2(n_137),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_189),
.A2(n_194),
.B1(n_207),
.B2(n_208),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_140),
.B(n_129),
.C(n_128),
.Y(n_190)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_208),
.B(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_195),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_136),
.B1(n_144),
.B2(n_118),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_154),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_138),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_179),
.B(n_153),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_162),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_165),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_212),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_139),
.B1(n_141),
.B2(n_132),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_160),
.A2(n_146),
.B1(n_115),
.B2(n_120),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_153),
.A2(n_115),
.B(n_124),
.C(n_146),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_184),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_213),
.B(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_156),
.C(n_181),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_221),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_199),
.Y(n_217)
);

AOI221xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_207),
.B1(n_196),
.B2(n_202),
.C(n_197),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_223),
.B1(n_194),
.B2(n_193),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_166),
.C(n_177),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_166),
.C(n_177),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_196),
.B1(n_188),
.B2(n_205),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_179),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_198),
.B(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_161),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_161),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_169),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

OAI322xp33_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_225),
.A3(n_227),
.B1(n_216),
.B2(n_220),
.C1(n_221),
.C2(n_228),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_167),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

A2O1A1O1Ixp25_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_190),
.B(n_187),
.C(n_189),
.D(n_201),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_223),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_243),
.B1(n_248),
.B2(n_214),
.Y(n_260)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_241),
.C(n_250),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_203),
.B(n_155),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_234),
.B(n_224),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_155),
.B1(n_167),
.B2(n_209),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_223),
.A2(n_168),
.B1(n_180),
.B2(n_158),
.Y(n_248)
);

OAI322xp33_ASAP7_75t_L g251 ( 
.A1(n_231),
.A2(n_203),
.A3(n_204),
.B1(n_159),
.B2(n_178),
.C1(n_110),
.C2(n_158),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_235),
.C(n_222),
.Y(n_264)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_234),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_252),
.Y(n_259)
);

NOR3xp33_ASAP7_75t_SL g253 ( 
.A(n_228),
.B(n_204),
.C(n_203),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_233),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_257),
.C(n_264),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_263),
.B1(n_265),
.B2(n_242),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_262),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_217),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_247),
.A2(n_224),
.B(n_215),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_214),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_215),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_246),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_269),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_236),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_254),
.A2(n_245),
.B1(n_236),
.B2(n_253),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_272),
.B(n_274),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_241),
.C(n_240),
.Y(n_274)
);

OAI31xp33_ASAP7_75t_L g275 ( 
.A1(n_266),
.A2(n_245),
.A3(n_237),
.B(n_248),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_275),
.A2(n_263),
.B(n_265),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_259),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_260),
.B1(n_259),
.B2(n_264),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_283),
.B1(n_272),
.B2(n_268),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_280),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_235),
.Y(n_280)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_282),
.A2(n_274),
.B(n_232),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_281),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_279),
.A2(n_270),
.B(n_273),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_287),
.C(n_267),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_277),
.B(n_281),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_232),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_289),
.A2(n_285),
.B(n_226),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_291),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_218),
.B1(n_226),
.B2(n_292),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_218),
.Y(n_295)
);


endmodule