module real_aes_2668_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_762;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_0), .B(n_482), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_1), .A2(n_481), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_2), .B(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_3), .B(n_271), .Y(n_507) );
INVx1_ASAP7_75t_L g145 ( .A(n_4), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_5), .B(n_164), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_6), .B(n_271), .Y(n_536) );
INVx1_ASAP7_75t_L g173 ( .A(n_7), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g780 ( .A(n_8), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_9), .Y(n_190) );
NAND2xp33_ASAP7_75t_L g577 ( .A(n_10), .B(n_268), .Y(n_577) );
INVx2_ASAP7_75t_L g134 ( .A(n_11), .Y(n_134) );
AOI221x1_ASAP7_75t_L g480 ( .A1(n_12), .A2(n_25), .B1(n_481), .B2(n_482), .C(n_483), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_13), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_14), .B(n_482), .Y(n_573) );
INVx1_ASAP7_75t_L g269 ( .A(n_15), .Y(n_269) );
AO21x2_ASAP7_75t_L g571 ( .A1(n_16), .A2(n_170), .B(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_17), .B(n_216), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_18), .B(n_271), .Y(n_560) );
AO21x1_ASAP7_75t_L g502 ( .A1(n_19), .A2(n_482), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g113 ( .A(n_20), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_21), .Y(n_115) );
INVx1_ASAP7_75t_L g266 ( .A(n_22), .Y(n_266) );
INVx1_ASAP7_75t_SL g231 ( .A(n_23), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_24), .B(n_151), .Y(n_252) );
AOI33xp33_ASAP7_75t_L g202 ( .A1(n_26), .A2(n_53), .A3(n_140), .B1(n_149), .B2(n_203), .B3(n_204), .Y(n_202) );
NAND2x1_ASAP7_75t_L g494 ( .A(n_27), .B(n_271), .Y(n_494) );
NAND2x1_ASAP7_75t_L g535 ( .A(n_28), .B(n_268), .Y(n_535) );
INVx1_ASAP7_75t_L g182 ( .A(n_29), .Y(n_182) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_30), .A2(n_85), .B(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g165 ( .A(n_30), .B(n_85), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_31), .B(n_159), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_32), .B(n_268), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_33), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_34), .B(n_271), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_35), .B(n_268), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_36), .A2(n_481), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g139 ( .A(n_37), .Y(n_139) );
AND2x2_ASAP7_75t_L g157 ( .A(n_37), .B(n_145), .Y(n_157) );
AND2x2_ASAP7_75t_L g163 ( .A(n_37), .B(n_142), .Y(n_163) );
OR2x6_ASAP7_75t_L g111 ( .A(n_38), .B(n_112), .Y(n_111) );
NOR3xp33_ASAP7_75t_L g778 ( .A(n_38), .B(n_779), .C(n_781), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_39), .Y(n_185) );
OAI22xp33_ASAP7_75t_L g769 ( .A1(n_40), .A2(n_473), .B1(n_759), .B2(n_770), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_40), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_41), .B(n_482), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_42), .B(n_159), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_43), .A2(n_132), .B1(n_164), .B2(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_44), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_45), .B(n_151), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_46), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_47), .B(n_268), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_48), .B(n_170), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_49), .B(n_151), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_50), .A2(n_481), .B(n_534), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_51), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_52), .B(n_268), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_54), .B(n_151), .Y(n_214) );
INVx1_ASAP7_75t_L g144 ( .A(n_55), .Y(n_144) );
INVx1_ASAP7_75t_L g153 ( .A(n_55), .Y(n_153) );
AND2x2_ASAP7_75t_L g215 ( .A(n_56), .B(n_216), .Y(n_215) );
AOI221xp5_ASAP7_75t_L g171 ( .A1(n_57), .A2(n_74), .B1(n_137), .B2(n_159), .C(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_58), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_59), .B(n_271), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_60), .B(n_132), .Y(n_192) );
AOI21xp5_ASAP7_75t_SL g136 ( .A1(n_61), .A2(n_137), .B(n_146), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_62), .A2(n_481), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g263 ( .A(n_63), .Y(n_263) );
AO21x1_ASAP7_75t_L g504 ( .A1(n_64), .A2(n_481), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_65), .B(n_482), .Y(n_525) );
INVx1_ASAP7_75t_L g213 ( .A(n_66), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_67), .B(n_482), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_68), .A2(n_137), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g518 ( .A(n_69), .B(n_217), .Y(n_518) );
INVx1_ASAP7_75t_L g142 ( .A(n_70), .Y(n_142) );
INVx1_ASAP7_75t_L g155 ( .A(n_70), .Y(n_155) );
AND2x2_ASAP7_75t_L g538 ( .A(n_71), .B(n_131), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_72), .B(n_159), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_73), .Y(n_783) );
AND2x2_ASAP7_75t_L g233 ( .A(n_75), .B(n_131), .Y(n_233) );
INVx1_ASAP7_75t_L g264 ( .A(n_76), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_77), .A2(n_137), .B(n_230), .Y(n_229) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_78), .A2(n_137), .B(n_197), .C(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g114 ( .A(n_79), .Y(n_114) );
AND2x2_ASAP7_75t_L g523 ( .A(n_80), .B(n_131), .Y(n_523) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_81), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_82), .B(n_482), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_83), .A2(n_137), .B1(n_200), .B2(n_201), .Y(n_199) );
AND2x2_ASAP7_75t_L g503 ( .A(n_84), .B(n_164), .Y(n_503) );
AND2x2_ASAP7_75t_L g497 ( .A(n_86), .B(n_131), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_87), .B(n_268), .Y(n_561) );
INVx1_ASAP7_75t_L g147 ( .A(n_88), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_89), .A2(n_755), .B1(n_757), .B2(n_762), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_90), .B(n_271), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_91), .B(n_268), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_92), .A2(n_481), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g206 ( .A(n_93), .B(n_131), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_94), .B(n_271), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_95), .A2(n_180), .B(n_181), .C(n_184), .Y(n_179) );
BUFx2_ASAP7_75t_L g118 ( .A(n_96), .Y(n_118) );
BUFx2_ASAP7_75t_SL g767 ( .A(n_96), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_97), .A2(n_481), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_98), .B(n_151), .Y(n_150) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_774), .B(n_782), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_119), .B(n_764), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g101 ( .A(n_102), .B(n_116), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_103), .A2(n_769), .B(n_771), .Y(n_768) );
NOR2xp33_ASAP7_75t_SL g103 ( .A(n_104), .B(n_115), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_R g773 ( .A(n_108), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
OR2x6_ASAP7_75t_SL g468 ( .A(n_109), .B(n_110), .Y(n_468) );
AND2x6_ASAP7_75t_SL g472 ( .A(n_109), .B(n_111), .Y(n_472) );
OR2x2_ASAP7_75t_L g763 ( .A(n_109), .B(n_111), .Y(n_763) );
CKINVDCx16_ASAP7_75t_R g781 ( .A(n_109), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_113), .B(n_114), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_755), .B(n_756), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_466), .B1(n_469), .B2(n_473), .Y(n_121) );
INVx2_ASAP7_75t_L g761 ( .A(n_122), .Y(n_761) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND3x1_ASAP7_75t_L g123 ( .A(n_124), .B(n_356), .C(n_421), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_310), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_255), .B(n_283), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_218), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_166), .Y(n_127) );
AOI21xp33_ASAP7_75t_L g357 ( .A1(n_128), .A2(n_358), .B(n_369), .Y(n_357) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_128), .B(n_299), .Y(n_392) );
AND2x2_ASAP7_75t_L g407 ( .A(n_128), .B(n_408), .Y(n_407) );
OR2x6_ASAP7_75t_L g417 ( .A(n_128), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g419 ( .A(n_128), .B(n_409), .Y(n_419) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g293 ( .A(n_129), .Y(n_293) );
AND2x2_ASAP7_75t_L g306 ( .A(n_129), .B(n_307), .Y(n_306) );
INVx4_ASAP7_75t_L g325 ( .A(n_129), .Y(n_325) );
AND2x2_ASAP7_75t_L g328 ( .A(n_129), .B(n_244), .Y(n_328) );
NOR2x1_ASAP7_75t_SL g331 ( .A(n_129), .B(n_259), .Y(n_331) );
AND2x4_ASAP7_75t_L g343 ( .A(n_129), .B(n_341), .Y(n_343) );
OR2x2_ASAP7_75t_L g353 ( .A(n_129), .B(n_225), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_129), .B(n_365), .Y(n_370) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_135), .Y(n_129) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_131), .A2(n_179), .B1(n_185), .B2(n_186), .Y(n_178) );
INVx3_ASAP7_75t_L g186 ( .A(n_131), .Y(n_186) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_132), .B(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx4f_ASAP7_75t_L g170 ( .A(n_133), .Y(n_170) );
AND2x4_ASAP7_75t_L g164 ( .A(n_134), .B(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_134), .B(n_165), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_158), .B(n_164), .Y(n_135) );
INVxp67_ASAP7_75t_L g191 ( .A(n_137), .Y(n_191) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_143), .Y(n_137) );
NOR2x1p5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
INVx1_ASAP7_75t_L g204 ( .A(n_140), .Y(n_204) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OR2x6_ASAP7_75t_L g148 ( .A(n_141), .B(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g268 ( .A(n_142), .B(n_152), .Y(n_268) );
AND2x6_ASAP7_75t_L g481 ( .A(n_143), .B(n_163), .Y(n_481) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
INVx2_ASAP7_75t_L g149 ( .A(n_144), .Y(n_149) );
AND2x4_ASAP7_75t_L g271 ( .A(n_144), .B(n_154), .Y(n_271) );
HB1xp67_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_150), .C(n_156), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_SL g172 ( .A1(n_148), .A2(n_156), .B(n_173), .C(n_174), .Y(n_172) );
INVxp67_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_148), .A2(n_156), .B(n_213), .C(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g230 ( .A1(n_148), .A2(n_156), .B(n_231), .C(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g254 ( .A(n_148), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_148), .A2(n_183), .B1(n_263), .B2(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g160 ( .A(n_149), .B(n_161), .Y(n_160) );
INVxp33_ASAP7_75t_L g203 ( .A(n_149), .Y(n_203) );
INVx1_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
AND2x4_ASAP7_75t_L g482 ( .A(n_151), .B(n_157), .Y(n_482) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_154), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_156), .A2(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_156), .B(n_164), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_156), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_156), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_156), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_156), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_156), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_156), .A2(n_535), .B(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_156), .A2(n_560), .B(n_561), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_156), .A2(n_576), .B(n_577), .Y(n_575) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_157), .Y(n_184) );
INVx1_ASAP7_75t_L g193 ( .A(n_159), .Y(n_193) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_162), .Y(n_159) );
INVx1_ASAP7_75t_L g247 ( .A(n_160), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_162), .Y(n_248) );
BUFx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_164), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_SL g556 ( .A(n_164), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_164), .A2(n_573), .B(n_574), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_166), .A2(n_299), .B1(n_394), .B2(n_395), .Y(n_393) );
INVx1_ASAP7_75t_SL g437 ( .A(n_166), .Y(n_437) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_194), .Y(n_166) );
INVx2_ASAP7_75t_L g368 ( .A(n_167), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_167), .B(n_314), .Y(n_440) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_176), .Y(n_167) );
BUFx3_ASAP7_75t_L g286 ( .A(n_168), .Y(n_286) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g279 ( .A(n_169), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_169), .B(n_196), .Y(n_301) );
AND2x4_ASAP7_75t_L g318 ( .A(n_169), .B(n_319), .Y(n_318) );
INVxp67_ASAP7_75t_L g334 ( .A(n_169), .Y(n_334) );
INVx2_ASAP7_75t_L g391 ( .A(n_169), .Y(n_391) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_175), .Y(n_169) );
INVx2_ASAP7_75t_SL g197 ( .A(n_170), .Y(n_197) );
AND2x2_ASAP7_75t_L g309 ( .A(n_176), .B(n_275), .Y(n_309) );
NOR2xp67_ASAP7_75t_L g355 ( .A(n_176), .B(n_278), .Y(n_355) );
AND2x2_ASAP7_75t_L g374 ( .A(n_176), .B(n_278), .Y(n_374) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g236 ( .A(n_177), .Y(n_236) );
INVx1_ASAP7_75t_L g317 ( .A(n_177), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_177), .B(n_208), .Y(n_336) );
AND2x4_ASAP7_75t_L g390 ( .A(n_177), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_187), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_186), .A2(n_209), .B(n_215), .Y(n_208) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_186), .A2(n_209), .B(n_215), .Y(n_278) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_186), .A2(n_491), .B(n_497), .Y(n_490) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_186), .A2(n_512), .B(n_518), .Y(n_511) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_186), .A2(n_512), .B(n_518), .Y(n_545) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_186), .A2(n_491), .B(n_497), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_187) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g349 ( .A(n_194), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_194), .B(n_407), .Y(n_406) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_207), .Y(n_194) );
AND2x2_ASAP7_75t_L g333 ( .A(n_195), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g373 ( .A(n_195), .Y(n_373) );
AND2x2_ASAP7_75t_L g378 ( .A(n_195), .B(n_278), .Y(n_378) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_196), .B(n_208), .Y(n_238) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_206), .Y(n_196) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_197), .A2(n_198), .B(n_206), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_199), .B(n_205), .Y(n_198) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g314 ( .A(n_207), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_207), .B(n_286), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_207), .B(n_236), .Y(n_453) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_208), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_216), .Y(n_226) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_216), .A2(n_480), .B(n_486), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_216), .A2(n_525), .B(n_526), .Y(n_524) );
OA21x2_ASAP7_75t_L g625 ( .A1(n_216), .A2(n_480), .B(n_486), .Y(n_625) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OAI21xp33_ASAP7_75t_SL g218 ( .A1(n_219), .A2(n_234), .B(n_239), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_221), .B(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g291 ( .A(n_222), .Y(n_291) );
AND2x2_ASAP7_75t_L g305 ( .A(n_222), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g339 ( .A(n_222), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g405 ( .A(n_222), .B(n_323), .Y(n_405) );
NOR3xp33_ASAP7_75t_L g451 ( .A(n_222), .B(n_452), .C(n_453), .Y(n_451) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_223), .Y(n_282) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_225), .B(n_259), .Y(n_304) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_225), .Y(n_315) );
AND2x2_ASAP7_75t_L g360 ( .A(n_225), .B(n_258), .Y(n_360) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_225), .Y(n_383) );
INVx1_ASAP7_75t_L g400 ( .A(n_225), .Y(n_400) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_233), .Y(n_225) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_226), .A2(n_532), .B(n_538), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g442 ( .A(n_234), .Y(n_442) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_235), .B(n_313), .Y(n_414) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g276 ( .A(n_236), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AOI211x1_ASAP7_75t_L g310 ( .A1(n_240), .A2(n_311), .B(n_320), .C(n_337), .Y(n_310) );
INVx2_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_SL g303 ( .A(n_241), .B(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g363 ( .A(n_241), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g299 ( .A(n_243), .B(n_258), .Y(n_299) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x4_ASAP7_75t_L g257 ( .A(n_244), .B(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_244), .Y(n_324) );
INVx1_ASAP7_75t_L g341 ( .A(n_244), .Y(n_341) );
AND2x2_ASAP7_75t_L g409 ( .A(n_244), .B(n_259), .Y(n_409) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
NOR3xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .C(n_249), .Y(n_246) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_273), .B(n_280), .Y(n_255) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_256), .B(n_325), .Y(n_428) );
INVx2_ASAP7_75t_L g460 ( .A(n_256), .Y(n_460) );
INVx4_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g292 ( .A(n_257), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g365 ( .A(n_258), .Y(n_365) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B(n_272), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B1(n_269), .B2(n_270), .Y(n_265) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
OR2x2_ASAP7_75t_L g367 ( .A(n_274), .B(n_368), .Y(n_367) );
NAND2x1_ASAP7_75t_SL g389 ( .A(n_274), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g289 ( .A(n_275), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g319 ( .A(n_275), .Y(n_319) );
INVx1_ASAP7_75t_L g443 ( .A(n_276), .Y(n_443) );
AND2x2_ASAP7_75t_L g308 ( .A(n_277), .B(n_309), .Y(n_308) );
NOR2x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx2_ASAP7_75t_L g290 ( .A(n_278), .Y(n_290) );
INVxp33_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g347 ( .A(n_282), .B(n_340), .Y(n_347) );
OAI211xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .B(n_294), .C(n_302), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g371 ( .A(n_285), .B(n_372), .Y(n_371) );
NOR2xp67_ASAP7_75t_SL g376 ( .A(n_285), .B(n_377), .Y(n_376) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_286), .B(n_373), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_288), .B(n_292), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
AND2x2_ASAP7_75t_L g420 ( .A(n_289), .B(n_390), .Y(n_420) );
AOI222xp33_ASAP7_75t_L g438 ( .A1(n_292), .A2(n_439), .B1(n_441), .B2(n_444), .C1(n_445), .C2(n_448), .Y(n_438) );
INVx1_ASAP7_75t_L g402 ( .A(n_293), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_300), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_298), .Y(n_329) );
AND2x4_ASAP7_75t_SL g364 ( .A(n_298), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g418 ( .A(n_299), .Y(n_418) );
AND2x2_ASAP7_75t_L g463 ( .A(n_299), .B(n_315), .Y(n_463) );
AND2x2_ASAP7_75t_L g344 ( .A(n_300), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g457 ( .A(n_301), .B(n_336), .Y(n_457) );
OAI21xp33_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_305), .B(n_308), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_303), .A2(n_323), .B(n_364), .Y(n_424) );
AND2x2_ASAP7_75t_L g448 ( .A(n_304), .B(n_325), .Y(n_448) );
NOR2xp33_ASAP7_75t_SL g458 ( .A(n_304), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g396 ( .A(n_307), .Y(n_396) );
NOR2x1_ASAP7_75t_L g401 ( .A(n_307), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g431 ( .A(n_309), .Y(n_431) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_316), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AND2x2_ASAP7_75t_L g434 ( .A(n_314), .B(n_318), .Y(n_434) );
BUFx2_ASAP7_75t_L g322 ( .A(n_315), .Y(n_322) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g345 ( .A(n_317), .Y(n_345) );
INVx2_ASAP7_75t_L g351 ( .A(n_317), .Y(n_351) );
AND2x2_ASAP7_75t_L g387 ( .A(n_317), .B(n_378), .Y(n_387) );
AND2x4_ASAP7_75t_L g354 ( .A(n_318), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g394 ( .A(n_318), .B(n_351), .Y(n_394) );
AND2x2_ASAP7_75t_L g445 ( .A(n_318), .B(n_446), .Y(n_445) );
AOI31xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_326), .A3(n_330), .B(n_332), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g342 ( .A(n_322), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_SL g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x4_ASAP7_75t_L g340 ( .A(n_325), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_328), .A2(n_380), .B1(n_411), .B2(n_414), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_328), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g465 ( .A(n_328), .B(n_381), .Y(n_465) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g380 ( .A(n_331), .B(n_381), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
AND2x2_ASAP7_75t_L g403 ( .A(n_333), .B(n_374), .Y(n_403) );
INVx1_ASAP7_75t_L g413 ( .A(n_335), .Y(n_413) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_346), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g436 ( .A(n_339), .Y(n_436) );
AND2x2_ASAP7_75t_L g444 ( .A(n_340), .B(n_396), .Y(n_444) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_340), .Y(n_450) );
AND2x2_ASAP7_75t_L g395 ( .A(n_343), .B(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_348), .B1(n_352), .B2(n_354), .Y(n_346) );
NOR2xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_350), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_349), .A2(n_368), .B1(n_462), .B2(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g361 ( .A(n_354), .Y(n_361) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_384), .Y(n_356) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OAI21xp33_ASAP7_75t_L g362 ( .A1(n_360), .A2(n_363), .B(n_366), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_363), .A2(n_387), .B1(n_388), .B2(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_375), .B2(n_379), .Y(n_369) );
INVx1_ASAP7_75t_L g404 ( .A(n_372), .Y(n_404) );
NAND2x1p5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g384 ( .A(n_385), .B(n_397), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_393), .Y(n_385) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
NAND2xp33_ASAP7_75t_SL g439 ( .A(n_389), .B(n_440), .Y(n_439) );
INVx3_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
INVx3_ASAP7_75t_L g426 ( .A(n_394), .Y(n_426) );
INVxp67_ASAP7_75t_L g455 ( .A(n_395), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g397 ( .A(n_398), .B(n_406), .C(n_410), .D(n_415), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_403), .B1(n_404), .B2(n_405), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
AND2x2_ASAP7_75t_L g408 ( .A(n_400), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g456 ( .A(n_404), .Y(n_456) );
NAND2xp33_ASAP7_75t_SL g411 ( .A(n_412), .B(n_413), .Y(n_411) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_419), .B(n_420), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND3x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_438), .C(n_449), .Y(n_421) );
AOI221x1_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_427), .B2(n_429), .C(n_435), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp33_ASAP7_75t_SL g429 ( .A(n_430), .B(n_433), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
NAND2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AOI211xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_454), .C(n_461), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_454) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_467), .Y(n_760) );
CKINVDCx11_ASAP7_75t_R g467 ( .A(n_468), .Y(n_467) );
CKINVDCx6p67_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
CKINVDCx11_ASAP7_75t_R g758 ( .A(n_470), .Y(n_758) );
INVx3_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g759 ( .A(n_473), .Y(n_759) );
NAND4xp75_ASAP7_75t_L g473 ( .A(n_474), .B(n_665), .C(n_705), .D(n_734), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_627), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_584), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_519), .B(n_539), .Y(n_476) );
AND2x2_ASAP7_75t_SL g477 ( .A(n_478), .B(n_487), .Y(n_477) );
AND2x4_ASAP7_75t_L g583 ( .A(n_478), .B(n_544), .Y(n_583) );
INVx1_ASAP7_75t_SL g636 ( .A(n_478), .Y(n_636) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_478), .A2(n_672), .B(n_675), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_SL g675 ( .A1(n_478), .A2(n_676), .B(n_677), .C(n_678), .Y(n_675) );
NAND2x1_ASAP7_75t_L g716 ( .A(n_478), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_478), .B(n_677), .Y(n_738) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g542 ( .A(n_479), .Y(n_542) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_479), .Y(n_615) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_498), .Y(n_487) );
AND2x2_ASAP7_75t_L g607 ( .A(n_488), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g688 ( .A(n_488), .B(n_544), .Y(n_688) );
INVx1_ASAP7_75t_L g748 ( .A(n_488), .Y(n_748) );
BUFx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g592 ( .A(n_489), .B(n_510), .Y(n_592) );
AND2x2_ASAP7_75t_L g717 ( .A(n_489), .B(n_511), .Y(n_717) );
AND2x2_ASAP7_75t_L g722 ( .A(n_489), .B(n_682), .Y(n_722) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVxp67_ASAP7_75t_L g598 ( .A(n_490), .Y(n_598) );
BUFx3_ASAP7_75t_L g631 ( .A(n_490), .Y(n_631) );
AND2x2_ASAP7_75t_L g677 ( .A(n_490), .B(n_511), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_496), .Y(n_491) );
AND2x2_ASAP7_75t_L g662 ( .A(n_498), .B(n_541), .Y(n_662) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
AND2x4_ASAP7_75t_L g544 ( .A(n_499), .B(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g654 ( .A(n_499), .B(n_638), .Y(n_654) );
AND2x2_ASAP7_75t_SL g697 ( .A(n_499), .B(n_625), .Y(n_697) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g633 ( .A(n_500), .Y(n_633) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g594 ( .A(n_501), .Y(n_594) );
OAI21x1_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_504), .B(n_508), .Y(n_501) );
INVx1_ASAP7_75t_L g509 ( .A(n_503), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_510), .B(n_594), .Y(n_597) );
AND2x2_ASAP7_75t_L g682 ( .A(n_510), .B(n_625), .Y(n_682) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g679 ( .A(n_511), .B(n_542), .Y(n_679) );
AND2x2_ASAP7_75t_L g699 ( .A(n_511), .B(n_625), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_513), .B(n_517), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_519), .B(n_588), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_519), .A2(n_711), .B1(n_712), .B2(n_713), .C(n_715), .Y(n_710) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI332xp33_ASAP7_75t_L g744 ( .A1(n_520), .A2(n_604), .A3(n_611), .B1(n_670), .B2(n_745), .B3(n_746), .C1(n_747), .C2(n_749), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
AND2x2_ASAP7_75t_L g550 ( .A(n_521), .B(n_531), .Y(n_550) );
AND2x2_ASAP7_75t_L g567 ( .A(n_521), .B(n_568), .Y(n_567) );
INVx4_ASAP7_75t_L g579 ( .A(n_521), .Y(n_579) );
AND2x2_ASAP7_75t_SL g639 ( .A(n_521), .B(n_580), .Y(n_639) );
INVx5_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NOR2x1_ASAP7_75t_SL g601 ( .A(n_522), .B(n_568), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_522), .B(n_530), .Y(n_605) );
AND2x2_ASAP7_75t_L g612 ( .A(n_522), .B(n_531), .Y(n_612) );
BUFx2_ASAP7_75t_L g647 ( .A(n_522), .Y(n_647) );
AND2x2_ASAP7_75t_L g702 ( .A(n_522), .B(n_571), .Y(n_702) );
OR2x6_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
OR2x2_ASAP7_75t_L g570 ( .A(n_530), .B(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g580 ( .A(n_530), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g620 ( .A(n_530), .Y(n_620) );
AND2x2_ASAP7_75t_L g690 ( .A(n_530), .B(n_589), .Y(n_690) );
AND2x2_ASAP7_75t_L g703 ( .A(n_530), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_530), .B(n_704), .Y(n_721) );
INVx4_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_531), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_537), .Y(n_532) );
OAI32xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_546), .A3(n_551), .B1(n_565), .B2(n_582), .Y(n_539) );
INVx2_ASAP7_75t_L g648 ( .A(n_540), .Y(n_648) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx1_ASAP7_75t_L g659 ( .A(n_541), .Y(n_659) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g593 ( .A(n_542), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g726 ( .A(n_542), .B(n_631), .Y(n_726) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g638 ( .A(n_545), .Y(n_638) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVx2_ASAP7_75t_L g626 ( .A(n_548), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_548), .B(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_SL g637 ( .A(n_549), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g714 ( .A(n_549), .Y(n_714) );
AND2x2_ASAP7_75t_L g732 ( .A(n_549), .B(n_594), .Y(n_732) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NOR2xp67_ASAP7_75t_SL g676 ( .A(n_552), .B(n_605), .Y(n_676) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_553), .B(n_587), .Y(n_674) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g750 ( .A(n_554), .B(n_620), .Y(n_750) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g581 ( .A(n_555), .Y(n_581) );
INVx2_ASAP7_75t_L g622 ( .A(n_555), .Y(n_622) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B(n_563), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_556), .B(n_564), .Y(n_563) );
AO21x2_ASAP7_75t_L g568 ( .A1(n_556), .A2(n_557), .B(n_563), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_562), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_578), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_566), .B(n_624), .Y(n_709) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
AND3x2_ASAP7_75t_L g664 ( .A(n_567), .B(n_611), .C(n_620), .Y(n_664) );
AND2x2_ASAP7_75t_L g588 ( .A(n_568), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_568), .B(n_571), .Y(n_645) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g599 ( .A(n_570), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g589 ( .A(n_571), .Y(n_589) );
INVx1_ASAP7_75t_L g604 ( .A(n_571), .Y(n_604) );
BUFx3_ASAP7_75t_L g611 ( .A(n_571), .Y(n_611) );
AND2x2_ASAP7_75t_L g621 ( .A(n_571), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AND2x4_ASAP7_75t_L g630 ( .A(n_579), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_579), .B(n_589), .Y(n_673) );
AND2x2_ASAP7_75t_L g629 ( .A(n_580), .B(n_604), .Y(n_629) );
INVx2_ASAP7_75t_L g656 ( .A(n_580), .Y(n_656) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AOI211xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_590), .B(n_595), .C(n_616), .Y(n_584) );
OAI21xp5_ASAP7_75t_L g736 ( .A1(n_585), .A2(n_712), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_588), .B(n_647), .Y(n_646) );
AOI211xp5_ASAP7_75t_SL g666 ( .A1(n_588), .A2(n_667), .B(n_671), .C(n_680), .Y(n_666) );
AND2x2_ASAP7_75t_L g652 ( .A(n_589), .B(n_612), .Y(n_652) );
OR2x2_ASAP7_75t_L g655 ( .A(n_589), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_592), .B(n_697), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_593), .B(n_638), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_593), .A2(n_619), .B1(n_699), .B2(n_702), .C(n_708), .Y(n_707) );
AND2x4_ASAP7_75t_L g624 ( .A(n_594), .B(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g670 ( .A(n_594), .B(n_625), .Y(n_670) );
OAI221xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_599), .B1(n_602), .B2(n_606), .C(n_609), .Y(n_595) );
AND2x2_ASAP7_75t_L g741 ( .A(n_596), .B(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g608 ( .A(n_597), .Y(n_608) );
INVx1_ASAP7_75t_L g694 ( .A(n_598), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_599), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g613 ( .A(n_601), .B(n_604), .Y(n_613) );
AND2x2_ASAP7_75t_L g689 ( .A(n_601), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g614 ( .A(n_608), .B(n_615), .Y(n_614) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_613), .B(n_614), .Y(n_609) );
INVx1_ASAP7_75t_L g733 ( .A(n_610), .Y(n_733) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g712 ( .A(n_611), .B(n_639), .Y(n_712) );
AND2x2_ASAP7_75t_SL g685 ( .A(n_612), .B(n_621), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_623), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_617), .A2(n_651), .B1(n_654), .B2(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g723 ( .A(n_617), .Y(n_723) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g643 ( .A(n_620), .Y(n_643) );
INVx1_ASAP7_75t_L g704 ( .A(n_622), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_624), .B(n_626), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g745 ( .A(n_624), .B(n_694), .Y(n_745) );
AND2x2_ASAP7_75t_L g713 ( .A(n_625), .B(n_714), .Y(n_713) );
OAI211xp5_ASAP7_75t_L g706 ( .A1(n_626), .A2(n_707), .B(n_710), .C(n_718), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_649), .Y(n_627) );
AOI322xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .A3(n_632), .B1(n_634), .B2(n_639), .C1(n_640), .C2(n_648), .Y(n_628) );
CKINVDCx16_ASAP7_75t_R g746 ( .A(n_630), .Y(n_746) );
AND2x2_ASAP7_75t_L g696 ( .A(n_631), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g730 ( .A(n_631), .Y(n_730) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_SL g681 ( .A(n_633), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_633), .B(n_679), .Y(n_687) );
AND2x2_ASAP7_75t_L g711 ( .A(n_633), .B(n_677), .Y(n_711) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g683 ( .A(n_637), .Y(n_683) );
NAND2xp33_ASAP7_75t_SL g640 ( .A(n_641), .B(n_646), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI221xp5_ASAP7_75t_SL g686 ( .A1(n_642), .A2(n_687), .B1(n_688), .B2(n_689), .C(n_691), .Y(n_686) );
AND2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVxp67_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g753 ( .A(n_645), .Y(n_753) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B(n_653), .C(n_657), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g728 ( .A(n_652), .Y(n_728) );
INVx1_ASAP7_75t_L g660 ( .A(n_654), .Y(n_660) );
OR2x2_ASAP7_75t_L g747 ( .A(n_654), .B(n_748), .Y(n_747) );
INVx2_ASAP7_75t_SL g743 ( .A(n_655), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B(n_663), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_659), .B(n_677), .Y(n_754) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_686), .Y(n_665) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_669), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
OR2x2_ASAP7_75t_L g720 ( .A(n_673), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI21xp33_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_683), .B(n_684), .Y(n_680) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AOI31xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .A3(n_698), .B(n_700), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_697), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_722), .B1(n_723), .B2(n_724), .C(n_727), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_731), .B2(n_733), .Y(n_727) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
NOR3xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_744), .C(n_751), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_736), .B(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_743), .Y(n_739) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OAI22x1_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_759), .B1(n_760), .B2(n_761), .Y(n_757) );
INVx3_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_765), .B(n_768), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g784 ( .A(n_775), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
AND2x4_ASAP7_75t_SL g776 ( .A(n_777), .B(n_778), .Y(n_776) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
endmodule