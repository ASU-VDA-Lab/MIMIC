module fake_jpeg_22633_n_304 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_SL g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_26),
.B1(n_40),
.B2(n_20),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_26),
.B1(n_20),
.B2(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_26),
.B1(n_34),
.B2(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_30),
.B1(n_26),
.B2(n_33),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_23),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_17),
.B1(n_42),
.B2(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_30),
.B1(n_37),
.B2(n_42),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_59),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_33),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_36),
.B1(n_24),
.B2(n_28),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_35),
.B1(n_37),
.B2(n_40),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_69),
.A2(n_64),
.B1(n_48),
.B2(n_57),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_32),
.B(n_22),
.C(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_70),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_75),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_72),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_77),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_83),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_39),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_37),
.C(n_19),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_27),
.B1(n_37),
.B2(n_39),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_95),
.Y(n_122)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_99),
.B(n_101),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_104),
.B(n_107),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_53),
.B(n_40),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_116),
.B1(n_77),
.B2(n_37),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_24),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_24),
.Y(n_111)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_37),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_41),
.Y(n_143)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_118),
.B1(n_36),
.B2(n_92),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_80),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_117),
.A2(n_81),
.B1(n_36),
.B2(n_29),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_119),
.Y(n_123)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_18),
.Y(n_121)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_110),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_132),
.B1(n_133),
.B2(n_149),
.Y(n_170)
);

XOR2x2_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_114),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_143),
.B(n_146),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_134),
.B1(n_150),
.B2(n_117),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_81),
.B1(n_82),
.B2(n_85),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_120),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_87),
.B1(n_69),
.B2(n_77),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_103),
.B(n_106),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_69),
.B(n_43),
.C(n_41),
.D(n_49),
.Y(n_139)
);

AOI221xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_116),
.B1(n_106),
.B2(n_112),
.C(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_107),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_19),
.B(n_21),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_41),
.B1(n_43),
.B2(n_36),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_91),
.B1(n_36),
.B2(n_43),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_45),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_180),
.B(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_155),
.B(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_159),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_136),
.A2(n_97),
.B(n_113),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_176),
.B(n_147),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_177),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_161),
.A2(n_126),
.B1(n_133),
.B2(n_98),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_102),
.A3(n_109),
.B1(n_110),
.B2(n_108),
.C1(n_122),
.C2(n_99),
.Y(n_162)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_169),
.B1(n_146),
.B2(n_132),
.C(n_143),
.Y(n_183)
);

BUFx24_ASAP7_75t_SL g163 ( 
.A(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_168),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_173),
.C(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_112),
.Y(n_172)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_116),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_112),
.C(n_106),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_145),
.C(n_141),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_136),
.A2(n_106),
.B(n_76),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_31),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_88),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_98),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_130),
.A2(n_19),
.B(n_21),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_138),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_96),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_156),
.A2(n_157),
.B1(n_130),
.B2(n_181),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_182),
.A2(n_203),
.B1(n_167),
.B2(n_175),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_183),
.B(n_194),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_184),
.A2(n_29),
.B(n_21),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_170),
.A2(n_128),
.B1(n_144),
.B2(n_139),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_200),
.B1(n_202),
.B2(n_155),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_176),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_187),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_205),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_123),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_170),
.A2(n_92),
.B1(n_119),
.B2(n_74),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_123),
.B1(n_96),
.B2(n_88),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_154),
.A2(n_28),
.B1(n_18),
.B2(n_29),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_72),
.Y(n_226)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_153),
.C(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_209),
.C(n_216),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_153),
.C(n_160),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_217),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_225),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_172),
.B1(n_167),
.B2(n_166),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_178),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_220),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_164),
.C(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_185),
.A2(n_158),
.B1(n_159),
.B2(n_180),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_177),
.B1(n_96),
.B2(n_18),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_203),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_177),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_46),
.C(n_45),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_223),
.C(n_229),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_222),
.B(n_202),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_45),
.C(n_62),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_227),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_28),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_8),
.B(n_15),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_62),
.C(n_43),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_43),
.C(n_41),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_189),
.C(n_188),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_237),
.Y(n_259)
);

AOI31xp67_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_187),
.A3(n_191),
.B(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_239),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_205),
.B(n_204),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_209),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_246),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_182),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_189),
.Y(n_241)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_241),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_190),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_249),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_250),
.C(n_216),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_231),
.A2(n_22),
.B(n_31),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_8),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_208),
.B(n_72),
.C(n_1),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_256),
.C(n_238),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_220),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_222),
.C(n_223),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_229),
.B1(n_230),
.B2(n_2),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_258),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_234),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_253),
.B1(n_255),
.B2(n_257),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_13),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_250),
.B(n_240),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_12),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_242),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_245),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_266),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_258),
.B(n_262),
.C(n_259),
.Y(n_280)
);

A2O1A1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_254),
.A2(n_237),
.B(n_246),
.C(n_242),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_276),
.B(n_259),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_9),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_236),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_272),
.C(n_273),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_240),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_11),
.B(n_10),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_274),
.A2(n_11),
.B(n_10),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_0),
.C(n_2),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_11),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_280),
.B(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_3),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_262),
.B(n_10),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_276),
.C(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_284),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_0),
.B(n_2),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_0),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_286),
.A2(n_268),
.B1(n_4),
.B2(n_5),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_289),
.C(n_3),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_285),
.A2(n_268),
.B1(n_270),
.B2(n_5),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_291),
.B(n_294),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_3),
.C(n_4),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_290),
.A2(n_284),
.B1(n_286),
.B2(n_6),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_7),
.B1(n_291),
.B2(n_290),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_3),
.B(n_5),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_7),
.B(n_299),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_293),
.C(n_6),
.Y(n_300)
);

AO21x2_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_296),
.Y(n_304)
);


endmodule