module fake_jpeg_1140_n_178 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_54),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_1),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_78),
.Y(n_85)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_42),
.B1(n_58),
.B2(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_49),
.B1(n_48),
.B2(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_55),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_62),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_88),
.B(n_93),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_84),
.B(n_92),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_68),
.B1(n_42),
.B2(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_89),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_59),
.B1(n_47),
.B2(n_43),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_91),
.B(n_46),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_65),
.B1(n_47),
.B2(n_59),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_49),
.B(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_50),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_79),
.A2(n_46),
.B(n_45),
.C(n_52),
.Y(n_94)
);

BUFx8_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_45),
.B(n_2),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_98),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_60),
.Y(n_98)
);

HAxp5_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_57),
.CON(n_99),
.SN(n_99)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_98),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_75),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_116),
.Y(n_134)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_114),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_81),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_97),
.C(n_87),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_136),
.C(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_129),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_94),
.B(n_76),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_102),
.B(n_107),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_104),
.B1(n_99),
.B2(n_108),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_89),
.B1(n_76),
.B2(n_3),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_1),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_4),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_111),
.B1(n_109),
.B2(n_105),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_31),
.C(n_30),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_137),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_147),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_141),
.B(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

OAI22x1_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_23),
.B1(n_22),
.B2(n_12),
.Y(n_161)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_151),
.B1(n_153),
.B2(n_128),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_28),
.C(n_27),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_149),
.C(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_120),
.B(n_123),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_24),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_123),
.C(n_135),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_122),
.B(n_119),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_7),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_145),
.C(n_21),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_161),
.B1(n_162),
.B2(n_14),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_157),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_138),
.C(n_147),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_165),
.Y(n_169)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_143),
.A3(n_149),
.B1(n_142),
.B2(n_137),
.C1(n_18),
.C2(n_14),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_168),
.C(n_158),
.Y(n_171)
);

OA21x2_ASAP7_75t_SL g170 ( 
.A1(n_167),
.A2(n_161),
.B(n_157),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_15),
.B(n_16),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.C(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_169),
.B(n_163),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_172),
.A2(n_173),
.B1(n_171),
.B2(n_166),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_15),
.B(n_16),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_17),
.C(n_19),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_17),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_19),
.Y(n_178)
);


endmodule