module fake_netlist_1_5875_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
BUFx8_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_9), .B(n_10), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
AND2x4_ASAP7_75t_SL g17 ( .A(n_13), .B(n_0), .Y(n_17) );
CKINVDCx16_ASAP7_75t_R g18 ( .A(n_11), .Y(n_18) );
AO21x2_ASAP7_75t_L g19 ( .A1(n_16), .A2(n_14), .B(n_11), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_15), .B(n_12), .Y(n_20) );
OR2x2_ASAP7_75t_L g21 ( .A(n_19), .B(n_18), .Y(n_21) );
NOR2x1_ASAP7_75t_L g22 ( .A(n_19), .B(n_18), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_19), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_19), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_20), .Y(n_25) );
AOI322xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_12), .A3(n_2), .B1(n_3), .B2(n_4), .C1(n_5), .C2(n_6), .Y(n_26) );
OAI21xp33_ASAP7_75t_SL g27 ( .A1(n_25), .A2(n_24), .B(n_20), .Y(n_27) );
OAI21xp33_ASAP7_75t_SL g28 ( .A1(n_25), .A2(n_20), .B(n_12), .Y(n_28) );
OAI221xp5_ASAP7_75t_SL g29 ( .A1(n_28), .A2(n_26), .B1(n_2), .B2(n_3), .C(n_4), .Y(n_29) );
AOI321xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_1), .A3(n_5), .B1(n_6), .B2(n_7), .C(n_8), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
HB1xp67_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
AOI21xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_7), .B(n_8), .Y(n_33) );
OAI21xp5_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_31), .B(n_32), .Y(n_34) );
endmodule