module fake_jpeg_28136_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_39),
.Y(n_61)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_46),
.Y(n_69)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_0),
.Y(n_65)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_16),
.B(n_0),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_28),
.B1(n_17),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_57),
.B1(n_66),
.B2(n_71),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_17),
.B1(n_28),
.B2(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_75),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_17),
.B1(n_28),
.B2(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_28),
.B1(n_18),
.B2(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_76),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_38),
.A2(n_25),
.B1(n_24),
.B2(n_18),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_43),
.B(n_45),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_24),
.B1(n_27),
.B2(n_35),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_78),
.B(n_82),
.Y(n_141)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_46),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_69),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_44),
.B(n_37),
.C(n_46),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_89),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_37),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_47),
.Y(n_90)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_91),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_97),
.B(n_102),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_54),
.B(n_19),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_19),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_35),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_111),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_22),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_22),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_72),
.C(n_58),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_15),
.Y(n_111)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_22),
.Y(n_114)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_31),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_52),
.Y(n_116)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_45),
.B1(n_39),
.B2(n_48),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_137),
.B1(n_107),
.B2(n_106),
.Y(n_160)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_136),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_48),
.Y(n_164)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_39),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_32),
.Y(n_171)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_45),
.B1(n_48),
.B2(n_16),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_81),
.B(n_53),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_103),
.B(n_110),
.Y(n_152)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_144),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_79),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_143),
.B(n_85),
.Y(n_161)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_83),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_148),
.B(n_154),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_83),
.B(n_101),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_151),
.A2(n_152),
.B(n_26),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_109),
.B1(n_95),
.B2(n_105),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_163),
.B1(n_168),
.B2(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_91),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_155),
.B(n_156),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_90),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_167),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_146),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_107),
.B(n_113),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_159),
.A2(n_32),
.B(n_26),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_175),
.B1(n_128),
.B2(n_136),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_96),
.Y(n_162)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_181),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_138),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_126),
.B(n_20),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_87),
.B1(n_93),
.B2(n_86),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_118),
.A2(n_80),
.B1(n_86),
.B2(n_93),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_173),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_171),
.B(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_34),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_176),
.Y(n_210)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_80),
.B1(n_116),
.B2(n_29),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_34),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_23),
.Y(n_177)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_96),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

NAND2x1_ASAP7_75t_SL g213 ( 
.A(n_180),
.B(n_2),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_118),
.B(n_23),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_148),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_187),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_149),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_120),
.C(n_121),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_153),
.C(n_164),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_140),
.B1(n_130),
.B2(n_122),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_191),
.A2(n_198),
.B1(n_204),
.B2(n_208),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_150),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_192),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_122),
.B1(n_144),
.B2(n_142),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_181),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_163),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_96),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_206),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_48),
.B1(n_23),
.B2(n_29),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_203),
.B(n_152),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_23),
.B1(n_29),
.B2(n_31),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_20),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_159),
.A2(n_31),
.B1(n_26),
.B2(n_20),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_168),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_228),
.C(n_187),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_220),
.B(n_223),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_184),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_221),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_177),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_172),
.B(n_167),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_225),
.A2(n_229),
.B(n_4),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_227),
.A2(n_189),
.B1(n_207),
.B2(n_204),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_156),
.C(n_166),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_155),
.B(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_211),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_186),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_233),
.Y(n_254)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_178),
.Y(n_234)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

OAI32xp33_ASAP7_75t_L g236 ( 
.A1(n_196),
.A2(n_178),
.A3(n_11),
.B1(n_12),
.B2(n_7),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_208),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_10),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_238),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_10),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_242),
.C(n_246),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_183),
.C(n_185),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_190),
.C(n_200),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_200),
.C(n_197),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_260),
.C(n_235),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_195),
.B1(n_209),
.B2(n_188),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_219),
.B1(n_223),
.B2(n_233),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_259),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_219),
.A2(n_210),
.B1(n_213),
.B2(n_198),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_210),
.B1(n_207),
.B2(n_206),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_257),
.A2(n_262),
.B1(n_217),
.B2(n_221),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_3),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_3),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_15),
.C(n_9),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_261),
.A2(n_226),
.B(n_229),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_217),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_275),
.B1(n_263),
.B2(n_252),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_272),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_228),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_271),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_225),
.C(n_224),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_278),
.C(n_280),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_270),
.A2(n_254),
.B(n_253),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_218),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_246),
.B(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_220),
.B(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_261),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_215),
.B1(n_240),
.B2(n_230),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_215),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_231),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_250),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_289),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_253),
.C(n_243),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_293),
.C(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_259),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_288),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_262),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_292),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_263),
.A2(n_243),
.B1(n_244),
.B2(n_262),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_264),
.C(n_268),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_264),
.C(n_267),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_296),
.B(n_297),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_276),
.C(n_244),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_274),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_302),
.B(n_260),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_255),
.Y(n_303)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_283),
.B(n_265),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_270),
.B(n_251),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_309),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_304),
.A2(n_291),
.B1(n_266),
.B2(n_292),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_258),
.B1(n_9),
.B2(n_11),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_283),
.C(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_13),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_13),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_298),
.B(n_295),
.Y(n_315)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_295),
.B1(n_302),
.B2(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_317),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_314),
.Y(n_323)
);

AOI211xp5_ASAP7_75t_L g325 ( 
.A1(n_323),
.A2(n_324),
.B(n_321),
.C(n_309),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_320),
.A2(n_316),
.B(n_308),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_307),
.B(n_319),
.Y(n_326)
);

OAI321xp33_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_319),
.A3(n_13),
.B1(n_14),
.B2(n_5),
.C(n_4),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_4),
.B(n_5),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_5),
.B1(n_14),
.B2(n_250),
.Y(n_329)
);


endmodule