module fake_jpeg_17448_n_245 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_245);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_45),
.Y(n_62)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_52),
.B1(n_26),
.B2(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_56),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx12_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_53),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_28),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_59),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_76),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_23),
.B1(n_15),
.B2(n_16),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_33),
.B1(n_30),
.B2(n_37),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_73),
.B1(n_45),
.B2(n_41),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_72),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_24),
.B1(n_26),
.B2(n_19),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_79),
.B1(n_19),
.B2(n_15),
.Y(n_84)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

AOI22x1_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_37),
.B1(n_35),
.B2(n_29),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_34),
.C(n_22),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_13),
.C(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_41),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_40),
.B(n_23),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_77),
.B(n_27),
.Y(n_82)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_78),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_40),
.A2(n_19),
.B1(n_45),
.B2(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_76),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_84),
.B1(n_60),
.B2(n_78),
.Y(n_105)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_44),
.B1(n_30),
.B2(n_35),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_88),
.A2(n_94),
.B1(n_95),
.B2(n_68),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_98),
.C(n_99),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_93),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_29),
.B1(n_42),
.B2(n_38),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_42),
.B1(n_38),
.B2(n_21),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_60),
.B1(n_17),
.B2(n_14),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_74),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_100),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_48),
.C(n_51),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_48),
.C(n_51),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_16),
.B(n_15),
.C(n_23),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_62),
.A2(n_16),
.B(n_18),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_14),
.B(n_17),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_112),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_114),
.B1(n_126),
.B2(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_62),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_64),
.B1(n_78),
.B2(n_60),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_125),
.B1(n_80),
.B2(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

BUFx4f_ASAP7_75t_SL g117 ( 
.A(n_86),
.Y(n_117)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_69),
.C(n_59),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_127),
.C(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_84),
.Y(n_145)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_82),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_83),
.A2(n_68),
.B1(n_63),
.B2(n_38),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_48),
.C(n_51),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_133),
.B1(n_86),
.B2(n_115),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_81),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_136),
.C(n_139),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_135),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_102),
.B(n_100),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_144),
.B(n_119),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_89),
.C(n_87),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_88),
.Y(n_139)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_80),
.B1(n_100),
.B2(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_121),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_147),
.B(n_145),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_68),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_68),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_79),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_136),
.C(n_144),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_150),
.B(n_151),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_125),
.A3(n_120),
.B1(n_104),
.B2(n_118),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_118),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_166),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_134),
.B(n_132),
.C(n_131),
.Y(n_177)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_94),
.B1(n_126),
.B2(n_120),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_171),
.B1(n_117),
.B2(n_65),
.Y(n_185)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_169),
.B(n_14),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_137),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_168),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_133),
.A2(n_146),
.B1(n_142),
.B2(n_149),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_170),
.B1(n_106),
.B2(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_110),
.B(n_124),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_86),
.B1(n_106),
.B2(n_123),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_158),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_141),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_162),
.B1(n_161),
.B2(n_171),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_49),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_182),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_117),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_181),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_48),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_183),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_188),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_74),
.C(n_13),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_153),
.C(n_163),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_169),
.A2(n_17),
.B1(n_21),
.B2(n_7),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_187),
.C(n_183),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_172),
.B1(n_21),
.B2(n_13),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_165),
.C(n_166),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_197),
.C(n_180),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_181),
.A2(n_159),
.B1(n_155),
.B2(n_156),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_185),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_195),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_165),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_161),
.C(n_155),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_199),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_7),
.B(n_12),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_200),
.A2(n_174),
.B(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_208),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_206),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_183),
.C(n_186),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_177),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_209),
.A2(n_191),
.B1(n_193),
.B2(n_199),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_210),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_0),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_213),
.B1(n_198),
.B2(n_10),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_22),
.C(n_21),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_0),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_217),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_201),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_220),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_191),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_223),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_212),
.B(n_203),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_227),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_213),
.Y(n_225)
);

AOI31xp67_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_10),
.A3(n_12),
.B(n_5),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_22),
.C(n_3),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_216),
.A2(n_218),
.B1(n_223),
.B2(n_221),
.Y(n_228)
);

BUFx12_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_235),
.Y(n_237)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_230),
.A2(n_218),
.B(n_4),
.C(n_5),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_229),
.Y(n_239)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_234),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_22),
.Y(n_235)
);

OAI21x1_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_228),
.B(n_227),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_239),
.A2(n_233),
.B(n_232),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_236),
.C(n_234),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_242),
.B(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_237),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_237),
.Y(n_245)
);


endmodule