module real_jpeg_8170_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_315, n_6, n_316, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_315;
input n_6;
input n_316;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_2),
.A2(n_66),
.B1(n_67),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_2),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_139),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_139),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_139),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_3),
.A2(n_51),
.B1(n_66),
.B2(n_67),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_5),
.A2(n_61),
.B1(n_66),
.B2(n_67),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_61),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_61),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_31),
.B(n_64),
.C(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_6),
.B(n_31),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_6),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_65)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_43),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_9),
.A2(n_43),
.B1(n_66),
.B2(n_67),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_11),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_79),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_79),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_79),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_12),
.A2(n_31),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_12),
.B(n_31),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_12),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_12),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_12),
.A2(n_27),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_12),
.B(n_27),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_12),
.B(n_52),
.Y(n_167)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_12),
.A2(n_28),
.B(n_47),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_12),
.A2(n_40),
.B1(n_41),
.B2(n_123),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_13),
.A2(n_66),
.B1(n_67),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_13),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_98),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_98),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_98),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_14),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_14),
.A2(n_66),
.B1(n_67),
.B2(n_110),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_110),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_110),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_15),
.A2(n_66),
.B1(n_67),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_15),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_103),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_103),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_103),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_17),
.A2(n_35),
.B1(n_66),
.B2(n_67),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_86),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_84),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_71),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_53),
.B1(n_54),
.B2(n_70),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_25),
.A2(n_30),
.B1(n_57),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_25),
.A2(n_30),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_25),
.A2(n_30),
.B1(n_148),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_25),
.A2(n_30),
.B1(n_164),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_25),
.A2(n_30),
.B1(n_204),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_25),
.A2(n_30),
.B1(n_215),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_25),
.A2(n_30),
.B1(n_241),
.B2(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_25),
.A2(n_30),
.B1(n_83),
.B2(n_259),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_27),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_49)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_29),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_30),
.B(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_31),
.B(n_33),
.Y(n_152)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_32),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_44),
.B1(n_50),
.B2(n_52),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_45),
.B1(n_49),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_46),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_41),
.A2(n_46),
.B(n_123),
.C(n_186),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_44),
.A2(n_52),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_49),
.B1(n_60),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_45),
.A2(n_49),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_45),
.A2(n_49),
.B1(n_219),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_45),
.A2(n_49),
.B1(n_244),
.B2(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_45),
.A2(n_49),
.B1(n_78),
.B2(n_262),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.C(n_62),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_56),
.B1(n_62),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_59),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_62),
.A2(n_76),
.B1(n_81),
.B2(n_82),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_65),
.B(n_69),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_65),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_63),
.A2(n_65),
.B1(n_109),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_63),
.A2(n_65),
.B1(n_136),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_63),
.A2(n_65),
.B1(n_144),
.B2(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_63),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_63),
.A2(n_65),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_63),
.A2(n_65),
.B1(n_227),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_63),
.A2(n_65),
.B1(n_236),
.B2(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_63),
.A2(n_65),
.B1(n_69),
.B2(n_268),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_65),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_65),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_66),
.B(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_66),
.B(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_67),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.C(n_80),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_302),
.Y(n_307)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_77),
.C(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_77),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_77),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_80),
.B(n_307),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_299),
.A3(n_308),
.B1(n_311),
.B2(n_312),
.C(n_315),
.Y(n_86)
);

AOI321xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_252),
.A3(n_287),
.B1(n_293),
.B2(n_298),
.C(n_316),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_209),
.C(n_248),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_179),
.B(n_208),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_158),
.B(n_178),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_141),
.B(n_157),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_130),
.B(n_140),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_116),
.B(n_129),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_95),
.B(n_104),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_97),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_99),
.A2(n_100),
.B1(n_156),
.B2(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_120),
.B1(n_121),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_111),
.B2(n_115),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_115),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_108),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_124),
.B(n_128),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_122),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_121),
.B1(n_138),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_120),
.A2(n_121),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_120),
.A2(n_121),
.B1(n_190),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_120),
.A2(n_121),
.B1(n_224),
.B2(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_120),
.A2(n_121),
.B(n_234),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_132),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_133),
.B(n_142),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.CI(n_137),
.CON(n_133),
.SN(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_145),
.CI(n_149),
.CON(n_142),
.SN(n_142)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_147),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_154),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_160),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_171),
.B2(n_172),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_174),
.C(n_176),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_165),
.B1(n_166),
.B2(n_170),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_168),
.C(n_170),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_180),
.B(n_181),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_194),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_183),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_193),
.C(n_194),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_188),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_191),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_205),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_202),
.B2(n_203),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_202),
.C(n_205),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_207),
.Y(n_218)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_210),
.A2(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_229),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_211),
.B(n_229),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_222),
.C(n_228),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_221),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_216),
.B1(n_217),
.B2(n_220),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_214),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_SL g246 ( 
.A(n_216),
.B(n_220),
.C(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_228),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_225),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_246),
.B2(n_247),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_232),
.B(n_237),
.C(n_247),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_235),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_242),
.C(n_245),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_242),
.B1(n_243),
.B2(n_245),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_240),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_246),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_249),
.B(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_271),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_253),
.B(n_271),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_264),
.C(n_270),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_254),
.A2(n_255),
.B1(n_264),
.B2(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_260),
.C(n_263),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_258),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_264),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_266),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_265),
.A2(n_281),
.B(n_283),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_267),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_267),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_285),
.B2(n_286),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_278),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_278),
.C(n_286),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B(n_277),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_301),
.C(n_305),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g310 ( 
.A(n_277),
.B(n_301),
.CI(n_305),
.CON(n_310),
.SN(n_310)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_281),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_294),
.B(n_297),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_290),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_306),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_306),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_309),
.B(n_310),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_310),
.Y(n_314)
);


endmodule