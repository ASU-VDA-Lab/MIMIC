module fake_ariane_420_n_2619 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_53, n_260, n_362, n_543, n_310, n_236, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_127, n_531, n_2619);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_127;
input n_531;

output n_2619;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_559;
wire n_2233;
wire n_2370;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_696;
wire n_1442;
wire n_798;
wire n_577;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2312;
wire n_670;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_604;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2599;
wire n_727;
wire n_699;
wire n_590;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_2606;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_907;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_596;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_574;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2275;
wire n_2205;
wire n_2183;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_2590;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_573;
wire n_796;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx2_ASAP7_75t_L g558 ( 
.A(n_532),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_180),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_546),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_401),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_523),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_556),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_159),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_481),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_403),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_451),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_195),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_538),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_310),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_72),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_525),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_421),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_284),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_312),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_372),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_166),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_376),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_366),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_128),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_551),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_321),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_490),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_86),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_362),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_25),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_347),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_340),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_487),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_493),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_112),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_550),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_164),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_312),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_259),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_519),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_192),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_334),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_1),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_435),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_234),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_486),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_111),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_132),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_275),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_449),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_303),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_0),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_468),
.Y(n_610)
);

BUFx10_ASAP7_75t_L g611 ( 
.A(n_343),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_58),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_196),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_251),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_74),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_416),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_439),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_354),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_310),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_502),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_555),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_324),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_151),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_552),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_541),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_422),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_93),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_234),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_211),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_537),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_338),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_252),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_554),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_54),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_430),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_303),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_557),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_268),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_41),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_44),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_364),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_549),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_512),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_299),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_5),
.Y(n_645)
);

CKINVDCx16_ASAP7_75t_R g646 ( 
.A(n_2),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_58),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_228),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_41),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_87),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_43),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_437),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_93),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_399),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_264),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_153),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_14),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_228),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_124),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_474),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_443),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_44),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_325),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_291),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_520),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_203),
.Y(n_666)
);

BUFx4f_ASAP7_75t_SL g667 ( 
.A(n_370),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_240),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_527),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_105),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_462),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_193),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_529),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_6),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_475),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_95),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_439),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_543),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_324),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_147),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_198),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_20),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_362),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_438),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_436),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_297),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_7),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_112),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_397),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_230),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_319),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_380),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_13),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_171),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_60),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_495),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_489),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_470),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_542),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_308),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_75),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_245),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_535),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_476),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_249),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_375),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_266),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_340),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_138),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_128),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_424),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_224),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_419),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_355),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_526),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_463),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_167),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_545),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_508),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_4),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_142),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_119),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_36),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_298),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_51),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_271),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_2),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_38),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_135),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_13),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_4),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_429),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_431),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_417),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_540),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_197),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_521),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_548),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_247),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_341),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_114),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_22),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_432),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_287),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_409),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_87),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_323),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_51),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_258),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_233),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_14),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_553),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_79),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_260),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_402),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_395),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_174),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_270),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_390),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_195),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_333),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_132),
.Y(n_762)
);

CKINVDCx14_ASAP7_75t_R g763 ( 
.A(n_343),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_215),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_384),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_471),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_247),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_107),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_501),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_544),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_192),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_3),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_161),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_91),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_273),
.Y(n_775)
);

CKINVDCx20_ASAP7_75t_R g776 ( 
.A(n_547),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_160),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_464),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_331),
.Y(n_779)
);

CKINVDCx16_ASAP7_75t_R g780 ( 
.A(n_503),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_374),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_465),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_539),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_249),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_276),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_378),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_348),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_434),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_511),
.Y(n_789)
);

INVxp33_ASAP7_75t_L g790 ( 
.A(n_759),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_564),
.Y(n_791)
);

BUFx6f_ASAP7_75t_L g792 ( 
.A(n_563),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_564),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_560),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_559),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_559),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_559),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_559),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_647),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_560),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_559),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_763),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_572),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_733),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_780),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_733),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_733),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_558),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_733),
.Y(n_809)
);

CKINVDCx16_ASAP7_75t_R g810 ( 
.A(n_646),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_583),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_647),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_653),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_733),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_602),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_602),
.Y(n_816)
);

INVxp33_ASAP7_75t_SL g817 ( 
.A(n_587),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_561),
.Y(n_818)
);

INVxp33_ASAP7_75t_SL g819 ( 
.A(n_561),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_653),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_578),
.Y(n_821)
);

BUFx8_ASAP7_75t_SL g822 ( 
.A(n_599),
.Y(n_822)
);

INVxp33_ASAP7_75t_L g823 ( 
.A(n_570),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_562),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_717),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_717),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_726),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_679),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_679),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_573),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_577),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_625),
.B(n_1),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_579),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_580),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_589),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_562),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_592),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_578),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_569),
.Y(n_839)
);

CKINVDCx16_ASAP7_75t_R g840 ( 
.A(n_611),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_594),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_778),
.Y(n_842)
);

CKINVDCx14_ASAP7_75t_R g843 ( 
.A(n_673),
.Y(n_843)
);

INVxp33_ASAP7_75t_SL g844 ( 
.A(n_566),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_778),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_726),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_727),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_727),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_734),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_650),
.Y(n_850)
);

CKINVDCx14_ASAP7_75t_R g851 ( 
.A(n_699),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_734),
.Y(n_852)
);

CKINVDCx16_ASAP7_75t_R g853 ( 
.A(n_611),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_757),
.Y(n_854)
);

INVxp33_ASAP7_75t_L g855 ( 
.A(n_598),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_566),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_757),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_784),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_784),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_569),
.Y(n_860)
);

INVxp33_ASAP7_75t_SL g861 ( 
.A(n_568),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_590),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_582),
.Y(n_863)
);

INVxp67_ASAP7_75t_SL g864 ( 
.A(n_605),
.Y(n_864)
);

INVxp67_ASAP7_75t_SL g865 ( 
.A(n_609),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_565),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_590),
.Y(n_867)
);

INVxp33_ASAP7_75t_SL g868 ( 
.A(n_568),
.Y(n_868)
);

CKINVDCx16_ASAP7_75t_R g869 ( 
.A(n_611),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_591),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_614),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_563),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_571),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_615),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_635),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_636),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_591),
.Y(n_877)
);

INVxp33_ASAP7_75t_SL g878 ( 
.A(n_571),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_574),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_621),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_704),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_685),
.Y(n_882)
);

INVxp33_ASAP7_75t_SL g883 ( 
.A(n_574),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_718),
.Y(n_884)
);

CKINVDCx16_ASAP7_75t_R g885 ( 
.A(n_685),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_621),
.Y(n_886)
);

INVxp33_ASAP7_75t_SL g887 ( 
.A(n_575),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_675),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_656),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_563),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_828),
.B(n_685),
.Y(n_891)
);

BUFx8_ASAP7_75t_L g892 ( 
.A(n_828),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_790),
.A2(n_639),
.B1(n_693),
.B2(n_622),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_802),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_792),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_795),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_795),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_794),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_792),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_792),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_792),
.Y(n_901)
);

BUFx12f_ASAP7_75t_L g902 ( 
.A(n_802),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_809),
.Y(n_903)
);

BUFx8_ASAP7_75t_SL g904 ( 
.A(n_822),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_794),
.B(n_650),
.Y(n_905)
);

XNOR2xp5_ASAP7_75t_L g906 ( 
.A(n_811),
.B(n_701),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_796),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_792),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_796),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_843),
.Y(n_910)
);

CKINVDCx6p67_ASAP7_75t_R g911 ( 
.A(n_810),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_872),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_805),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_797),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_800),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_797),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_817),
.A2(n_724),
.B1(n_779),
.B2(n_712),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_872),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_872),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_798),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_872),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_872),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_890),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_890),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_890),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_858),
.B(n_740),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_890),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_823),
.A2(n_576),
.B1(n_581),
.B2(n_575),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_805),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_798),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_890),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_809),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_801),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_862),
.A2(n_675),
.B(n_607),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_801),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_808),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_800),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_824),
.Y(n_938)
);

AOI22x1_ASAP7_75t_SL g939 ( 
.A1(n_803),
.A2(n_581),
.B1(n_585),
.B2(n_576),
.Y(n_939)
);

OA21x2_ASAP7_75t_L g940 ( 
.A1(n_862),
.A2(n_610),
.B(n_593),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_821),
.B(n_689),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_808),
.A2(n_776),
.B1(n_682),
.B2(n_764),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_804),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_818),
.Y(n_944)
);

OAI22x1_ASAP7_75t_SL g945 ( 
.A1(n_881),
.A2(n_586),
.B1(n_588),
.B2(n_585),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_804),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_821),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_806),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_838),
.B(n_661),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_838),
.B(n_789),
.Y(n_950)
);

BUFx12f_ASAP7_75t_L g951 ( 
.A(n_824),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_856),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_806),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_807),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_832),
.A2(n_627),
.B1(n_588),
.B2(n_586),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_936),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_R g957 ( 
.A(n_910),
.B(n_851),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_896),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_938),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_896),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_898),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_897),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_892),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_937),
.B(n_836),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_937),
.B(n_915),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_904),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_938),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_897),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_913),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_907),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_915),
.B(n_898),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_892),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_912),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_907),
.Y(n_974)
);

XNOR2xp5_ASAP7_75t_L g975 ( 
.A(n_917),
.B(n_884),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_954),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_935),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_909),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_951),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_915),
.B(n_836),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_913),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_892),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_951),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_926),
.B(n_793),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_892),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_929),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_906),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_935),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_934),
.A2(n_866),
.B(n_814),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_909),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_898),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_906),
.Y(n_992)
);

CKINVDCx16_ASAP7_75t_R g993 ( 
.A(n_902),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_891),
.B(n_839),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_929),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_891),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_944),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_954),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_947),
.B(n_799),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_935),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_951),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_902),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_914),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_952),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_917),
.Y(n_1005)
);

AND2x6_ASAP7_75t_L g1006 ( 
.A(n_926),
.B(n_563),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_911),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_943),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_916),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_916),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_920),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_940),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_947),
.B(n_812),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_894),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_894),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_943),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_902),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_893),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_905),
.B(n_813),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_920),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_911),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_930),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_930),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_911),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_893),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_942),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_945),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_933),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_947),
.B(n_820),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_943),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_945),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_954),
.Y(n_1032)
);

OA21x2_ASAP7_75t_L g1033 ( 
.A1(n_934),
.A2(n_870),
.B(n_867),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_933),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_946),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_946),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_950),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_950),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_948),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_934),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_942),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_939),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_939),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_948),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1037),
.B(n_839),
.Y(n_1045)
);

AND2x2_ASAP7_75t_SL g1046 ( 
.A(n_993),
.B(n_1018),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_977),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_977),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_988),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_988),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_958),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_1040),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_984),
.B(n_905),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1038),
.B(n_860),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_964),
.B(n_860),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_995),
.B(n_819),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_960),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_986),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_984),
.B(n_863),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_1000),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_994),
.B(n_844),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_999),
.B(n_863),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_980),
.B(n_861),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_976),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1039),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1000),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_973),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1008),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1008),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1044),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_1041),
.A2(n_955),
.B1(n_928),
.B2(n_941),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_1005),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1016),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_999),
.B(n_1013),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1016),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_962),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_968),
.Y(n_1077)
);

NAND3xp33_ASAP7_75t_L g1078 ( 
.A(n_967),
.B(n_955),
.C(n_928),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1030),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_999),
.B(n_868),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_996),
.B(n_878),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1030),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_970),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_974),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1013),
.B(n_905),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_959),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_989),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_961),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_989),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_961),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_956),
.B(n_883),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_978),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1033),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_990),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_997),
.B(n_887),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_973),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_973),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_1013),
.B(n_1029),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1029),
.B(n_840),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1004),
.B(n_853),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_969),
.B(n_879),
.C(n_873),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1029),
.B(n_905),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1041),
.A2(n_941),
.B1(n_940),
.B2(n_949),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1033),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1033),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1014),
.B(n_1015),
.Y(n_1106)
);

OR2x2_ASAP7_75t_L g1107 ( 
.A(n_981),
.B(n_869),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1003),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1009),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1019),
.B(n_941),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1010),
.Y(n_1111)
);

INVx5_ASAP7_75t_L g1112 ( 
.A(n_976),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1011),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_1040),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_976),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_1019),
.B(n_941),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1006),
.B(n_949),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_966),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1020),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1022),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_979),
.B(n_882),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1023),
.A2(n_751),
.B1(n_753),
.B2(n_674),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_979),
.B(n_885),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1028),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1034),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1006),
.B(n_866),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_991),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1001),
.B(n_855),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_991),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_976),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_965),
.B(n_864),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_971),
.B(n_865),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1035),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1036),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_983),
.B(n_874),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1006),
.B(n_842),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_983),
.B(n_582),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1012),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1006),
.B(n_842),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1012),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1012),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_976),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_998),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_998),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1002),
.B(n_667),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_998),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1006),
.B(n_845),
.Y(n_1147)
);

NAND2xp33_ASAP7_75t_L g1148 ( 
.A(n_998),
.B(n_674),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_998),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1006),
.B(n_845),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_966),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1024),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1024),
.Y(n_1153)
);

NOR2x1p5_ASAP7_75t_L g1154 ( 
.A(n_1002),
.B(n_751),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_1007),
.B(n_689),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1032),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1032),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_957),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1017),
.B(n_753),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1032),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_1032),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_SL g1162 ( 
.A(n_1007),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1032),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1017),
.B(n_755),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1026),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1025),
.B(n_755),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1026),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1025),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_1005),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_963),
.B(n_756),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_963),
.B(n_756),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1021),
.Y(n_1172)
);

BUFx8_ASAP7_75t_SL g1173 ( 
.A(n_1021),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_972),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_972),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_975),
.B(n_791),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_982),
.Y(n_1177)
);

NAND2xp33_ASAP7_75t_SL g1178 ( 
.A(n_982),
.B(n_758),
.Y(n_1178)
);

NAND2xp33_ASAP7_75t_L g1179 ( 
.A(n_1042),
.B(n_758),
.Y(n_1179)
);

NAND2xp33_ASAP7_75t_SL g1180 ( 
.A(n_985),
.B(n_765),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1027),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_985),
.B(n_940),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1131),
.B(n_867),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1092),
.Y(n_1184)
);

NOR2xp67_ASAP7_75t_L g1185 ( 
.A(n_1158),
.B(n_1118),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1047),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1058),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1086),
.B(n_975),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1045),
.B(n_584),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_1128),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1092),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1054),
.B(n_584),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1047),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1166),
.B(n_987),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1094),
.Y(n_1195)
);

NAND3xp33_ASAP7_75t_L g1196 ( 
.A(n_1055),
.B(n_831),
.C(n_830),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1048),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1056),
.B(n_1168),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1048),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1095),
.B(n_992),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1094),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_SL g1202 ( 
.A(n_1152),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1074),
.B(n_1108),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1108),
.B(n_940),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1109),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1109),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_1158),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1078),
.A2(n_633),
.B(n_643),
.C(n_630),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1049),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1128),
.B(n_850),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1050),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1176),
.B(n_829),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1110),
.B(n_870),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1091),
.B(n_987),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1135),
.B(n_992),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1100),
.B(n_1081),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1053),
.B(n_877),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1050),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1169),
.B(n_1027),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1059),
.B(n_766),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_R g1221 ( 
.A(n_1118),
.B(n_1031),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1111),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1111),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1053),
.B(n_1116),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1116),
.B(n_877),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1116),
.B(n_880),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_1088),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1113),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1106),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1062),
.B(n_766),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1132),
.B(n_880),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1113),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1098),
.B(n_886),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1120),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1071),
.A2(n_782),
.B1(n_783),
.B2(n_770),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1107),
.B(n_1031),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1120),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1085),
.B(n_886),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1102),
.B(n_888),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1051),
.B(n_888),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_1173),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1107),
.B(n_1042),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1176),
.B(n_833),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1080),
.B(n_1043),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1057),
.B(n_765),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1124),
.B(n_948),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_1169),
.Y(n_1247)
);

NOR2xp67_ASAP7_75t_L g1248 ( 
.A(n_1151),
.B(n_1043),
.Y(n_1248)
);

INVx4_ASAP7_75t_L g1249 ( 
.A(n_1088),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1090),
.B(n_770),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1090),
.B(n_782),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1124),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1152),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1076),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1060),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1077),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_SL g1257 ( 
.A(n_1153),
.B(n_567),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1130),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1083),
.B(n_953),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1161),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1084),
.B(n_953),
.Y(n_1261)
);

INVx5_ASAP7_75t_L g1262 ( 
.A(n_1052),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1161),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1119),
.B(n_903),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1125),
.B(n_903),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1133),
.B(n_903),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_L g1267 ( 
.A(n_1159),
.B(n_767),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1164),
.B(n_767),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1061),
.B(n_768),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1099),
.B(n_1170),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1046),
.B(n_834),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1134),
.B(n_903),
.Y(n_1272)
);

OR2x6_ASAP7_75t_L g1273 ( 
.A(n_1155),
.B(n_1153),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1171),
.B(n_768),
.Y(n_1274)
);

NOR3xp33_ASAP7_75t_L g1275 ( 
.A(n_1145),
.B(n_658),
.C(n_657),
.Y(n_1275)
);

NOR2xp67_ASAP7_75t_L g1276 ( 
.A(n_1151),
.B(n_1101),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1066),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1063),
.B(n_771),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1121),
.B(n_771),
.Y(n_1279)
);

INVx2_ASAP7_75t_SL g1280 ( 
.A(n_1172),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1066),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1065),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1065),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1070),
.B(n_1103),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1123),
.B(n_773),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1070),
.Y(n_1286)
);

A2O1A1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1138),
.A2(n_660),
.B(n_671),
.C(n_669),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1068),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1068),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1173),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1069),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1165),
.B(n_835),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1067),
.B(n_773),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1174),
.B(n_775),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1069),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1064),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1073),
.Y(n_1297)
);

BUFx6f_ASAP7_75t_L g1298 ( 
.A(n_1161),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1174),
.B(n_775),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1127),
.B(n_783),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1073),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1172),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1075),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1127),
.B(n_777),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1129),
.B(n_777),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1161),
.Y(n_1306)
);

BUFx5_ASAP7_75t_L g1307 ( 
.A(n_1138),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1129),
.B(n_781),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1052),
.B(n_781),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1075),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1148),
.B(n_841),
.C(n_837),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1067),
.B(n_786),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1067),
.B(n_786),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1079),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1096),
.B(n_659),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1096),
.B(n_664),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1082),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1096),
.B(n_677),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1161),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1130),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1046),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1126),
.Y(n_1322)
);

INVxp33_ASAP7_75t_L g1323 ( 
.A(n_1165),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1175),
.B(n_1177),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1097),
.B(n_680),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1072),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1182),
.A2(n_762),
.B1(n_740),
.B2(n_694),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_1167),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1097),
.B(n_684),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1052),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1146),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1175),
.B(n_595),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1146),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1167),
.B(n_871),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1052),
.B(n_1114),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1087),
.A2(n_715),
.B(n_698),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1130),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1156),
.Y(n_1338)
);

NOR3xp33_ASAP7_75t_L g1339 ( 
.A(n_1137),
.B(n_1180),
.C(n_1178),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1140),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_SL g1341 ( 
.A(n_1052),
.B(n_567),
.Y(n_1341)
);

AND2x6_ASAP7_75t_L g1342 ( 
.A(n_1114),
.B(n_752),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1140),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1114),
.B(n_596),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1141),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1097),
.B(n_709),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1154),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1157),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1177),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1155),
.B(n_600),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1064),
.B(n_601),
.Y(n_1351)
);

INVxp67_ASAP7_75t_L g1352 ( 
.A(n_1178),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1157),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1141),
.B(n_1093),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1155),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1093),
.B(n_932),
.Y(n_1356)
);

BUFx5_ASAP7_75t_L g1357 ( 
.A(n_1142),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1104),
.B(n_932),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1136),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1142),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_SL g1361 ( 
.A(n_1155),
.Y(n_1361)
);

AND2x2_ASAP7_75t_SL g1362 ( 
.A(n_1179),
.B(n_1181),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1143),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1104),
.B(n_932),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1139),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1105),
.B(n_1117),
.Y(n_1366)
);

INVxp33_ASAP7_75t_L g1367 ( 
.A(n_1122),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1162),
.B(n_604),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1162),
.B(n_606),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1064),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1105),
.B(n_769),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1143),
.B(n_912),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1147),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1162),
.B(n_608),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1064),
.B(n_612),
.Y(n_1375)
);

BUFx5_ASAP7_75t_L g1376 ( 
.A(n_1144),
.Y(n_1376)
);

AND2x4_ASAP7_75t_SL g1377 ( 
.A(n_1072),
.B(n_740),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1064),
.B(n_613),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1144),
.B(n_912),
.Y(n_1379)
);

OR2x2_ASAP7_75t_SL g1380 ( 
.A(n_1290),
.B(n_1219),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1184),
.Y(n_1381)
);

AO22x2_ASAP7_75t_L g1382 ( 
.A1(n_1321),
.A2(n_1181),
.B1(n_1180),
.B2(n_1179),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1221),
.Y(n_1383)
);

NAND2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1227),
.B(n_1181),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1224),
.B(n_1112),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1191),
.Y(n_1386)
);

OAI221xp5_ASAP7_75t_L g1387 ( 
.A1(n_1274),
.A2(n_1148),
.B1(n_889),
.B2(n_876),
.C(n_875),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1216),
.B(n_762),
.Y(n_1388)
);

AO22x2_ASAP7_75t_L g1389 ( 
.A1(n_1271),
.A2(n_1150),
.B1(n_1160),
.B2(n_816),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1186),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1267),
.A2(n_1160),
.B1(n_1163),
.B2(n_1149),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1268),
.A2(n_1149),
.B1(n_1115),
.B2(n_617),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1195),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1201),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1254),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1256),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1205),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1193),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1206),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1222),
.Y(n_1400)
);

CKINVDCx20_ASAP7_75t_R g1401 ( 
.A(n_1241),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1187),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1273),
.B(n_1115),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1198),
.B(n_1243),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1197),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1269),
.A2(n_1149),
.B1(n_1115),
.B2(n_618),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_1377),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1223),
.Y(n_1408)
);

AO22x2_ASAP7_75t_L g1409 ( 
.A1(n_1284),
.A2(n_816),
.B1(n_825),
.B2(n_815),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1326),
.Y(n_1410)
);

AOI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1194),
.A2(n_619),
.B1(n_623),
.B2(n_616),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1188),
.B(n_762),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1215),
.B(n_1112),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1247),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1212),
.B(n_1112),
.Y(n_1415)
);

AO22x2_ASAP7_75t_L g1416 ( 
.A1(n_1284),
.A2(n_825),
.B1(n_826),
.B2(n_815),
.Y(n_1416)
);

BUFx8_ASAP7_75t_L g1417 ( 
.A(n_1361),
.Y(n_1417)
);

NAND2x1p5_ASAP7_75t_L g1418 ( 
.A(n_1227),
.B(n_1112),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1334),
.B(n_1112),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1190),
.Y(n_1420)
);

OAI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1200),
.A2(n_1214),
.B1(n_1350),
.B2(n_1235),
.C(n_1270),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1257),
.B(n_626),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1228),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1210),
.B(n_826),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1232),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1326),
.B(n_827),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1199),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1292),
.B(n_827),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1367),
.B(n_628),
.Y(n_1429)
);

BUFx8_ASAP7_75t_L g1430 ( 
.A(n_1361),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1242),
.A2(n_629),
.B1(n_632),
.B2(n_631),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1234),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1237),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1252),
.Y(n_1434)
);

AO22x2_ASAP7_75t_L g1435 ( 
.A1(n_1339),
.A2(n_847),
.B1(n_848),
.B2(n_846),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1253),
.Y(n_1436)
);

OAI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1278),
.A2(n_728),
.B1(n_741),
.B2(n_721),
.C(n_711),
.Y(n_1437)
);

OAI221xp5_ASAP7_75t_L g1438 ( 
.A1(n_1275),
.A2(n_761),
.B1(n_772),
.B2(n_760),
.C(n_754),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1207),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1282),
.Y(n_1440)
);

NAND2xp33_ASAP7_75t_L g1441 ( 
.A(n_1307),
.B(n_1357),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1203),
.B(n_634),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1203),
.B(n_638),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1183),
.B(n_640),
.Y(n_1444)
);

AO22x2_ASAP7_75t_L g1445 ( 
.A1(n_1355),
.A2(n_847),
.B1(n_848),
.B2(n_846),
.Y(n_1445)
);

OAI221xp5_ASAP7_75t_L g1446 ( 
.A1(n_1279),
.A2(n_787),
.B1(n_788),
.B2(n_785),
.C(n_774),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1283),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1328),
.B(n_641),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1324),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1286),
.Y(n_1450)
);

AO22x2_ASAP7_75t_L g1451 ( 
.A1(n_1349),
.A2(n_849),
.B1(n_854),
.B2(n_852),
.Y(n_1451)
);

BUFx8_ASAP7_75t_L g1452 ( 
.A(n_1202),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1236),
.B(n_849),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1273),
.B(n_852),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1352),
.B(n_644),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1233),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1264),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1217),
.B(n_645),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1264),
.Y(n_1459)
);

OAI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1285),
.A2(n_652),
.B1(n_654),
.B2(n_651),
.C(n_648),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1229),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1257),
.B(n_649),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1265),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1265),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1362),
.B(n_655),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1209),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1208),
.A2(n_1311),
.B(n_1196),
.C(n_1287),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1276),
.A2(n_1244),
.B1(n_1185),
.B2(n_1273),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1207),
.B(n_662),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1249),
.B(n_1262),
.Y(n_1470)
);

OAI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1294),
.A2(n_666),
.B1(n_670),
.B2(n_668),
.C(n_663),
.Y(n_1471)
);

AO22x2_ASAP7_75t_L g1472 ( 
.A1(n_1280),
.A2(n_854),
.B1(n_859),
.B2(n_857),
.Y(n_1472)
);

AO22x2_ASAP7_75t_L g1473 ( 
.A1(n_1302),
.A2(n_857),
.B1(n_859),
.B2(n_1087),
.Y(n_1473)
);

NAND2x1p5_ASAP7_75t_L g1474 ( 
.A(n_1249),
.B(n_1262),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1225),
.B(n_672),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1347),
.B(n_1089),
.Y(n_1476)
);

NAND2xp33_ASAP7_75t_L g1477 ( 
.A(n_1307),
.B(n_1089),
.Y(n_1477)
);

NAND2x1p5_ASAP7_75t_L g1478 ( 
.A(n_1262),
.B(n_954),
.Y(n_1478)
);

AO22x2_ASAP7_75t_L g1479 ( 
.A1(n_1311),
.A2(n_624),
.B1(n_814),
.B2(n_807),
.Y(n_1479)
);

AO22x2_ASAP7_75t_L g1480 ( 
.A1(n_1196),
.A2(n_624),
.B1(n_912),
.B2(n_5),
.Y(n_1480)
);

OAI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1299),
.A2(n_683),
.B1(n_687),
.B2(n_686),
.C(n_676),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1266),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1266),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1272),
.Y(n_1484)
);

BUFx8_ASAP7_75t_L g1485 ( 
.A(n_1202),
.Y(n_1485)
);

AO22x2_ASAP7_75t_L g1486 ( 
.A1(n_1340),
.A2(n_6),
.B1(n_0),
.B2(n_3),
.Y(n_1486)
);

NAND2x1p5_ASAP7_75t_L g1487 ( 
.A(n_1296),
.B(n_954),
.Y(n_1487)
);

AO22x2_ASAP7_75t_L g1488 ( 
.A1(n_1343),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_1488)
);

AO22x2_ASAP7_75t_L g1489 ( 
.A1(n_1345),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1332),
.B(n_1368),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1272),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1240),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1369),
.B(n_681),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1374),
.B(n_688),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1245),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1226),
.B(n_690),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1211),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1259),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1231),
.B(n_691),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1248),
.A2(n_695),
.B1(n_700),
.B2(n_692),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1296),
.B(n_954),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1218),
.Y(n_1502)
);

AO22x2_ASAP7_75t_L g1503 ( 
.A1(n_1366),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1213),
.B(n_1323),
.Y(n_1504)
);

OAI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1220),
.A2(n_706),
.B1(n_707),
.B2(n_705),
.C(n_702),
.Y(n_1505)
);

AO22x2_ASAP7_75t_L g1506 ( 
.A1(n_1366),
.A2(n_15),
.B1(n_11),
.B2(n_12),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1255),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1260),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1259),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1261),
.Y(n_1510)
);

OAI221xp5_ASAP7_75t_L g1511 ( 
.A1(n_1230),
.A2(n_713),
.B1(n_714),
.B2(n_710),
.C(n_708),
.Y(n_1511)
);

AO22x2_ASAP7_75t_L g1512 ( 
.A1(n_1288),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1261),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1238),
.B(n_720),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1289),
.Y(n_1515)
);

NAND2x1p5_ASAP7_75t_L g1516 ( 
.A(n_1370),
.B(n_901),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1304),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1291),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1297),
.Y(n_1519)
);

NAND2x1p5_ASAP7_75t_L g1520 ( 
.A(n_1370),
.B(n_901),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1258),
.B(n_901),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1189),
.A2(n_723),
.B1(n_725),
.B2(n_722),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1192),
.A2(n_730),
.B1(n_731),
.B2(n_729),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1301),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1239),
.B(n_750),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1303),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1258),
.B(n_1320),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1305),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1315),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1260),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1308),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1354),
.A2(n_736),
.B1(n_739),
.B2(n_732),
.Y(n_1532)
);

OA22x2_ASAP7_75t_L g1533 ( 
.A1(n_1250),
.A2(n_743),
.B1(n_744),
.B2(n_742),
.Y(n_1533)
);

AO22x2_ASAP7_75t_L g1534 ( 
.A1(n_1354),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1534)
);

AO22x2_ASAP7_75t_L g1535 ( 
.A1(n_1277),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1251),
.B(n_745),
.Y(n_1536)
);

AO22x2_ASAP7_75t_L g1537 ( 
.A1(n_1281),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1327),
.B(n_746),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1260),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1316),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1309),
.B(n_563),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1318),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1293),
.B(n_1312),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1325),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1329),
.Y(n_1545)
);

NAND3xp33_ASAP7_75t_SL g1546 ( 
.A(n_1313),
.B(n_748),
.C(n_747),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1346),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1295),
.Y(n_1548)
);

AO22x2_ASAP7_75t_L g1549 ( 
.A1(n_1310),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1314),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1360),
.B(n_749),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1363),
.B(n_23),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1317),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1246),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1300),
.B(n_597),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1320),
.B(n_918),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1246),
.Y(n_1557)
);

AO22x2_ASAP7_75t_L g1558 ( 
.A1(n_1322),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1558)
);

AO22x2_ASAP7_75t_L g1559 ( 
.A1(n_1371),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1331),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1333),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1338),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1330),
.B(n_637),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1263),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1263),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1348),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1353),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1344),
.B(n_603),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_L g1569 ( 
.A(n_1341),
.B(n_620),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1371),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1204),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1341),
.A2(n_642),
.B1(n_678),
.B2(n_665),
.Y(n_1572)
);

AO22x2_ASAP7_75t_L g1573 ( 
.A1(n_1359),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1204),
.Y(n_1574)
);

OAI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1351),
.A2(n_697),
.B1(n_716),
.B2(n_703),
.C(n_696),
.Y(n_1575)
);

OAI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1375),
.A2(n_735),
.B1(n_738),
.B2(n_737),
.C(n_719),
.Y(n_1576)
);

AO22x2_ASAP7_75t_L g1577 ( 
.A1(n_1365),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1336),
.B(n_30),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1372),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1373),
.A2(n_752),
.B1(n_637),
.B2(n_918),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1357),
.A2(n_752),
.B1(n_637),
.B2(n_918),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1404),
.B(n_1357),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1421),
.A2(n_1337),
.B1(n_1330),
.B2(n_1378),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1449),
.B(n_1357),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1402),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1388),
.B(n_31),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1477),
.A2(n_1335),
.B(n_1298),
.Y(n_1587)
);

INVx3_ASAP7_75t_L g1588 ( 
.A(n_1564),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1490),
.B(n_1357),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1424),
.B(n_1376),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1453),
.B(n_32),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1412),
.B(n_1376),
.Y(n_1592)
);

INVx4_ASAP7_75t_L g1593 ( 
.A(n_1383),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1441),
.A2(n_1298),
.B(n_1263),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1543),
.A2(n_1306),
.B(n_1298),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1429),
.A2(n_1413),
.B1(n_1494),
.B2(n_1407),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1460),
.A2(n_1379),
.B(n_1337),
.C(n_1358),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1492),
.B(n_1376),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_R g1599 ( 
.A(n_1401),
.B(n_1306),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1471),
.A2(n_1379),
.B(n_1358),
.C(n_1364),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1498),
.A2(n_1319),
.B(n_1306),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1390),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1509),
.A2(n_1319),
.B(n_1330),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1510),
.A2(n_1319),
.B(n_1356),
.Y(n_1604)
);

OR2x6_ASAP7_75t_L g1605 ( 
.A(n_1403),
.B(n_1356),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1398),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1467),
.A2(n_1342),
.B(n_1364),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1495),
.A2(n_1307),
.B1(n_1336),
.B2(n_1376),
.Y(n_1608)
);

BUFx4f_ASAP7_75t_L g1609 ( 
.A(n_1403),
.Y(n_1609)
);

AO22x1_ASAP7_75t_L g1610 ( 
.A1(n_1417),
.A2(n_1430),
.B1(n_1485),
.B2(n_1452),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1513),
.A2(n_1307),
.B(n_1376),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1405),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1406),
.A2(n_1307),
.B1(n_1342),
.B2(n_752),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1414),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1426),
.B(n_32),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1428),
.B(n_1342),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1395),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1504),
.B(n_1342),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1508),
.B(n_919),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1410),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1530),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1414),
.B(n_33),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1420),
.B(n_33),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1396),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1461),
.B(n_34),
.Y(n_1625)
);

BUFx8_ASAP7_75t_SL g1626 ( 
.A(n_1436),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1385),
.B(n_922),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1569),
.A2(n_752),
.B1(n_637),
.B2(n_925),
.Y(n_1628)
);

BUFx4f_ASAP7_75t_L g1629 ( 
.A(n_1436),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1529),
.B(n_34),
.Y(n_1630)
);

AOI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1473),
.A2(n_925),
.B(n_899),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1385),
.B(n_1527),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1444),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1540),
.B(n_35),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1427),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1481),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1422),
.B(n_39),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1570),
.A2(n_899),
.B(n_895),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1462),
.B(n_40),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_1417),
.Y(n_1640)
);

O2A1O1Ixp5_ASAP7_75t_L g1641 ( 
.A1(n_1465),
.A2(n_43),
.B(n_40),
.C(n_42),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1571),
.A2(n_899),
.B(n_895),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1542),
.B(n_42),
.Y(n_1643)
);

AOI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1574),
.A2(n_931),
.B(n_899),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1544),
.B(n_45),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1454),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1457),
.A2(n_924),
.B(n_899),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1439),
.Y(n_1648)
);

NAND3xp33_ASAP7_75t_L g1649 ( 
.A(n_1431),
.B(n_899),
.C(n_895),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1459),
.A2(n_900),
.B(n_895),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1463),
.A2(n_900),
.B(n_895),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1455),
.B(n_45),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1381),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1545),
.A2(n_1547),
.B(n_1536),
.C(n_1555),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1456),
.B(n_46),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1527),
.B(n_1419),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1493),
.B(n_46),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1464),
.A2(n_900),
.B(n_895),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1482),
.A2(n_931),
.B(n_908),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1486),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1483),
.A2(n_924),
.B(n_908),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1484),
.A2(n_931),
.B(n_908),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1546),
.B(n_47),
.C(n_48),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1415),
.B(n_900),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1386),
.B(n_49),
.Y(n_1665)
);

AOI22x1_ASAP7_75t_L g1666 ( 
.A1(n_1480),
.A2(n_908),
.B1(n_921),
.B2(n_900),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1564),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1393),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1491),
.A2(n_908),
.B(n_900),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1394),
.B(n_50),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1539),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1469),
.A2(n_931),
.B1(n_921),
.B2(n_923),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1551),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1448),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1440),
.B(n_50),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1476),
.B(n_440),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1554),
.A2(n_931),
.B(n_921),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1447),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1450),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_SL g1680 ( 
.A1(n_1552),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1391),
.A2(n_924),
.B(n_921),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1468),
.B(n_908),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1466),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1499),
.B(n_52),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1497),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1392),
.B(n_921),
.Y(n_1686)
);

A2O1A1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1568),
.A2(n_923),
.B(n_927),
.C(n_921),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1442),
.B(n_53),
.Y(n_1688)
);

AO21x1_ASAP7_75t_L g1689 ( 
.A1(n_1578),
.A2(n_55),
.B(n_56),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1397),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1443),
.B(n_55),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1476),
.B(n_441),
.Y(n_1692)
);

OAI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1557),
.A2(n_924),
.B(n_923),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1579),
.A2(n_924),
.B(n_923),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1502),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1539),
.B(n_923),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1563),
.A2(n_927),
.B(n_923),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1563),
.A2(n_931),
.B(n_927),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1507),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1384),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1387),
.A2(n_59),
.B(n_56),
.C(n_57),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1458),
.B(n_57),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1411),
.B(n_1382),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1565),
.B(n_927),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1446),
.A2(n_927),
.B(n_924),
.C(n_61),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1501),
.A2(n_927),
.B(n_924),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1501),
.A2(n_444),
.B(n_442),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1382),
.B(n_59),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1514),
.A2(n_446),
.B(n_445),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1517),
.B(n_60),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1525),
.B(n_61),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1475),
.B(n_62),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1521),
.A2(n_448),
.B(n_447),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1521),
.A2(n_452),
.B(n_450),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1496),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1715)
);

AND2x2_ASAP7_75t_SL g1716 ( 
.A(n_1535),
.B(n_63),
.Y(n_1716)
);

AOI33xp33_ASAP7_75t_L g1717 ( 
.A1(n_1522),
.A2(n_66),
.A3(n_68),
.B1(n_64),
.B2(n_65),
.B3(n_67),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1418),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1399),
.B(n_65),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1400),
.B(n_66),
.Y(n_1720)
);

A2O1A1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1437),
.A2(n_1438),
.B(n_1538),
.C(n_1531),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1528),
.B(n_67),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1556),
.A2(n_454),
.B(n_453),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1408),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1423),
.B(n_68),
.Y(n_1725)
);

NAND2xp33_ASAP7_75t_L g1726 ( 
.A(n_1470),
.B(n_69),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1425),
.B(n_69),
.Y(n_1727)
);

O2A1O1Ixp5_ASAP7_75t_L g1728 ( 
.A1(n_1532),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1486),
.A2(n_73),
.B1(n_70),
.B2(n_71),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1432),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1572),
.B(n_1556),
.Y(n_1731)
);

BUFx12f_ASAP7_75t_L g1732 ( 
.A(n_1380),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1433),
.B(n_73),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1505),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1500),
.B(n_76),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1434),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1435),
.A2(n_456),
.B(n_455),
.Y(n_1737)
);

OA22x2_ASAP7_75t_L g1738 ( 
.A1(n_1541),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1511),
.B(n_77),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1488),
.B(n_78),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1435),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1451),
.B(n_80),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1581),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1451),
.B(n_81),
.Y(n_1744)
);

BUFx4f_ASAP7_75t_L g1745 ( 
.A(n_1474),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1515),
.A2(n_1519),
.B(n_1518),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1488),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1524),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1526),
.B(n_83),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1480),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1548),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1487),
.A2(n_85),
.B(n_88),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1550),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1473),
.A2(n_1520),
.B(n_1516),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1533),
.B(n_88),
.Y(n_1755)
);

A2O1A1Ixp33_ASAP7_75t_L g1756 ( 
.A1(n_1523),
.A2(n_91),
.B(n_89),
.C(n_90),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1472),
.B(n_89),
.Y(n_1757)
);

NOR3xp33_ASAP7_75t_L g1758 ( 
.A(n_1575),
.B(n_90),
.C(n_92),
.Y(n_1758)
);

AOI21xp33_ASAP7_75t_L g1759 ( 
.A1(n_1389),
.A2(n_92),
.B(n_94),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1561),
.B(n_94),
.Y(n_1760)
);

OAI321xp33_ASAP7_75t_L g1761 ( 
.A1(n_1541),
.A2(n_97),
.A3(n_99),
.B1(n_95),
.B2(n_96),
.C(n_98),
.Y(n_1761)
);

O2A1O1Ixp33_ASAP7_75t_L g1762 ( 
.A1(n_1576),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_1762)
);

CKINVDCx20_ASAP7_75t_R g1763 ( 
.A(n_1560),
.Y(n_1763)
);

NAND2xp33_ASAP7_75t_R g1764 ( 
.A(n_1562),
.B(n_457),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1478),
.A2(n_459),
.B(n_458),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1566),
.B(n_99),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1534),
.A2(n_461),
.B(n_460),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1553),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1567),
.B(n_100),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1489),
.A2(n_1573),
.B1(n_1577),
.B2(n_1558),
.Y(n_1770)
);

INVx5_ASAP7_75t_L g1771 ( 
.A(n_1472),
.Y(n_1771)
);

AO22x1_ASAP7_75t_L g1772 ( 
.A1(n_1740),
.A2(n_1489),
.B1(n_1512),
.B2(n_1558),
.Y(n_1772)
);

BUFx12f_ASAP7_75t_L g1773 ( 
.A(n_1640),
.Y(n_1773)
);

INVx5_ASAP7_75t_L g1774 ( 
.A(n_1626),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1591),
.B(n_1573),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1751),
.Y(n_1776)
);

BUFx4f_ASAP7_75t_L g1777 ( 
.A(n_1732),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_R g1778 ( 
.A(n_1629),
.B(n_466),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1614),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1611),
.A2(n_1559),
.B(n_1534),
.Y(n_1780)
);

O2A1O1Ixp33_ASAP7_75t_SL g1781 ( 
.A1(n_1652),
.A2(n_1512),
.B(n_1506),
.C(n_1503),
.Y(n_1781)
);

A2O1A1Ixp33_ASAP7_75t_L g1782 ( 
.A1(n_1770),
.A2(n_1577),
.B(n_1537),
.C(n_1549),
.Y(n_1782)
);

AOI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1660),
.A2(n_1559),
.B1(n_1506),
.B2(n_1503),
.C(n_1537),
.Y(n_1783)
);

AO21x1_ASAP7_75t_L g1784 ( 
.A1(n_1660),
.A2(n_1549),
.B(n_1535),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1615),
.B(n_1445),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1609),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1617),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1629),
.Y(n_1788)
);

OAI22xp5_ASAP7_75t_L g1789 ( 
.A1(n_1735),
.A2(n_1445),
.B1(n_1389),
.B2(n_1479),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1596),
.B(n_1580),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1610),
.Y(n_1791)
);

NAND3xp33_ASAP7_75t_SL g1792 ( 
.A(n_1750),
.B(n_100),
.C(n_101),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1594),
.A2(n_1416),
.B(n_1409),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1593),
.B(n_101),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1620),
.B(n_1409),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1620),
.B(n_1416),
.Y(n_1796)
);

A2O1A1Ixp33_ASAP7_75t_L g1797 ( 
.A1(n_1654),
.A2(n_1479),
.B(n_104),
.C(n_102),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1585),
.B(n_102),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1592),
.B(n_103),
.Y(n_1799)
);

INVxp67_ASAP7_75t_L g1800 ( 
.A(n_1671),
.Y(n_1800)
);

OR2x6_ASAP7_75t_L g1801 ( 
.A(n_1621),
.B(n_1676),
.Y(n_1801)
);

A2O1A1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1701),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1589),
.B(n_106),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1673),
.B(n_106),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_L g1805 ( 
.A(n_1609),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1646),
.B(n_1674),
.Y(n_1806)
);

A2O1A1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1739),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_SL g1808 ( 
.A1(n_1729),
.A2(n_108),
.B(n_109),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1586),
.B(n_110),
.Y(n_1809)
);

HB1xp67_ASAP7_75t_L g1810 ( 
.A(n_1590),
.Y(n_1810)
);

NAND2xp33_ASAP7_75t_R g1811 ( 
.A(n_1599),
.B(n_467),
.Y(n_1811)
);

A2O1A1Ixp33_ASAP7_75t_L g1812 ( 
.A1(n_1636),
.A2(n_113),
.B(n_110),
.C(n_111),
.Y(n_1812)
);

BUFx2_ASAP7_75t_L g1813 ( 
.A(n_1588),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1624),
.B(n_113),
.Y(n_1814)
);

O2A1O1Ixp33_ASAP7_75t_SL g1815 ( 
.A1(n_1756),
.A2(n_1734),
.B(n_1747),
.C(n_1729),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1607),
.A2(n_114),
.B(n_115),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1676),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1763),
.Y(n_1818)
);

NAND2x1p5_ASAP7_75t_L g1819 ( 
.A(n_1745),
.B(n_469),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1653),
.B(n_115),
.Y(n_1820)
);

O2A1O1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1721),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1668),
.B(n_116),
.Y(n_1822)
);

AND2x6_ASAP7_75t_L g1823 ( 
.A(n_1708),
.B(n_1692),
.Y(n_1823)
);

OAI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1738),
.A2(n_1747),
.B1(n_1761),
.B2(n_1771),
.Y(n_1824)
);

BUFx4f_ASAP7_75t_L g1825 ( 
.A(n_1692),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1678),
.B(n_117),
.Y(n_1826)
);

O2A1O1Ixp5_ASAP7_75t_L g1827 ( 
.A1(n_1767),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_1827)
);

NOR3xp33_ASAP7_75t_L g1828 ( 
.A(n_1761),
.B(n_120),
.C(n_121),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1679),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1607),
.A2(n_121),
.B(n_122),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1690),
.B(n_1724),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1730),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1588),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1587),
.A2(n_122),
.B(n_123),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1736),
.B(n_123),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1593),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1748),
.B(n_124),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1716),
.B(n_125),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1764),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1630),
.B(n_125),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1768),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1705),
.A2(n_126),
.B(n_127),
.Y(n_1842)
);

NAND2x1p5_ASAP7_75t_L g1843 ( 
.A(n_1745),
.B(n_1667),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1648),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1753),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1681),
.A2(n_1582),
.B(n_1598),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1681),
.A2(n_126),
.B(n_127),
.Y(n_1847)
);

AO32x1_ASAP7_75t_L g1848 ( 
.A1(n_1608),
.A2(n_131),
.A3(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1622),
.B(n_129),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1657),
.B(n_130),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1613),
.A2(n_131),
.B(n_133),
.Y(n_1851)
);

OAI21x1_ASAP7_75t_L g1852 ( 
.A1(n_1642),
.A2(n_473),
.B(n_472),
.Y(n_1852)
);

A2O1A1Ixp33_ASAP7_75t_L g1853 ( 
.A1(n_1762),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1602),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1634),
.B(n_134),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1647),
.A2(n_136),
.B(n_137),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1667),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1643),
.B(n_137),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1710),
.B(n_138),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1583),
.B(n_139),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1606),
.Y(n_1861)
);

CKINVDCx20_ASAP7_75t_R g1862 ( 
.A(n_1623),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1647),
.A2(n_139),
.B(n_140),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1718),
.Y(n_1864)
);

AND2x4_ASAP7_75t_SL g1865 ( 
.A(n_1605),
.B(n_1718),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1645),
.B(n_140),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1584),
.Y(n_1867)
);

BUFx6f_ASAP7_75t_L g1868 ( 
.A(n_1605),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1625),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1655),
.B(n_141),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1722),
.B(n_1637),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1661),
.A2(n_141),
.B(n_142),
.Y(n_1872)
);

O2A1O1Ixp5_ASAP7_75t_SL g1873 ( 
.A1(n_1759),
.A2(n_145),
.B(n_143),
.C(n_144),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1612),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1635),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1661),
.A2(n_143),
.B(n_144),
.Y(n_1876)
);

NAND2x1_ASAP7_75t_L g1877 ( 
.A(n_1583),
.B(n_477),
.Y(n_1877)
);

O2A1O1Ixp33_ASAP7_75t_SL g1878 ( 
.A1(n_1684),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_1878)
);

OAI21xp33_ASAP7_75t_SL g1879 ( 
.A1(n_1738),
.A2(n_146),
.B(n_148),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1683),
.Y(n_1880)
);

A2O1A1Ixp33_ASAP7_75t_L g1881 ( 
.A1(n_1688),
.A2(n_150),
.B(n_148),
.C(n_149),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1685),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1639),
.B(n_149),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_SL g1884 ( 
.A1(n_1771),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_1884)
);

O2A1O1Ixp33_ASAP7_75t_SL g1885 ( 
.A1(n_1743),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_1885)
);

NAND2xp33_ASAP7_75t_SL g1886 ( 
.A(n_1717),
.B(n_154),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1605),
.Y(n_1887)
);

O2A1O1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1758),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_1888)
);

NOR3xp33_ASAP7_75t_SL g1889 ( 
.A(n_1633),
.B(n_155),
.C(n_156),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1632),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1691),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1693),
.A2(n_158),
.B(n_160),
.Y(n_1892)
);

NOR2xp67_ASAP7_75t_L g1893 ( 
.A(n_1700),
.B(n_478),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1749),
.B(n_161),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1695),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1766),
.B(n_162),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_L g1897 ( 
.A1(n_1711),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_1897)
);

NOR3xp33_ASAP7_75t_L g1898 ( 
.A(n_1715),
.B(n_1663),
.C(n_1755),
.Y(n_1898)
);

INVxp67_ASAP7_75t_L g1899 ( 
.A(n_1712),
.Y(n_1899)
);

INVx2_ASAP7_75t_SL g1900 ( 
.A(n_1699),
.Y(n_1900)
);

O2A1O1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1702),
.A2(n_166),
.B(n_163),
.C(n_165),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_SL g1902 ( 
.A(n_1616),
.B(n_165),
.Y(n_1902)
);

O2A1O1Ixp33_ASAP7_75t_L g1903 ( 
.A1(n_1680),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_1903)
);

O2A1O1Ixp33_ASAP7_75t_L g1904 ( 
.A1(n_1726),
.A2(n_1744),
.B(n_1757),
.C(n_1742),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1771),
.B(n_168),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1746),
.B(n_169),
.Y(n_1906)
);

INVx8_ASAP7_75t_L g1907 ( 
.A(n_1771),
.Y(n_1907)
);

OAI21x1_ASAP7_75t_L g1908 ( 
.A1(n_1644),
.A2(n_480),
.B(n_479),
.Y(n_1908)
);

CKINVDCx6p67_ASAP7_75t_R g1909 ( 
.A(n_1665),
.Y(n_1909)
);

AOI21xp33_ASAP7_75t_L g1910 ( 
.A1(n_1703),
.A2(n_170),
.B(n_171),
.Y(n_1910)
);

A2O1A1Ixp33_ASAP7_75t_SL g1911 ( 
.A1(n_1752),
.A2(n_173),
.B(n_170),
.C(n_172),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1693),
.A2(n_172),
.B(n_173),
.Y(n_1912)
);

A2O1A1Ixp33_ASAP7_75t_L g1913 ( 
.A1(n_1737),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1746),
.Y(n_1914)
);

O2A1O1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1752),
.A2(n_177),
.B(n_175),
.C(n_176),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1769),
.B(n_177),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1670),
.B(n_178),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1675),
.Y(n_1918)
);

INVx5_ASAP7_75t_L g1919 ( 
.A(n_1666),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1741),
.B(n_178),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1597),
.A2(n_179),
.B(n_180),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1656),
.B(n_179),
.Y(n_1922)
);

OR2x6_ASAP7_75t_L g1923 ( 
.A(n_1731),
.B(n_482),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1719),
.B(n_181),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1720),
.B(n_181),
.Y(n_1925)
);

INVxp67_ASAP7_75t_L g1926 ( 
.A(n_1725),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1727),
.B(n_182),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_SL g1928 ( 
.A1(n_1649),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_1928)
);

O2A1O1Ixp5_ASAP7_75t_SL g1929 ( 
.A1(n_1682),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1733),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1618),
.B(n_185),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1754),
.B(n_186),
.Y(n_1932)
);

INVx6_ASAP7_75t_L g1933 ( 
.A(n_1619),
.Y(n_1933)
);

NOR2x1_ASAP7_75t_L g1934 ( 
.A(n_1595),
.B(n_186),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1689),
.Y(n_1935)
);

OAI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1672),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_1936)
);

OA22x2_ASAP7_75t_L g1937 ( 
.A1(n_1760),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1696),
.B(n_190),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1600),
.B(n_190),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1603),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1694),
.Y(n_1941)
);

BUFx6f_ASAP7_75t_L g1942 ( 
.A(n_1619),
.Y(n_1942)
);

OAI21x1_ASAP7_75t_L g1943 ( 
.A1(n_1793),
.A2(n_1631),
.B(n_1650),
.Y(n_1943)
);

AO22x2_ASAP7_75t_L g1944 ( 
.A1(n_1789),
.A2(n_1601),
.B1(n_1604),
.B2(n_1627),
.Y(n_1944)
);

OAI21xp5_ASAP7_75t_L g1945 ( 
.A1(n_1871),
.A2(n_1728),
.B(n_1641),
.Y(n_1945)
);

AND2x6_ASAP7_75t_L g1946 ( 
.A(n_1817),
.B(n_1628),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1779),
.Y(n_1947)
);

INVxp67_ASAP7_75t_L g1948 ( 
.A(n_1806),
.Y(n_1948)
);

OAI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1859),
.A2(n_1709),
.B1(n_1686),
.B2(n_1713),
.Y(n_1949)
);

AO21x2_ASAP7_75t_L g1950 ( 
.A1(n_1780),
.A2(n_1638),
.B(n_1677),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1787),
.Y(n_1951)
);

OA21x2_ASAP7_75t_L g1952 ( 
.A1(n_1935),
.A2(n_1687),
.B(n_1658),
.Y(n_1952)
);

INVx3_ASAP7_75t_L g1953 ( 
.A(n_1868),
.Y(n_1953)
);

O2A1O1Ixp5_ASAP7_75t_L g1954 ( 
.A1(n_1816),
.A2(n_1830),
.B(n_1860),
.C(n_1824),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1829),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1832),
.Y(n_1956)
);

AOI221x1_ASAP7_75t_L g1957 ( 
.A1(n_1828),
.A2(n_1662),
.B1(n_1669),
.B2(n_1659),
.C(n_1651),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1801),
.B(n_1868),
.Y(n_1958)
);

AOI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1919),
.A2(n_1694),
.B(n_1664),
.Y(n_1959)
);

O2A1O1Ixp5_ASAP7_75t_L g1960 ( 
.A1(n_1784),
.A2(n_1714),
.B(n_1723),
.C(n_1707),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1776),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1825),
.B(n_1765),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1845),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1810),
.B(n_191),
.Y(n_1964)
);

AOI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1919),
.A2(n_1698),
.B(n_1697),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1774),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1786),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1800),
.B(n_191),
.Y(n_1968)
);

A2O1A1Ixp33_ASAP7_75t_L g1969 ( 
.A1(n_1821),
.A2(n_1706),
.B(n_1704),
.C(n_196),
.Y(n_1969)
);

BUFx12f_ASAP7_75t_L g1970 ( 
.A(n_1774),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1919),
.A2(n_193),
.B(n_194),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1838),
.B(n_194),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1918),
.B(n_197),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1831),
.B(n_1795),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1844),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1914),
.Y(n_1976)
);

OAI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1847),
.A2(n_198),
.B(n_199),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1930),
.B(n_199),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1786),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_L g1980 ( 
.A1(n_1877),
.A2(n_484),
.B(n_483),
.Y(n_1980)
);

OAI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1921),
.A2(n_200),
.B(n_201),
.Y(n_1981)
);

OAI21x1_ASAP7_75t_L g1982 ( 
.A1(n_1852),
.A2(n_488),
.B(n_485),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1846),
.A2(n_200),
.B(n_201),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1815),
.A2(n_202),
.B(n_203),
.Y(n_1984)
);

OAI21x1_ASAP7_75t_L g1985 ( 
.A1(n_1908),
.A2(n_492),
.B(n_491),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1867),
.Y(n_1986)
);

NAND2xp33_ASAP7_75t_L g1987 ( 
.A(n_1836),
.B(n_202),
.Y(n_1987)
);

O2A1O1Ixp5_ASAP7_75t_L g1988 ( 
.A1(n_1772),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_1988)
);

BUFx3_ASAP7_75t_L g1989 ( 
.A(n_1774),
.Y(n_1989)
);

A2O1A1Ixp33_ASAP7_75t_L g1990 ( 
.A1(n_1783),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1781),
.A2(n_207),
.B(n_208),
.Y(n_1991)
);

NAND3xp33_ASAP7_75t_L g1992 ( 
.A(n_1807),
.B(n_207),
.C(n_208),
.Y(n_1992)
);

NAND3x1_ASAP7_75t_L g1993 ( 
.A(n_1850),
.B(n_1883),
.C(n_1775),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1841),
.Y(n_1994)
);

O2A1O1Ixp5_ASAP7_75t_L g1995 ( 
.A1(n_1842),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1926),
.B(n_209),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1869),
.B(n_210),
.Y(n_1997)
);

OAI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1915),
.A2(n_212),
.B(n_213),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1848),
.A2(n_1801),
.B(n_1856),
.Y(n_1999)
);

OA21x2_ASAP7_75t_L g2000 ( 
.A1(n_1827),
.A2(n_1782),
.B(n_1939),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1785),
.B(n_212),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1920),
.B(n_213),
.Y(n_2002)
);

OAI21xp5_ASAP7_75t_SL g2003 ( 
.A1(n_1792),
.A2(n_214),
.B(n_215),
.Y(n_2003)
);

OAI21x1_ASAP7_75t_L g2004 ( 
.A1(n_1934),
.A2(n_1872),
.B(n_1863),
.Y(n_2004)
);

AOI221x1_ASAP7_75t_L g2005 ( 
.A1(n_1898),
.A2(n_217),
.B1(n_214),
.B2(n_216),
.C(n_218),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1848),
.A2(n_216),
.B(n_217),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1854),
.Y(n_2007)
);

OAI21x1_ASAP7_75t_L g2008 ( 
.A1(n_1876),
.A2(n_496),
.B(n_494),
.Y(n_2008)
);

OAI21x1_ASAP7_75t_L g2009 ( 
.A1(n_1892),
.A2(n_498),
.B(n_497),
.Y(n_2009)
);

AO31x2_ASAP7_75t_L g2010 ( 
.A1(n_1797),
.A2(n_500),
.A3(n_504),
.B(n_499),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1861),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1899),
.B(n_1823),
.Y(n_2012)
);

AO21x2_ASAP7_75t_L g2013 ( 
.A1(n_1796),
.A2(n_506),
.B(n_505),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1813),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1823),
.B(n_218),
.Y(n_2015)
);

OAI22x1_ASAP7_75t_L g2016 ( 
.A1(n_1839),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1848),
.A2(n_219),
.B(n_220),
.Y(n_2017)
);

OAI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1812),
.A2(n_221),
.B(n_222),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1874),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1833),
.B(n_222),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1786),
.Y(n_2021)
);

OAI21x1_ASAP7_75t_L g2022 ( 
.A1(n_1912),
.A2(n_509),
.B(n_507),
.Y(n_2022)
);

CKINVDCx20_ASAP7_75t_R g2023 ( 
.A(n_1791),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1880),
.Y(n_2024)
);

AOI21xp33_ASAP7_75t_L g2025 ( 
.A1(n_1904),
.A2(n_223),
.B(n_224),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1823),
.B(n_1906),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1857),
.Y(n_2027)
);

BUFx5_ASAP7_75t_L g2028 ( 
.A(n_1823),
.Y(n_2028)
);

A2O1A1Ixp33_ASAP7_75t_L g2029 ( 
.A1(n_1888),
.A2(n_226),
.B(n_223),
.C(n_225),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1894),
.B(n_1909),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1940),
.B(n_510),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1851),
.A2(n_225),
.B(n_226),
.Y(n_2032)
);

NAND2x1p5_ASAP7_75t_L g2033 ( 
.A(n_1805),
.B(n_513),
.Y(n_2033)
);

AOI21xp5_ASAP7_75t_L g2034 ( 
.A1(n_1817),
.A2(n_227),
.B(n_229),
.Y(n_2034)
);

OA21x2_ASAP7_75t_L g2035 ( 
.A1(n_1913),
.A2(n_227),
.B(n_229),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1773),
.Y(n_2036)
);

A2O1A1Ixp33_ASAP7_75t_L g2037 ( 
.A1(n_1924),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1875),
.Y(n_2038)
);

OAI21x1_ASAP7_75t_L g2039 ( 
.A1(n_1834),
.A2(n_515),
.B(n_514),
.Y(n_2039)
);

OAI21x1_ASAP7_75t_L g2040 ( 
.A1(n_1932),
.A2(n_518),
.B(n_516),
.Y(n_2040)
);

CKINVDCx16_ASAP7_75t_R g2041 ( 
.A(n_1811),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1896),
.B(n_1818),
.Y(n_2042)
);

OAI21x1_ASAP7_75t_L g2043 ( 
.A1(n_1929),
.A2(n_1873),
.B(n_1931),
.Y(n_2043)
);

OAI21x1_ASAP7_75t_L g2044 ( 
.A1(n_1803),
.A2(n_524),
.B(n_522),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1882),
.Y(n_2045)
);

OAI21x1_ASAP7_75t_L g2046 ( 
.A1(n_1864),
.A2(n_530),
.B(n_528),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_1777),
.Y(n_2047)
);

O2A1O1Ixp33_ASAP7_75t_SL g2048 ( 
.A1(n_1881),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_2048)
);

NAND3xp33_ASAP7_75t_L g2049 ( 
.A(n_1889),
.B(n_235),
.C(n_236),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1868),
.B(n_531),
.Y(n_2050)
);

CKINVDCx6p67_ASAP7_75t_R g2051 ( 
.A(n_1862),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1895),
.Y(n_2052)
);

AOI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1925),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_2053)
);

NAND3x1_ASAP7_75t_L g2054 ( 
.A(n_1794),
.B(n_237),
.C(n_238),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1941),
.Y(n_2055)
);

AOI21x1_ASAP7_75t_L g2056 ( 
.A1(n_1905),
.A2(n_238),
.B(n_239),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1814),
.B(n_239),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_1949),
.A2(n_1960),
.B(n_1959),
.Y(n_2058)
);

OAI21x1_ASAP7_75t_L g2059 ( 
.A1(n_1943),
.A2(n_1903),
.B(n_1808),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_2028),
.B(n_1887),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2019),
.Y(n_2061)
);

OAI21x1_ASAP7_75t_L g2062 ( 
.A1(n_1965),
.A2(n_1799),
.B(n_1937),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2019),
.Y(n_2063)
);

OAI21x1_ASAP7_75t_L g2064 ( 
.A1(n_2004),
.A2(n_1902),
.B(n_1936),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2045),
.Y(n_2065)
);

O2A1O1Ixp33_ASAP7_75t_SL g2066 ( 
.A1(n_2003),
.A2(n_1911),
.B(n_1802),
.C(n_1853),
.Y(n_2066)
);

NAND3xp33_ASAP7_75t_L g2067 ( 
.A(n_2037),
.B(n_1927),
.C(n_1849),
.Y(n_2067)
);

OA21x2_ASAP7_75t_L g2068 ( 
.A1(n_1999),
.A2(n_1910),
.B(n_1822),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_2055),
.B(n_1887),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_2014),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2045),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1954),
.A2(n_1923),
.B(n_1885),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1951),
.Y(n_2073)
);

OAI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_2053),
.A2(n_1884),
.B1(n_1916),
.B2(n_1923),
.Y(n_2074)
);

O2A1O1Ixp33_ASAP7_75t_L g2075 ( 
.A1(n_1987),
.A2(n_1901),
.B(n_1897),
.C(n_1891),
.Y(n_2075)
);

OAI211xp5_ASAP7_75t_L g2076 ( 
.A1(n_1998),
.A2(n_2018),
.B(n_2005),
.C(n_1977),
.Y(n_2076)
);

OAI21x1_ASAP7_75t_L g2077 ( 
.A1(n_1957),
.A2(n_1826),
.B(n_1820),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2038),
.Y(n_2078)
);

OAI21x1_ASAP7_75t_L g2079 ( 
.A1(n_1952),
.A2(n_1837),
.B(n_1835),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_2055),
.B(n_1887),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_1947),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1948),
.B(n_1798),
.Y(n_2082)
);

CKINVDCx6p67_ASAP7_75t_R g2083 ( 
.A(n_1970),
.Y(n_2083)
);

OAI21x1_ASAP7_75t_L g2084 ( 
.A1(n_1952),
.A2(n_1864),
.B(n_1819),
.Y(n_2084)
);

OAI21x1_ASAP7_75t_L g2085 ( 
.A1(n_1982),
.A2(n_1917),
.B(n_1855),
.Y(n_2085)
);

CKINVDCx20_ASAP7_75t_R g2086 ( 
.A(n_2023),
.Y(n_2086)
);

BUFx2_ASAP7_75t_L g2087 ( 
.A(n_1966),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1955),
.Y(n_2088)
);

OAI21x1_ASAP7_75t_L g2089 ( 
.A1(n_1985),
.A2(n_1858),
.B(n_1840),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_2015),
.B(n_1866),
.Y(n_2090)
);

AOI22xp33_ASAP7_75t_L g2091 ( 
.A1(n_1992),
.A2(n_1886),
.B1(n_1790),
.B2(n_1879),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1956),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1963),
.Y(n_2093)
);

BUFx8_ASAP7_75t_SL g2094 ( 
.A(n_2036),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_L g2095 ( 
.A1(n_2008),
.A2(n_1870),
.B(n_1938),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_1989),
.Y(n_2096)
);

OAI21x1_ASAP7_75t_L g2097 ( 
.A1(n_1983),
.A2(n_1843),
.B(n_1893),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1961),
.Y(n_2098)
);

OAI21xp5_ASAP7_75t_L g2099 ( 
.A1(n_1984),
.A2(n_1988),
.B(n_1991),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_2051),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1986),
.B(n_1922),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2007),
.Y(n_2102)
);

AO21x2_ASAP7_75t_L g2103 ( 
.A1(n_1950),
.A2(n_1878),
.B(n_1809),
.Y(n_2103)
);

AOI21xp5_ASAP7_75t_L g2104 ( 
.A1(n_1962),
.A2(n_1907),
.B(n_1928),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_1958),
.B(n_1922),
.Y(n_2105)
);

INVx3_ASAP7_75t_L g2106 ( 
.A(n_2028),
.Y(n_2106)
);

OAI21x1_ASAP7_75t_L g2107 ( 
.A1(n_2009),
.A2(n_1804),
.B(n_1907),
.Y(n_2107)
);

INVx2_ASAP7_75t_SL g2108 ( 
.A(n_2027),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2030),
.B(n_1865),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2011),
.Y(n_2110)
);

AO32x2_ASAP7_75t_L g2111 ( 
.A1(n_1974),
.A2(n_1900),
.A3(n_1788),
.B1(n_1890),
.B2(n_1933),
.Y(n_2111)
);

O2A1O1Ixp33_ASAP7_75t_SL g2112 ( 
.A1(n_2029),
.A2(n_1778),
.B(n_242),
.C(n_240),
.Y(n_2112)
);

AOI21xp33_ASAP7_75t_L g2113 ( 
.A1(n_2000),
.A2(n_1890),
.B(n_1805),
.Y(n_2113)
);

OAI221xp5_ASAP7_75t_L g2114 ( 
.A1(n_1990),
.A2(n_1890),
.B1(n_1805),
.B2(n_1933),
.C(n_1942),
.Y(n_2114)
);

OR2x6_ASAP7_75t_L g2115 ( 
.A(n_2026),
.B(n_1942),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_2012),
.B(n_1976),
.Y(n_2116)
);

AO21x2_ASAP7_75t_L g2117 ( 
.A1(n_1945),
.A2(n_2013),
.B(n_1981),
.Y(n_2117)
);

CKINVDCx11_ASAP7_75t_R g2118 ( 
.A(n_1975),
.Y(n_2118)
);

OAI21x1_ASAP7_75t_L g2119 ( 
.A1(n_2022),
.A2(n_1942),
.B(n_534),
.Y(n_2119)
);

OAI21x1_ASAP7_75t_L g2120 ( 
.A1(n_1980),
.A2(n_536),
.B(n_533),
.Y(n_2120)
);

AO21x2_ASAP7_75t_L g2121 ( 
.A1(n_2025),
.A2(n_241),
.B(n_242),
.Y(n_2121)
);

O2A1O1Ixp33_ASAP7_75t_L g2122 ( 
.A1(n_2048),
.A2(n_244),
.B(n_241),
.C(n_243),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_1976),
.Y(n_2123)
);

A2O1A1Ixp33_ASAP7_75t_L g2124 ( 
.A1(n_1995),
.A2(n_245),
.B(n_243),
.C(n_244),
.Y(n_2124)
);

INVx1_ASAP7_75t_SL g2125 ( 
.A(n_2042),
.Y(n_2125)
);

INVx2_ASAP7_75t_SL g2126 ( 
.A(n_1967),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2024),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_1953),
.B(n_246),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2052),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2001),
.B(n_1972),
.Y(n_2130)
);

OAI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_2074),
.A2(n_2041),
.B1(n_2000),
.B2(n_2035),
.Y(n_2131)
);

INVx1_ASAP7_75t_SL g2132 ( 
.A(n_2118),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2081),
.B(n_1964),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2110),
.Y(n_2134)
);

BUFx8_ASAP7_75t_L g2135 ( 
.A(n_2128),
.Y(n_2135)
);

INVxp67_ASAP7_75t_L g2136 ( 
.A(n_2081),
.Y(n_2136)
);

AOI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_2067),
.A2(n_2016),
.B1(n_2035),
.B2(n_2049),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2110),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_SL g2139 ( 
.A1(n_2117),
.A2(n_2028),
.B1(n_1944),
.B2(n_1993),
.Y(n_2139)
);

AOI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_2091),
.A2(n_2002),
.B1(n_2057),
.B2(n_1973),
.Y(n_2140)
);

INVx6_ASAP7_75t_L g2141 ( 
.A(n_2105),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2127),
.Y(n_2142)
);

AOI22xp5_ASAP7_75t_SL g2143 ( 
.A1(n_2086),
.A2(n_2100),
.B1(n_2090),
.B2(n_2130),
.Y(n_2143)
);

AOI22xp33_ASAP7_75t_SL g2144 ( 
.A1(n_2117),
.A2(n_2028),
.B1(n_1944),
.B2(n_1946),
.Y(n_2144)
);

INVx2_ASAP7_75t_SL g2145 ( 
.A(n_2087),
.Y(n_2145)
);

INVx4_ASAP7_75t_L g2146 ( 
.A(n_2100),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2127),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2061),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2091),
.A2(n_2099),
.B1(n_2072),
.B2(n_2068),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2078),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2063),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_L g2152 ( 
.A1(n_2068),
.A2(n_2032),
.B1(n_2017),
.B2(n_2006),
.Y(n_2152)
);

CKINVDCx11_ASAP7_75t_R g2153 ( 
.A(n_2086),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2065),
.Y(n_2154)
);

CKINVDCx11_ASAP7_75t_R g2155 ( 
.A(n_2118),
.Y(n_2155)
);

BUFx2_ASAP7_75t_SL g2156 ( 
.A(n_2108),
.Y(n_2156)
);

INVx6_ASAP7_75t_L g2157 ( 
.A(n_2105),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2071),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2078),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2123),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2123),
.Y(n_2161)
);

AND2x4_ASAP7_75t_L g2162 ( 
.A(n_2106),
.B(n_1953),
.Y(n_2162)
);

OAI21xp5_ASAP7_75t_L g2163 ( 
.A1(n_2076),
.A2(n_2054),
.B(n_1971),
.Y(n_2163)
);

OAI22xp33_ASAP7_75t_SL g2164 ( 
.A1(n_2082),
.A2(n_1994),
.B1(n_1996),
.B2(n_1997),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2073),
.Y(n_2165)
);

AOI21x1_ASAP7_75t_L g2166 ( 
.A1(n_2058),
.A2(n_1968),
.B(n_1978),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2088),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2098),
.Y(n_2168)
);

INVx3_ASAP7_75t_L g2169 ( 
.A(n_2116),
.Y(n_2169)
);

OAI21x1_ASAP7_75t_L g2170 ( 
.A1(n_2084),
.A2(n_2043),
.B(n_2046),
.Y(n_2170)
);

INVx2_ASAP7_75t_SL g2171 ( 
.A(n_2096),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_2068),
.A2(n_2028),
.B1(n_1946),
.B2(n_2031),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2098),
.Y(n_2173)
);

OAI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_2124),
.A2(n_2034),
.B(n_1969),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2092),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2093),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2070),
.B(n_2020),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2116),
.B(n_1946),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2102),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_L g2180 ( 
.A1(n_2090),
.A2(n_1946),
.B1(n_2047),
.B2(n_1979),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2129),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2169),
.B(n_2116),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2142),
.Y(n_2183)
);

INVx2_ASAP7_75t_SL g2184 ( 
.A(n_2141),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2160),
.Y(n_2185)
);

INVxp67_ASAP7_75t_L g2186 ( 
.A(n_2156),
.Y(n_2186)
);

AOI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_2131),
.A2(n_2112),
.B1(n_2066),
.B2(n_2121),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2169),
.B(n_2125),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2161),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2142),
.Y(n_2190)
);

BUFx4f_ASAP7_75t_L g2191 ( 
.A(n_2141),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2150),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2149),
.A2(n_2124),
.B1(n_2128),
.B2(n_2104),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2169),
.B(n_2109),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_L g2195 ( 
.A1(n_2149),
.A2(n_2128),
.B1(n_2075),
.B2(n_2122),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2134),
.Y(n_2196)
);

AOI22xp33_ASAP7_75t_L g2197 ( 
.A1(n_2163),
.A2(n_2103),
.B1(n_2121),
.B2(n_2113),
.Y(n_2197)
);

CKINVDCx11_ASAP7_75t_R g2198 ( 
.A(n_2153),
.Y(n_2198)
);

OAI21xp5_ASAP7_75t_SL g2199 ( 
.A1(n_2137),
.A2(n_2056),
.B(n_2105),
.Y(n_2199)
);

OAI22xp33_ASAP7_75t_L g2200 ( 
.A1(n_2178),
.A2(n_2174),
.B1(n_2166),
.B2(n_2114),
.Y(n_2200)
);

BUFx2_ASAP7_75t_L g2201 ( 
.A(n_2135),
.Y(n_2201)
);

INVx4_ASAP7_75t_SL g2202 ( 
.A(n_2141),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_2137),
.A2(n_2103),
.B1(n_2095),
.B2(n_2079),
.Y(n_2203)
);

INVx5_ASAP7_75t_L g2204 ( 
.A(n_2146),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2138),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_2153),
.Y(n_2206)
);

CKINVDCx20_ASAP7_75t_R g2207 ( 
.A(n_2155),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_2182),
.B(n_2145),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2182),
.B(n_2171),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_R g2210 ( 
.A(n_2207),
.B(n_2155),
.Y(n_2210)
);

OR2x6_ASAP7_75t_L g2211 ( 
.A(n_2199),
.B(n_2060),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2194),
.B(n_2184),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2196),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2202),
.B(n_2162),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2194),
.B(n_2177),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_2201),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2185),
.B(n_2181),
.Y(n_2217)
);

AND2x4_ASAP7_75t_L g2218 ( 
.A(n_2202),
.B(n_2162),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2196),
.Y(n_2219)
);

BUFx3_ASAP7_75t_L g2220 ( 
.A(n_2198),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2217),
.B(n_2133),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2212),
.B(n_2201),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2213),
.Y(n_2223)
);

BUFx3_ASAP7_75t_L g2224 ( 
.A(n_2220),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2213),
.B(n_2185),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2215),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2222),
.B(n_2214),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2223),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2221),
.B(n_2216),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2226),
.B(n_2214),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2224),
.A2(n_2187),
.B1(n_2193),
.B2(n_2200),
.Y(n_2231)
);

HB1xp67_ASAP7_75t_L g2232 ( 
.A(n_2225),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2223),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2224),
.Y(n_2234)
);

BUFx3_ASAP7_75t_L g2235 ( 
.A(n_2225),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2223),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2236),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2227),
.B(n_2220),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2236),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2235),
.B(n_2215),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2228),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2228),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2233),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2232),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2235),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2234),
.Y(n_2246)
);

INVx2_ASAP7_75t_SL g2247 ( 
.A(n_2234),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2230),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2247),
.B(n_2231),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2238),
.B(n_2220),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2247),
.B(n_2229),
.Y(n_2251)
);

AND2x4_ASAP7_75t_L g2252 ( 
.A(n_2238),
.B(n_2227),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_2248),
.B(n_2230),
.Y(n_2253)
);

AND2x4_ASAP7_75t_L g2254 ( 
.A(n_2248),
.B(n_2206),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2241),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2240),
.B(n_2217),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2246),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2250),
.B(n_2245),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_2253),
.B(n_2246),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2253),
.B(n_2244),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2257),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2259),
.B(n_2252),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2258),
.B(n_2252),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2260),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_2261),
.B(n_2254),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2263),
.Y(n_2266)
);

OAI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2262),
.A2(n_2251),
.B1(n_2249),
.B2(n_2254),
.Y(n_2267)
);

AO22x2_ASAP7_75t_L g2268 ( 
.A1(n_2265),
.A2(n_2255),
.B1(n_2237),
.B2(n_2239),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2264),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2263),
.Y(n_2270)
);

AOI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2265),
.A2(n_2243),
.B1(n_2242),
.B2(n_2255),
.Y(n_2271)
);

NAND3xp33_ASAP7_75t_SL g2272 ( 
.A(n_2267),
.B(n_2256),
.C(n_2210),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2266),
.B(n_2206),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2268),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2270),
.A2(n_2211),
.B1(n_2195),
.B2(n_2140),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2271),
.B(n_2269),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2268),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2268),
.B(n_2143),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_2266),
.B(n_2132),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2268),
.Y(n_2280)
);

NAND2x1_ASAP7_75t_L g2281 ( 
.A(n_2268),
.B(n_2146),
.Y(n_2281)
);

NOR4xp25_ASAP7_75t_L g2282 ( 
.A(n_2274),
.B(n_2140),
.C(n_2112),
.D(n_2186),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2278),
.A2(n_2279),
.B1(n_2276),
.B2(n_2277),
.Y(n_2283)
);

OAI22xp33_ASAP7_75t_SL g2284 ( 
.A1(n_2280),
.A2(n_2211),
.B1(n_2146),
.B2(n_2204),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2273),
.B(n_2212),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2275),
.B(n_2219),
.Y(n_2286)
);

AOI221xp5_ASAP7_75t_L g2287 ( 
.A1(n_2272),
.A2(n_2197),
.B1(n_2203),
.B2(n_2066),
.C(n_2164),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_2281),
.B(n_2204),
.Y(n_2288)
);

AOI221xp5_ASAP7_75t_L g2289 ( 
.A1(n_2274),
.A2(n_2152),
.B1(n_2219),
.B2(n_2139),
.C(n_2172),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2273),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2273),
.B(n_2211),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_L g2292 ( 
.A(n_2281),
.B(n_2094),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_2281),
.A2(n_2211),
.B(n_2094),
.Y(n_2293)
);

INVxp67_ASAP7_75t_SL g2294 ( 
.A(n_2273),
.Y(n_2294)
);

AOI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2294),
.A2(n_2211),
.B(n_2214),
.Y(n_2295)
);

INVxp67_ASAP7_75t_L g2296 ( 
.A(n_2292),
.Y(n_2296)
);

NOR3x1_ASAP7_75t_L g2297 ( 
.A(n_2283),
.B(n_2083),
.C(n_2189),
.Y(n_2297)
);

NAND4xp25_ASAP7_75t_L g2298 ( 
.A(n_2293),
.B(n_2214),
.C(n_2218),
.D(n_2152),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2290),
.Y(n_2299)
);

BUFx2_ASAP7_75t_L g2300 ( 
.A(n_2285),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2291),
.B(n_2204),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2282),
.B(n_2218),
.Y(n_2302)
);

AOI211xp5_ASAP7_75t_L g2303 ( 
.A1(n_2284),
.A2(n_2218),
.B(n_2085),
.C(n_2089),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_2286),
.B(n_2204),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2288),
.B(n_2208),
.Y(n_2305)
);

AOI221xp5_ASAP7_75t_L g2306 ( 
.A1(n_2287),
.A2(n_2289),
.B1(n_2172),
.B2(n_2218),
.C(n_2144),
.Y(n_2306)
);

NOR4xp75_ASAP7_75t_L g2307 ( 
.A(n_2283),
.B(n_2209),
.C(n_2208),
.D(n_2204),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2285),
.Y(n_2308)
);

NOR3xp33_ASAP7_75t_L g2309 ( 
.A(n_2283),
.B(n_2089),
.C(n_2085),
.Y(n_2309)
);

O2A1O1Ixp33_ASAP7_75t_L g2310 ( 
.A1(n_2299),
.A2(n_2033),
.B(n_250),
.C(n_246),
.Y(n_2310)
);

NAND3xp33_ASAP7_75t_L g2311 ( 
.A(n_2300),
.B(n_2204),
.C(n_2135),
.Y(n_2311)
);

AOI22xp33_ASAP7_75t_SL g2312 ( 
.A1(n_2302),
.A2(n_2135),
.B1(n_2095),
.B2(n_1979),
.Y(n_2312)
);

AOI21xp33_ASAP7_75t_L g2313 ( 
.A1(n_2296),
.A2(n_2301),
.B(n_2308),
.Y(n_2313)
);

NOR4xp25_ASAP7_75t_L g2314 ( 
.A(n_2304),
.B(n_2188),
.C(n_2189),
.D(n_2209),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2295),
.B(n_2136),
.Y(n_2315)
);

OAI221xp5_ASAP7_75t_SL g2316 ( 
.A1(n_2309),
.A2(n_2180),
.B1(n_2184),
.B2(n_2101),
.C(n_2175),
.Y(n_2316)
);

NOR3xp33_ASAP7_75t_L g2317 ( 
.A(n_2306),
.B(n_2050),
.C(n_2077),
.Y(n_2317)
);

OAI221xp5_ASAP7_75t_L g2318 ( 
.A1(n_2303),
.A2(n_2298),
.B1(n_2305),
.B2(n_2307),
.C(n_2297),
.Y(n_2318)
);

NOR3xp33_ASAP7_75t_L g2319 ( 
.A(n_2299),
.B(n_2050),
.C(n_2120),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2300),
.B(n_2202),
.Y(n_2320)
);

OAI211xp5_ASAP7_75t_L g2321 ( 
.A1(n_2300),
.A2(n_251),
.B(n_248),
.C(n_250),
.Y(n_2321)
);

AOI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2302),
.A2(n_2188),
.B1(n_1979),
.B2(n_2021),
.Y(n_2322)
);

OAI211xp5_ASAP7_75t_L g2323 ( 
.A1(n_2300),
.A2(n_253),
.B(n_248),
.C(n_252),
.Y(n_2323)
);

A2O1A1Ixp33_ASAP7_75t_L g2324 ( 
.A1(n_2310),
.A2(n_2318),
.B(n_2313),
.C(n_2322),
.Y(n_2324)
);

AOI222xp33_ASAP7_75t_L g2325 ( 
.A1(n_2315),
.A2(n_2320),
.B1(n_2323),
.B2(n_2321),
.C1(n_2311),
.C2(n_2317),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2314),
.B(n_2205),
.Y(n_2326)
);

AOI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2312),
.A2(n_2205),
.B1(n_2176),
.B2(n_2179),
.C(n_2167),
.Y(n_2327)
);

AOI221xp5_ASAP7_75t_L g2328 ( 
.A1(n_2316),
.A2(n_2165),
.B1(n_2154),
.B2(n_2158),
.C(n_2151),
.Y(n_2328)
);

O2A1O1Ixp33_ASAP7_75t_L g2329 ( 
.A1(n_2319),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2320),
.B(n_2202),
.Y(n_2330)
);

NAND3xp33_ASAP7_75t_SL g2331 ( 
.A(n_2321),
.B(n_2180),
.C(n_254),
.Y(n_2331)
);

OAI21xp33_ASAP7_75t_L g2332 ( 
.A1(n_2311),
.A2(n_2162),
.B(n_2148),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2314),
.B(n_255),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2314),
.B(n_256),
.Y(n_2334)
);

AOI211x1_ASAP7_75t_SL g2335 ( 
.A1(n_2313),
.A2(n_258),
.B(n_256),
.C(n_257),
.Y(n_2335)
);

AOI221xp5_ASAP7_75t_L g2336 ( 
.A1(n_2318),
.A2(n_2190),
.B1(n_2183),
.B2(n_2192),
.C(n_260),
.Y(n_2336)
);

OAI211xp5_ASAP7_75t_SL g2337 ( 
.A1(n_2313),
.A2(n_261),
.B(n_257),
.C(n_259),
.Y(n_2337)
);

NAND3xp33_ASAP7_75t_L g2338 ( 
.A(n_2313),
.B(n_2021),
.C(n_1967),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2320),
.A2(n_261),
.B(n_262),
.Y(n_2339)
);

NAND3xp33_ASAP7_75t_L g2340 ( 
.A(n_2313),
.B(n_2021),
.C(n_1967),
.Y(n_2340)
);

NOR3xp33_ASAP7_75t_L g2341 ( 
.A(n_2313),
.B(n_2097),
.C(n_2039),
.Y(n_2341)
);

OAI22xp33_ASAP7_75t_L g2342 ( 
.A1(n_2322),
.A2(n_2191),
.B1(n_2190),
.B2(n_2183),
.Y(n_2342)
);

AOI322xp5_ASAP7_75t_L g2343 ( 
.A1(n_2317),
.A2(n_2010),
.A3(n_2192),
.B1(n_2060),
.B2(n_2080),
.C1(n_2069),
.C2(n_2126),
.Y(n_2343)
);

NAND4xp25_ASAP7_75t_L g2344 ( 
.A(n_2313),
.B(n_264),
.C(n_262),
.D(n_263),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2314),
.B(n_263),
.Y(n_2345)
);

OAI22xp33_ASAP7_75t_L g2346 ( 
.A1(n_2333),
.A2(n_2191),
.B1(n_2106),
.B2(n_2157),
.Y(n_2346)
);

OR2x2_ASAP7_75t_L g2347 ( 
.A(n_2334),
.B(n_265),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_L g2348 ( 
.A(n_2345),
.B(n_265),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2344),
.B(n_266),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2335),
.Y(n_2350)
);

AOI21xp33_ASAP7_75t_L g2351 ( 
.A1(n_2325),
.A2(n_267),
.B(n_268),
.Y(n_2351)
);

NAND4xp25_ASAP7_75t_L g2352 ( 
.A(n_2324),
.B(n_270),
.C(n_267),
.D(n_269),
.Y(n_2352)
);

O2A1O1Ixp5_ASAP7_75t_L g2353 ( 
.A1(n_2339),
.A2(n_272),
.B(n_269),
.C(n_271),
.Y(n_2353)
);

NAND2xp33_ASAP7_75t_SL g2354 ( 
.A(n_2330),
.B(n_272),
.Y(n_2354)
);

OAI321xp33_ASAP7_75t_L g2355 ( 
.A1(n_2336),
.A2(n_2147),
.A3(n_2115),
.B1(n_275),
.B2(n_276),
.C(n_277),
.Y(n_2355)
);

NOR3xp33_ASAP7_75t_L g2356 ( 
.A(n_2337),
.B(n_273),
.C(n_274),
.Y(n_2356)
);

OAI221xp5_ASAP7_75t_SL g2357 ( 
.A1(n_2329),
.A2(n_274),
.B1(n_277),
.B2(n_278),
.C(n_279),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2326),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2331),
.Y(n_2359)
);

AOI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_2341),
.A2(n_2170),
.B1(n_2107),
.B2(n_2064),
.Y(n_2360)
);

AOI221xp5_ASAP7_75t_L g2361 ( 
.A1(n_2342),
.A2(n_278),
.B1(n_279),
.B2(n_280),
.C(n_281),
.Y(n_2361)
);

INVx1_ASAP7_75t_SL g2362 ( 
.A(n_2338),
.Y(n_2362)
);

AOI211xp5_ASAP7_75t_L g2363 ( 
.A1(n_2340),
.A2(n_282),
.B(n_280),
.C(n_281),
.Y(n_2363)
);

OAI211xp5_ASAP7_75t_L g2364 ( 
.A1(n_2327),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_2364)
);

A2O1A1O1Ixp25_ASAP7_75t_L g2365 ( 
.A1(n_2332),
.A2(n_283),
.B(n_285),
.C(n_286),
.D(n_287),
.Y(n_2365)
);

AOI322xp5_ASAP7_75t_L g2366 ( 
.A1(n_2343),
.A2(n_2010),
.A3(n_2069),
.B1(n_2080),
.B2(n_2062),
.C1(n_2159),
.C2(n_2173),
.Y(n_2366)
);

AOI211xp5_ASAP7_75t_L g2367 ( 
.A1(n_2328),
.A2(n_288),
.B(n_285),
.C(n_286),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_2333),
.B(n_288),
.Y(n_2368)
);

OAI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_2324),
.A2(n_2044),
.B(n_2107),
.Y(n_2369)
);

NOR2x1p5_ASAP7_75t_L g2370 ( 
.A(n_2344),
.B(n_289),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2335),
.B(n_289),
.Y(n_2371)
);

AOI211xp5_ASAP7_75t_L g2372 ( 
.A1(n_2333),
.A2(n_292),
.B(n_290),
.C(n_291),
.Y(n_2372)
);

O2A1O1Ixp33_ASAP7_75t_L g2373 ( 
.A1(n_2324),
.A2(n_293),
.B(n_290),
.C(n_292),
.Y(n_2373)
);

AOI311xp33_ASAP7_75t_L g2374 ( 
.A1(n_2324),
.A2(n_293),
.A3(n_294),
.B(n_295),
.C(n_296),
.Y(n_2374)
);

OAI211xp5_ASAP7_75t_L g2375 ( 
.A1(n_2333),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_2375)
);

AOI221xp5_ASAP7_75t_L g2376 ( 
.A1(n_2333),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.C(n_300),
.Y(n_2376)
);

A2O1A1Ixp33_ASAP7_75t_L g2377 ( 
.A1(n_2339),
.A2(n_2170),
.B(n_2040),
.C(n_2191),
.Y(n_2377)
);

OAI211xp5_ASAP7_75t_L g2378 ( 
.A1(n_2333),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_2378)
);

OAI211xp5_ASAP7_75t_L g2379 ( 
.A1(n_2333),
.A2(n_304),
.B(n_301),
.C(n_302),
.Y(n_2379)
);

CKINVDCx20_ASAP7_75t_R g2380 ( 
.A(n_2333),
.Y(n_2380)
);

AOI221xp5_ASAP7_75t_L g2381 ( 
.A1(n_2333),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.C(n_307),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2330),
.B(n_2157),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2374),
.B(n_2157),
.Y(n_2383)
);

BUFx5_ASAP7_75t_L g2384 ( 
.A(n_2359),
.Y(n_2384)
);

AOI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2380),
.A2(n_2059),
.B1(n_2119),
.B2(n_2084),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2371),
.Y(n_2386)
);

NOR2x1_ASAP7_75t_L g2387 ( 
.A(n_2352),
.B(n_305),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2382),
.B(n_306),
.Y(n_2388)
);

AND4x1_ASAP7_75t_L g2389 ( 
.A(n_2372),
.B(n_2348),
.C(n_2363),
.D(n_2353),
.Y(n_2389)
);

AOI21xp5_ASAP7_75t_L g2390 ( 
.A1(n_2373),
.A2(n_307),
.B(n_308),
.Y(n_2390)
);

NOR3x1_ASAP7_75t_L g2391 ( 
.A(n_2375),
.B(n_309),
.C(n_311),
.Y(n_2391)
);

AND2x4_ASAP7_75t_L g2392 ( 
.A(n_2370),
.B(n_2362),
.Y(n_2392)
);

NOR2x1_ASAP7_75t_L g2393 ( 
.A(n_2358),
.B(n_309),
.Y(n_2393)
);

NAND3xp33_ASAP7_75t_SL g2394 ( 
.A(n_2350),
.B(n_2362),
.C(n_2376),
.Y(n_2394)
);

NOR2xp67_ASAP7_75t_SL g2395 ( 
.A(n_2347),
.B(n_311),
.Y(n_2395)
);

NAND3xp33_ASAP7_75t_L g2396 ( 
.A(n_2354),
.B(n_2351),
.C(n_2381),
.Y(n_2396)
);

INVx2_ASAP7_75t_SL g2397 ( 
.A(n_2368),
.Y(n_2397)
);

NOR2xp67_ASAP7_75t_L g2398 ( 
.A(n_2364),
.B(n_313),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2349),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2356),
.B(n_313),
.Y(n_2400)
);

NAND4xp75_ASAP7_75t_L g2401 ( 
.A(n_2361),
.B(n_314),
.C(n_315),
.D(n_316),
.Y(n_2401)
);

NAND3xp33_ASAP7_75t_L g2402 ( 
.A(n_2365),
.B(n_314),
.C(n_315),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2378),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2360),
.Y(n_2404)
);

NOR3x2_ASAP7_75t_L g2405 ( 
.A(n_2357),
.B(n_316),
.C(n_317),
.Y(n_2405)
);

OR2x2_ASAP7_75t_L g2406 ( 
.A(n_2379),
.B(n_317),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2367),
.Y(n_2407)
);

NOR3x1_ASAP7_75t_L g2408 ( 
.A(n_2369),
.B(n_2355),
.C(n_2346),
.Y(n_2408)
);

NAND3xp33_ASAP7_75t_L g2409 ( 
.A(n_2377),
.B(n_2366),
.C(n_318),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_2371),
.B(n_318),
.Y(n_2410)
);

AOI22xp5_ASAP7_75t_L g2411 ( 
.A1(n_2380),
.A2(n_2059),
.B1(n_2069),
.B2(n_2080),
.Y(n_2411)
);

NAND3xp33_ASAP7_75t_L g2412 ( 
.A(n_2348),
.B(n_319),
.C(n_320),
.Y(n_2412)
);

NAND4xp75_ASAP7_75t_L g2413 ( 
.A(n_2351),
.B(n_320),
.C(n_321),
.D(n_322),
.Y(n_2413)
);

NOR2x1_ASAP7_75t_L g2414 ( 
.A(n_2352),
.B(n_322),
.Y(n_2414)
);

NOR2x1_ASAP7_75t_L g2415 ( 
.A(n_2394),
.B(n_323),
.Y(n_2415)
);

NOR2x1_ASAP7_75t_SL g2416 ( 
.A(n_2401),
.B(n_325),
.Y(n_2416)
);

NOR2x1_ASAP7_75t_L g2417 ( 
.A(n_2410),
.B(n_326),
.Y(n_2417)
);

NOR2x1_ASAP7_75t_L g2418 ( 
.A(n_2392),
.B(n_326),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2391),
.Y(n_2419)
);

NAND3x1_ASAP7_75t_SL g2420 ( 
.A(n_2393),
.B(n_327),
.C(n_328),
.Y(n_2420)
);

AND2x4_ASAP7_75t_L g2421 ( 
.A(n_2383),
.B(n_2388),
.Y(n_2421)
);

OR2x2_ASAP7_75t_L g2422 ( 
.A(n_2402),
.B(n_2406),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2384),
.B(n_327),
.Y(n_2423)
);

NAND2x1_ASAP7_75t_SL g2424 ( 
.A(n_2387),
.B(n_328),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2395),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2384),
.Y(n_2426)
);

INVxp67_ASAP7_75t_L g2427 ( 
.A(n_2397),
.Y(n_2427)
);

NOR3xp33_ASAP7_75t_L g2428 ( 
.A(n_2386),
.B(n_329),
.C(n_330),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2384),
.Y(n_2429)
);

NOR2x1_ASAP7_75t_L g2430 ( 
.A(n_2412),
.B(n_329),
.Y(n_2430)
);

NOR2x1_ASAP7_75t_L g2431 ( 
.A(n_2413),
.B(n_2403),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_SL g2432 ( 
.A(n_2384),
.B(n_330),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_2389),
.B(n_331),
.Y(n_2433)
);

NOR2x1_ASAP7_75t_L g2434 ( 
.A(n_2399),
.B(n_332),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2414),
.B(n_332),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2405),
.Y(n_2436)
);

NOR2x1_ASAP7_75t_L g2437 ( 
.A(n_2396),
.B(n_333),
.Y(n_2437)
);

OR2x2_ASAP7_75t_L g2438 ( 
.A(n_2400),
.B(n_334),
.Y(n_2438)
);

NAND2x1p5_ASAP7_75t_L g2439 ( 
.A(n_2407),
.B(n_335),
.Y(n_2439)
);

NOR3xp33_ASAP7_75t_SL g2440 ( 
.A(n_2390),
.B(n_335),
.C(n_336),
.Y(n_2440)
);

OR2x2_ASAP7_75t_L g2441 ( 
.A(n_2398),
.B(n_336),
.Y(n_2441)
);

NAND4xp75_ASAP7_75t_L g2442 ( 
.A(n_2408),
.B(n_337),
.C(n_338),
.D(n_339),
.Y(n_2442)
);

NOR2x1p5_ASAP7_75t_L g2443 ( 
.A(n_2404),
.B(n_337),
.Y(n_2443)
);

NOR2xp67_ASAP7_75t_SL g2444 ( 
.A(n_2409),
.B(n_339),
.Y(n_2444)
);

NOR2x1_ASAP7_75t_L g2445 ( 
.A(n_2411),
.B(n_341),
.Y(n_2445)
);

NOR2x1_ASAP7_75t_L g2446 ( 
.A(n_2385),
.B(n_342),
.Y(n_2446)
);

NOR2xp67_ASAP7_75t_L g2447 ( 
.A(n_2402),
.B(n_342),
.Y(n_2447)
);

NOR3xp33_ASAP7_75t_SL g2448 ( 
.A(n_2394),
.B(n_344),
.C(n_345),
.Y(n_2448)
);

NAND3x2_ASAP7_75t_L g2449 ( 
.A(n_2399),
.B(n_344),
.C(n_345),
.Y(n_2449)
);

INVx3_ASAP7_75t_SL g2450 ( 
.A(n_2384),
.Y(n_2450)
);

NOR2x1_ASAP7_75t_L g2451 ( 
.A(n_2394),
.B(n_346),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2384),
.B(n_346),
.Y(n_2452)
);

NAND3x1_ASAP7_75t_SL g2453 ( 
.A(n_2393),
.B(n_347),
.C(n_348),
.Y(n_2453)
);

NAND3xp33_ASAP7_75t_SL g2454 ( 
.A(n_2410),
.B(n_349),
.C(n_350),
.Y(n_2454)
);

AND2x4_ASAP7_75t_L g2455 ( 
.A(n_2392),
.B(n_349),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2384),
.B(n_350),
.Y(n_2456)
);

OR2x2_ASAP7_75t_L g2457 ( 
.A(n_2402),
.B(n_351),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_2384),
.B(n_351),
.Y(n_2458)
);

NAND4xp75_ASAP7_75t_L g2459 ( 
.A(n_2393),
.B(n_352),
.C(n_353),
.D(n_354),
.Y(n_2459)
);

NAND4xp75_ASAP7_75t_L g2460 ( 
.A(n_2393),
.B(n_352),
.C(n_353),
.D(n_355),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2393),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2450),
.B(n_356),
.Y(n_2462)
);

AND2x4_ASAP7_75t_L g2463 ( 
.A(n_2421),
.B(n_356),
.Y(n_2463)
);

AOI22xp33_ASAP7_75t_L g2464 ( 
.A1(n_2419),
.A2(n_2173),
.B1(n_2168),
.B2(n_2159),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2424),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2434),
.B(n_357),
.Y(n_2466)
);

AND2x4_ASAP7_75t_L g2467 ( 
.A(n_2421),
.B(n_357),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2461),
.B(n_358),
.Y(n_2468)
);

AOI221xp5_ASAP7_75t_L g2469 ( 
.A1(n_2427),
.A2(n_358),
.B1(n_359),
.B2(n_360),
.C(n_361),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2418),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2420),
.Y(n_2471)
);

NOR3xp33_ASAP7_75t_L g2472 ( 
.A(n_2426),
.B(n_359),
.C(n_360),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2439),
.Y(n_2473)
);

OAI221xp5_ASAP7_75t_L g2474 ( 
.A1(n_2429),
.A2(n_361),
.B1(n_363),
.B2(n_364),
.C(n_365),
.Y(n_2474)
);

NAND3xp33_ASAP7_75t_L g2475 ( 
.A(n_2415),
.B(n_363),
.C(n_365),
.Y(n_2475)
);

NOR3x1_ASAP7_75t_L g2476 ( 
.A(n_2442),
.B(n_366),
.C(n_367),
.Y(n_2476)
);

NAND4xp75_ASAP7_75t_L g2477 ( 
.A(n_2451),
.B(n_367),
.C(n_368),
.D(n_369),
.Y(n_2477)
);

NOR3xp33_ASAP7_75t_L g2478 ( 
.A(n_2423),
.B(n_368),
.C(n_369),
.Y(n_2478)
);

OAI211xp5_ASAP7_75t_SL g2479 ( 
.A1(n_2431),
.A2(n_370),
.B(n_371),
.C(n_372),
.Y(n_2479)
);

OR2x2_ASAP7_75t_L g2480 ( 
.A(n_2441),
.B(n_371),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_L g2481 ( 
.A(n_2455),
.B(n_373),
.Y(n_2481)
);

NAND3xp33_ASAP7_75t_SL g2482 ( 
.A(n_2422),
.B(n_373),
.C(n_374),
.Y(n_2482)
);

NAND2x1p5_ASAP7_75t_L g2483 ( 
.A(n_2455),
.B(n_375),
.Y(n_2483)
);

NOR2xp67_ASAP7_75t_L g2484 ( 
.A(n_2456),
.B(n_376),
.Y(n_2484)
);

HB1xp67_ASAP7_75t_L g2485 ( 
.A(n_2443),
.Y(n_2485)
);

XNOR2xp5_ASAP7_75t_L g2486 ( 
.A(n_2453),
.B(n_377),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2417),
.Y(n_2487)
);

NAND4xp75_ASAP7_75t_L g2488 ( 
.A(n_2437),
.B(n_377),
.C(n_378),
.D(n_379),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2435),
.Y(n_2489)
);

NAND3xp33_ASAP7_75t_L g2490 ( 
.A(n_2433),
.B(n_379),
.C(n_380),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2416),
.Y(n_2491)
);

NAND2xp33_ASAP7_75t_R g2492 ( 
.A(n_2448),
.B(n_2457),
.Y(n_2492)
);

NAND3x1_ASAP7_75t_L g2493 ( 
.A(n_2428),
.B(n_381),
.C(n_382),
.Y(n_2493)
);

AOI22xp33_ASAP7_75t_SL g2494 ( 
.A1(n_2436),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_2494)
);

O2A1O1Ixp33_ASAP7_75t_L g2495 ( 
.A1(n_2432),
.A2(n_383),
.B(n_384),
.C(n_385),
.Y(n_2495)
);

AOI221x1_ASAP7_75t_L g2496 ( 
.A1(n_2425),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.C(n_388),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_2440),
.Y(n_2497)
);

OR4x2_ASAP7_75t_L g2498 ( 
.A(n_2454),
.B(n_386),
.C(n_387),
.D(n_388),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2459),
.Y(n_2499)
);

OR2x2_ASAP7_75t_L g2500 ( 
.A(n_2449),
.B(n_2452),
.Y(n_2500)
);

AND2x4_ASAP7_75t_L g2501 ( 
.A(n_2447),
.B(n_389),
.Y(n_2501)
);

NAND3xp33_ASAP7_75t_L g2502 ( 
.A(n_2458),
.B(n_389),
.C(n_390),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_2438),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2460),
.Y(n_2504)
);

NAND2xp33_ASAP7_75t_SL g2505 ( 
.A(n_2462),
.B(n_2444),
.Y(n_2505)
);

NAND3xp33_ASAP7_75t_L g2506 ( 
.A(n_2465),
.B(n_2430),
.C(n_2446),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2484),
.B(n_2445),
.Y(n_2507)
);

NAND2xp33_ASAP7_75t_SL g2508 ( 
.A(n_2500),
.B(n_391),
.Y(n_2508)
);

NOR2xp33_ASAP7_75t_R g2509 ( 
.A(n_2492),
.B(n_391),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_R g2510 ( 
.A(n_2471),
.B(n_392),
.Y(n_2510)
);

NOR2xp33_ASAP7_75t_R g2511 ( 
.A(n_2482),
.B(n_392),
.Y(n_2511)
);

NAND3xp33_ASAP7_75t_L g2512 ( 
.A(n_2487),
.B(n_393),
.C(n_394),
.Y(n_2512)
);

NAND2xp33_ASAP7_75t_SL g2513 ( 
.A(n_2486),
.B(n_393),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2463),
.B(n_394),
.Y(n_2514)
);

XOR2xp5_ASAP7_75t_L g2515 ( 
.A(n_2503),
.B(n_395),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2485),
.B(n_396),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_R g2517 ( 
.A(n_2497),
.B(n_396),
.Y(n_2517)
);

NOR3xp33_ASAP7_75t_SL g2518 ( 
.A(n_2491),
.B(n_2470),
.C(n_2489),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_SL g2519 ( 
.A(n_2463),
.B(n_397),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_R g2520 ( 
.A(n_2499),
.B(n_398),
.Y(n_2520)
);

NAND2xp33_ASAP7_75t_SL g2521 ( 
.A(n_2467),
.B(n_398),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2473),
.B(n_2483),
.Y(n_2522)
);

NAND2xp33_ASAP7_75t_SL g2523 ( 
.A(n_2467),
.B(n_399),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2481),
.B(n_400),
.Y(n_2524)
);

XOR2x2_ASAP7_75t_L g2525 ( 
.A(n_2493),
.B(n_400),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_SL g2526 ( 
.A(n_2501),
.B(n_401),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2501),
.B(n_402),
.Y(n_2527)
);

OAI21xp33_ASAP7_75t_L g2528 ( 
.A1(n_2504),
.A2(n_403),
.B(n_404),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_R g2529 ( 
.A(n_2468),
.B(n_404),
.Y(n_2529)
);

NAND3xp33_ASAP7_75t_SL g2530 ( 
.A(n_2480),
.B(n_405),
.C(n_406),
.Y(n_2530)
);

NAND2xp33_ASAP7_75t_SL g2531 ( 
.A(n_2466),
.B(n_405),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_2479),
.B(n_406),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_SL g2533 ( 
.A(n_2494),
.B(n_407),
.Y(n_2533)
);

NAND2xp33_ASAP7_75t_SL g2534 ( 
.A(n_2498),
.B(n_407),
.Y(n_2534)
);

XNOR2xp5_ASAP7_75t_L g2535 ( 
.A(n_2477),
.B(n_2488),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_SL g2536 ( 
.A(n_2472),
.B(n_408),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_R g2537 ( 
.A(n_2476),
.B(n_408),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2475),
.B(n_409),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2478),
.B(n_410),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_R g2540 ( 
.A(n_2495),
.B(n_410),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2525),
.Y(n_2541)
);

HB1xp67_ASAP7_75t_L g2542 ( 
.A(n_2509),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2507),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2534),
.Y(n_2544)
);

AOI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2518),
.A2(n_2490),
.B1(n_2502),
.B2(n_2474),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2527),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2515),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2522),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2535),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2526),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2514),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2521),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2519),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2524),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2523),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2516),
.Y(n_2556)
);

INVxp67_ASAP7_75t_L g2557 ( 
.A(n_2513),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2506),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2508),
.Y(n_2559)
);

AO22x2_ASAP7_75t_L g2560 ( 
.A1(n_2530),
.A2(n_2539),
.B1(n_2538),
.B2(n_2536),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2532),
.Y(n_2561)
);

OAI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2558),
.A2(n_2549),
.B1(n_2548),
.B2(n_2541),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2542),
.Y(n_2563)
);

AOI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2544),
.A2(n_2505),
.B1(n_2528),
.B2(n_2531),
.Y(n_2564)
);

OAI22xp5_ASAP7_75t_L g2565 ( 
.A1(n_2541),
.A2(n_2512),
.B1(n_2533),
.B2(n_2469),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2552),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2560),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2555),
.Y(n_2568)
);

AOI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2543),
.A2(n_2537),
.B1(n_2510),
.B2(n_2520),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2560),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2559),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2546),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2554),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2550),
.Y(n_2574)
);

AO22x2_ASAP7_75t_L g2575 ( 
.A1(n_2551),
.A2(n_2496),
.B1(n_2517),
.B2(n_2529),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2553),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2547),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2557),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2556),
.Y(n_2579)
);

AND3x1_ASAP7_75t_L g2580 ( 
.A(n_2545),
.B(n_2511),
.C(n_2540),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2561),
.Y(n_2581)
);

OAI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_2570),
.A2(n_2464),
.B1(n_412),
.B2(n_413),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2575),
.B(n_2111),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2575),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2566),
.Y(n_2585)
);

AND2x2_ASAP7_75t_SL g2586 ( 
.A(n_2580),
.B(n_411),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2567),
.B(n_411),
.Y(n_2587)
);

OR4x1_ASAP7_75t_L g2588 ( 
.A(n_2578),
.B(n_412),
.C(n_413),
.D(n_414),
.Y(n_2588)
);

AOI21xp5_ASAP7_75t_L g2589 ( 
.A1(n_2562),
.A2(n_414),
.B(n_415),
.Y(n_2589)
);

INVx3_ASAP7_75t_L g2590 ( 
.A(n_2573),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2569),
.Y(n_2591)
);

HB1xp67_ASAP7_75t_L g2592 ( 
.A(n_2574),
.Y(n_2592)
);

OA21x2_ASAP7_75t_L g2593 ( 
.A1(n_2568),
.A2(n_415),
.B(n_416),
.Y(n_2593)
);

OR4x1_ASAP7_75t_L g2594 ( 
.A(n_2563),
.B(n_417),
.C(n_418),
.D(n_419),
.Y(n_2594)
);

OAI22xp5_ASAP7_75t_SL g2595 ( 
.A1(n_2585),
.A2(n_2576),
.B1(n_2572),
.B2(n_2579),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2592),
.Y(n_2596)
);

AO22x2_ASAP7_75t_L g2597 ( 
.A1(n_2584),
.A2(n_2571),
.B1(n_2577),
.B2(n_2581),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2590),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2586),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2596),
.Y(n_2600)
);

BUFx2_ASAP7_75t_L g2601 ( 
.A(n_2597),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2598),
.A2(n_2564),
.B1(n_2591),
.B2(n_2587),
.Y(n_2602)
);

NAND3xp33_ASAP7_75t_L g2603 ( 
.A(n_2599),
.B(n_2565),
.C(n_2589),
.Y(n_2603)
);

AOI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2601),
.A2(n_2595),
.B1(n_2593),
.B2(n_2582),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2600),
.Y(n_2605)
);

OAI21x1_ASAP7_75t_L g2606 ( 
.A1(n_2602),
.A2(n_2583),
.B(n_2594),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2605),
.A2(n_2603),
.B(n_2588),
.Y(n_2607)
);

XNOR2xp5_ASAP7_75t_L g2608 ( 
.A(n_2604),
.B(n_418),
.Y(n_2608)
);

O2A1O1Ixp33_ASAP7_75t_L g2609 ( 
.A1(n_2606),
.A2(n_420),
.B(n_421),
.C(n_422),
.Y(n_2609)
);

OAI22xp5_ASAP7_75t_L g2610 ( 
.A1(n_2605),
.A2(n_420),
.B1(n_423),
.B2(n_424),
.Y(n_2610)
);

NAND3xp33_ASAP7_75t_L g2611 ( 
.A(n_2607),
.B(n_423),
.C(n_425),
.Y(n_2611)
);

NAND3xp33_ASAP7_75t_L g2612 ( 
.A(n_2608),
.B(n_425),
.C(n_426),
.Y(n_2612)
);

NAND3xp33_ASAP7_75t_L g2613 ( 
.A(n_2609),
.B(n_426),
.C(n_427),
.Y(n_2613)
);

OAI21xp5_ASAP7_75t_L g2614 ( 
.A1(n_2612),
.A2(n_2610),
.B(n_428),
.Y(n_2614)
);

OAI21xp5_ASAP7_75t_L g2615 ( 
.A1(n_2613),
.A2(n_427),
.B(n_428),
.Y(n_2615)
);

OAI211xp5_ASAP7_75t_L g2616 ( 
.A1(n_2615),
.A2(n_2611),
.B(n_430),
.C(n_431),
.Y(n_2616)
);

OR2x6_ASAP7_75t_L g2617 ( 
.A(n_2616),
.B(n_2614),
.Y(n_2617)
);

AOI21xp5_ASAP7_75t_L g2618 ( 
.A1(n_2617),
.A2(n_429),
.B(n_432),
.Y(n_2618)
);

AOI211xp5_ASAP7_75t_L g2619 ( 
.A1(n_2618),
.A2(n_433),
.B(n_434),
.C(n_435),
.Y(n_2619)
);


endmodule