module fake_jpeg_13447_n_211 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_211);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_211;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_5),
.B(n_6),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_21),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_48),
.B(n_55),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_21),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_26),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_60),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_12),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_11),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_57),
.B(n_58),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_11),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_59),
.B(n_64),
.Y(n_114)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_2),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_69),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_2),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_70),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_2),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_73),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_74),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_3),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_27),
.B(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_76),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_30),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_35),
.B1(n_72),
.B2(n_42),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_77),
.A2(n_91),
.B1(n_113),
.B2(n_81),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_34),
.B1(n_16),
.B2(n_38),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_79),
.A2(n_90),
.B1(n_95),
.B2(n_102),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_40),
.A2(n_16),
.B(n_17),
.C(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_84),
.B(n_110),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_28),
.B1(n_37),
.B2(n_32),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_88),
.A2(n_110),
.B1(n_81),
.B2(n_108),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_46),
.A2(n_28),
.B1(n_37),
.B2(n_32),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_27),
.B1(n_31),
.B2(n_38),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_53),
.B1(n_76),
.B2(n_65),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_31),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_54),
.A2(n_4),
.B1(n_7),
.B2(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_56),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_123),
.Y(n_143)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_40),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_83),
.B(n_89),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_137),
.B(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_142),
.Y(n_153)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_136),
.B1(n_138),
.B2(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_90),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_141),
.Y(n_158)
);

OA22x2_ASAP7_75t_SL g135 ( 
.A1(n_79),
.A2(n_101),
.B1(n_111),
.B2(n_110),
.Y(n_135)
);

AO22x1_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_85),
.B1(n_106),
.B2(n_86),
.Y(n_159)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_109),
.B1(n_105),
.B2(n_114),
.Y(n_156)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_123),
.B(n_92),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_157),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_156),
.A2(n_160),
.B1(n_121),
.B2(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_144),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_105),
.B1(n_109),
.B2(n_86),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_169),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_SL g163 ( 
.A(n_143),
.B(n_119),
.C(n_115),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_164),
.C(n_167),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_124),
.C(n_118),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_165),
.A2(n_157),
.B(n_161),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

XOR2x2_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_139),
.B1(n_135),
.B2(n_136),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_171),
.B1(n_150),
.B2(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_170),
.B(n_174),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_160),
.B1(n_158),
.B2(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_100),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_179),
.B(n_183),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_178),
.A2(n_182),
.B1(n_170),
.B2(n_151),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_167),
.A2(n_159),
.B(n_146),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_158),
.B1(n_159),
.B2(n_127),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_159),
.B(n_149),
.Y(n_183)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_146),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_166),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_164),
.C(n_163),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_187),
.C(n_191),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_161),
.C(n_171),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_193),
.B1(n_182),
.B2(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_149),
.C(n_155),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_145),
.C(n_117),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_175),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_185),
.A2(n_151),
.B1(n_120),
.B2(n_126),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_180),
.B1(n_185),
.B2(n_176),
.Y(n_197)
);

AOI31xp67_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_184),
.A3(n_179),
.B(n_183),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_199),
.A2(n_198),
.B1(n_190),
.B2(n_196),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_196),
.C(n_194),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_204),
.Y(n_206)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_180),
.C(n_176),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_206),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_208),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_151),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_145),
.B(n_85),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_132),
.Y(n_211)
);


endmodule