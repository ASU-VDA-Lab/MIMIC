module fake_jpeg_2718_n_650 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_650);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_650;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_58),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_59),
.B(n_82),
.Y(n_137)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_62),
.Y(n_151)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_65),
.Y(n_164)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_66),
.Y(n_206)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_67),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_68),
.Y(n_227)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_69),
.Y(n_172)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_70),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_72),
.Y(n_168)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_74),
.Y(n_183)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_75),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_20),
.B(n_10),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_77),
.B(n_81),
.Y(n_163)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_78),
.Y(n_174)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_10),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_119),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_9),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_85),
.B(n_87),
.Y(n_192)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_26),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_26),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_88),
.B(n_91),
.Y(n_209)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_32),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_89),
.Y(n_134)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_22),
.B(n_9),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_92),
.Y(n_179)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_93),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_94),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_96),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_9),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_97),
.B(n_98),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_23),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

BUFx16f_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_9),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_105),
.B(n_111),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_107),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_110),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_37),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_112),
.Y(n_154)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_115),
.Y(n_166)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_118),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_48),
.B(n_11),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_37),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_120),
.B(n_38),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_49),
.B(n_8),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_51),
.Y(n_150)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_125),
.Y(n_216)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_24),
.Y(n_126)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_127),
.Y(n_217)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_42),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_23),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_85),
.B(n_56),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_136),
.B(n_226),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_104),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_142),
.B(n_150),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_97),
.A2(n_51),
.B1(n_55),
.B2(n_54),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_143),
.A2(n_203),
.B(n_23),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_89),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_146),
.B(n_213),
.Y(n_231)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_162),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_105),
.B(n_56),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_167),
.B(n_184),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_70),
.B(n_52),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_169),
.B(n_199),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g170 ( 
.A(n_64),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g239 ( 
.A(n_170),
.Y(n_239)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_171),
.Y(n_258)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_61),
.Y(n_175)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_79),
.Y(n_176)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_60),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_185),
.Y(n_298)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_80),
.Y(n_188)
);

INVx3_ASAP7_75t_SL g295 ( 
.A(n_188),
.Y(n_295)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_108),
.Y(n_190)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_190),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_127),
.A2(n_39),
.B1(n_52),
.B2(n_54),
.Y(n_194)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_194),
.A2(n_200),
.B1(n_221),
.B2(n_24),
.Y(n_241)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_195),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_130),
.B(n_55),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_106),
.A2(n_39),
.B1(n_43),
.B2(n_33),
.Y(n_200)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_201),
.Y(n_308)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_96),
.Y(n_202)
);

CKINVDCx9p33_ASAP7_75t_R g242 ( 
.A(n_202),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_100),
.A2(n_38),
.B(n_33),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_212),
.Y(n_259)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_66),
.B(n_14),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_69),
.Y(n_240)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_99),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_67),
.A2(n_23),
.B1(n_41),
.B2(n_24),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_68),
.B(n_13),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_222),
.B(n_2),
.Y(n_268)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_101),
.Y(n_224)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_224),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_122),
.B(n_13),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_121),
.B1(n_114),
.B2(n_110),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_228),
.A2(n_152),
.B1(n_206),
.B2(n_187),
.Y(n_327)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_243),
.Y(n_312)
);

NOR2x1_ASAP7_75t_R g337 ( 
.A(n_232),
.B(n_147),
.Y(n_337)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_233),
.Y(n_315)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_148),
.Y(n_234)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_234),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_236),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_238),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_240),
.B(n_251),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_241),
.A2(n_299),
.B1(n_300),
.B2(n_303),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_173),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_209),
.A2(n_95),
.B1(n_94),
.B2(n_92),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_244),
.A2(n_276),
.B1(n_280),
.B2(n_215),
.Y(n_318)
);

CKINVDCx12_ASAP7_75t_R g245 ( 
.A(n_157),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_245),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_211),
.A2(n_84),
.B1(n_76),
.B2(n_71),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_246),
.Y(n_340)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_247),
.Y(n_319)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_250),
.B(n_256),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_141),
.B(n_12),
.Y(n_251)
);

AO22x1_ASAP7_75t_L g252 ( 
.A1(n_192),
.A2(n_39),
.B1(n_45),
.B2(n_41),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_252),
.B(n_296),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_167),
.B(n_0),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_254),
.Y(n_341)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_148),
.Y(n_255)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_255),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_45),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_257),
.B(n_272),
.Y(n_338)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_137),
.B(n_45),
.C(n_41),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_261),
.B(n_269),
.C(n_278),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_216),
.A2(n_221),
.B1(n_166),
.B2(n_208),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_263),
.Y(n_339)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_144),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_219),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_266),
.A2(n_284),
.B1(n_160),
.B2(n_187),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_268),
.B(n_271),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_182),
.B(n_2),
.C(n_4),
.Y(n_269)
);

CKINVDCx12_ASAP7_75t_R g270 ( 
.A(n_157),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_270),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_163),
.B(n_5),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_136),
.B(n_5),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_216),
.A2(n_221),
.B1(n_166),
.B2(n_225),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_273),
.Y(n_342)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_193),
.Y(n_275)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_275),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_163),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_183),
.Y(n_277)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_277),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_6),
.C(n_8),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_173),
.Y(n_279)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_194),
.A2(n_6),
.B1(n_12),
.B2(n_15),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_177),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_281),
.B(n_289),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_140),
.B(n_6),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_292),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_156),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_284)
);

HAxp5_ASAP7_75t_SL g285 ( 
.A(n_134),
.B(n_15),
.CON(n_285),
.SN(n_285)
);

OR2x2_ASAP7_75t_SL g335 ( 
.A(n_285),
.B(n_132),
.Y(n_335)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_198),
.Y(n_287)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_287),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_288),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_154),
.B(n_15),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_154),
.Y(n_290)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_290),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_153),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_291),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_161),
.B(n_16),
.Y(n_292)
);

INVx6_ASAP7_75t_L g293 ( 
.A(n_218),
.Y(n_293)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_215),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_294),
.Y(n_356)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_172),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_153),
.A2(n_17),
.B1(n_18),
.B2(n_131),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_159),
.A2(n_177),
.B1(n_210),
.B2(n_189),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_164),
.B(n_178),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_302),
.Y(n_336)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_172),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_138),
.A2(n_17),
.B1(n_196),
.B2(n_200),
.Y(n_303)
);

BUFx12_ASAP7_75t_L g304 ( 
.A(n_135),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_304),
.B(n_306),
.Y(n_371)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_170),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_309),
.Y(n_347)
);

CKINVDCx12_ASAP7_75t_R g306 ( 
.A(n_135),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_168),
.B(n_186),
.Y(n_309)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_152),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_310),
.B(n_311),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_149),
.B(n_151),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_267),
.B(n_191),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_316),
.B(n_361),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_317),
.B(n_325),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_318),
.A2(n_328),
.B1(n_350),
.B2(n_351),
.Y(n_391)
);

AND2x4_ASAP7_75t_SL g320 ( 
.A(n_244),
.B(n_280),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_320),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_252),
.A2(n_207),
.B1(n_204),
.B2(n_206),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_327),
.A2(n_238),
.B1(n_279),
.B2(n_298),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_241),
.A2(n_181),
.B1(n_179),
.B2(n_160),
.Y(n_328)
);

AOI32xp33_ASAP7_75t_L g329 ( 
.A1(n_261),
.A2(n_135),
.A3(n_179),
.B1(n_181),
.B2(n_139),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_329),
.A2(n_349),
.B(n_346),
.C(n_339),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_L g332 ( 
.A1(n_246),
.A2(n_139),
.B1(n_155),
.B2(n_147),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_332),
.A2(n_344),
.B1(n_346),
.B2(n_328),
.Y(n_406)
);

OR2x2_ASAP7_75t_SL g409 ( 
.A(n_335),
.B(n_337),
.Y(n_409)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_284),
.A2(n_147),
.B1(n_212),
.B2(n_155),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_241),
.A2(n_212),
.B1(n_133),
.B2(n_145),
.Y(n_346)
);

AOI32xp33_ASAP7_75t_L g349 ( 
.A1(n_231),
.A2(n_132),
.A3(n_133),
.B1(n_145),
.B2(n_307),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_241),
.A2(n_132),
.B1(n_133),
.B2(n_145),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_242),
.A2(n_274),
.B1(n_302),
.B2(n_296),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_254),
.B(n_264),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_354),
.B(n_369),
.C(n_297),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_242),
.A2(n_277),
.B1(n_265),
.B2(n_258),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_254),
.B(n_276),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_269),
.B(n_278),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_341),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_233),
.A2(n_247),
.B1(n_258),
.B2(n_297),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_367),
.A2(n_293),
.B1(n_234),
.B2(n_255),
.Y(n_393)
);

MAJx2_ASAP7_75t_L g369 ( 
.A(n_283),
.B(n_266),
.C(n_260),
.Y(n_369)
);

MAJx2_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_323),
.C(n_363),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_372),
.B(n_373),
.C(n_395),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_287),
.C(n_262),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_360),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_375),
.B(n_377),
.Y(n_424)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_357),
.Y(n_376)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_360),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_365),
.Y(n_378)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_378),
.Y(n_422)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_379),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_347),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_380),
.B(n_388),
.Y(n_445)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_321),
.B(n_295),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_383),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_384),
.B(n_389),
.Y(n_447)
);

BUFx12_ASAP7_75t_L g385 ( 
.A(n_331),
.Y(n_385)
);

BUFx4f_ASAP7_75t_L g428 ( 
.A(n_385),
.Y(n_428)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_386),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_387),
.B(n_393),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_285),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_322),
.B(n_298),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_390),
.B(n_407),
.Y(n_426)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_392),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_330),
.A2(n_308),
.B(n_237),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_394),
.A2(n_345),
.B(n_319),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_295),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_330),
.A2(n_239),
.B(n_235),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_396),
.B(n_401),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_358),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_408),
.Y(n_423)
);

BUFx2_ASAP7_75t_SL g398 ( 
.A(n_333),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_398),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g401 ( 
.A(n_330),
.B(n_239),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_402),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_313),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_403),
.B(n_404),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_312),
.Y(n_404)
);

INVx8_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_405),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_406),
.A2(n_418),
.B1(n_340),
.B2(n_339),
.Y(n_427)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_349),
.B(n_305),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_324),
.B(n_286),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g410 ( 
.A(n_314),
.B(n_275),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_410),
.B(n_411),
.Y(n_432)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_315),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_341),
.B(n_249),
.C(n_235),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_417),
.C(n_335),
.Y(n_438)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_413),
.B(n_414),
.Y(n_440)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_326),
.Y(n_414)
);

BUFx12_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_416),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_336),
.B(n_310),
.Y(n_416)
);

MAJx2_ASAP7_75t_L g417 ( 
.A(n_321),
.B(n_308),
.C(n_236),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_399),
.A2(n_318),
.B1(n_340),
.B2(n_342),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_419),
.A2(n_431),
.B1(n_396),
.B2(n_389),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_427),
.A2(n_417),
.B1(n_412),
.B2(n_416),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_406),
.A2(n_342),
.B1(n_352),
.B2(n_320),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_384),
.A2(n_320),
.B1(n_325),
.B2(n_329),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_434),
.A2(n_436),
.B1(n_437),
.B2(n_442),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_382),
.A2(n_320),
.B1(n_314),
.B2(n_364),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_382),
.A2(n_364),
.B1(n_368),
.B2(n_317),
.Y(n_437)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_425),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_387),
.A2(n_368),
.B(n_371),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_439),
.A2(n_334),
.B(n_230),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_382),
.A2(n_338),
.B1(n_369),
.B2(n_356),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_374),
.B(n_369),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_443),
.B(n_452),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_394),
.A2(n_312),
.B(n_333),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_449),
.A2(n_455),
.B(n_458),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_391),
.A2(n_370),
.B1(n_343),
.B2(n_353),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_450),
.A2(n_453),
.B1(n_378),
.B2(n_392),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_374),
.B(n_322),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_397),
.A2(n_370),
.B1(n_343),
.B2(n_353),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_395),
.B(n_338),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_401),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_372),
.B(n_362),
.C(n_345),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_403),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_408),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_459),
.B(n_469),
.Y(n_499)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_460),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_425),
.B(n_373),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_461),
.B(n_489),
.C(n_447),
.Y(n_500)
);

CKINVDCx11_ASAP7_75t_R g462 ( 
.A(n_436),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_462),
.B(n_475),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_463),
.A2(n_467),
.B1(n_471),
.B2(n_476),
.Y(n_511)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_422),
.Y(n_464)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_464),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_468),
.B(n_490),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_362),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_470),
.B(n_487),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_431),
.A2(n_407),
.B1(n_396),
.B2(n_418),
.Y(n_471)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_472),
.Y(n_505)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_446),
.Y(n_473)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_473),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_452),
.B(n_423),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_474),
.B(n_481),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_426),
.B(n_410),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_434),
.A2(n_388),
.B1(n_409),
.B2(n_400),
.Y(n_476)
);

AND2x2_ASAP7_75t_SL g478 ( 
.A(n_458),
.B(n_409),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_478),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_479),
.B(n_435),
.Y(n_515)
);

BUFx12_ASAP7_75t_L g480 ( 
.A(n_428),
.Y(n_480)
);

INVx13_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_423),
.B(n_411),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_440),
.Y(n_482)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_482),
.B(n_485),
.C(n_492),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_455),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_483),
.B(n_486),
.Y(n_526)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_446),
.Y(n_484)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_484),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_440),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_435),
.B(n_386),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_426),
.A2(n_400),
.B1(n_405),
.B2(n_379),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_451),
.A2(n_359),
.B1(n_366),
.B2(n_294),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_488),
.B(n_450),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_447),
.B(n_415),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_445),
.B(n_415),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_SL g491 ( 
.A1(n_419),
.A2(n_334),
.B1(n_248),
.B2(n_359),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_491),
.A2(n_451),
.B(n_427),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_439),
.A2(n_449),
.B(n_451),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_493),
.A2(n_449),
.B(n_421),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_429),
.Y(n_494)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_494),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_454),
.B(n_442),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_495),
.B(n_470),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_500),
.B(n_506),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_486),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_504),
.B(n_513),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_457),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_466),
.B(n_429),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_509),
.B(n_519),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_472),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_461),
.B(n_438),
.C(n_443),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_514),
.B(n_522),
.C(n_524),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_515),
.B(n_492),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_516),
.A2(n_487),
.B(n_488),
.Y(n_548)
);

OAI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_518),
.A2(n_480),
.B1(n_248),
.B2(n_288),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_466),
.B(n_453),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_521),
.B(n_527),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_479),
.B(n_432),
.C(n_421),
.Y(n_522)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_523),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_478),
.B(n_432),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_468),
.B(n_441),
.C(n_437),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_525),
.B(n_528),
.C(n_530),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_482),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_430),
.Y(n_528)
);

OA21x2_ASAP7_75t_L g529 ( 
.A1(n_465),
.A2(n_430),
.B(n_420),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_529),
.B(n_428),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_468),
.B(n_441),
.C(n_420),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_505),
.A2(n_467),
.B1(n_471),
.B2(n_462),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_531),
.A2(n_551),
.B1(n_518),
.B2(n_512),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_501),
.A2(n_485),
.B1(n_465),
.B2(n_476),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_535),
.A2(n_543),
.B1(n_547),
.B2(n_549),
.Y(n_561)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_498),
.Y(n_536)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_536),
.Y(n_564)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_498),
.Y(n_538)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_538),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_539),
.B(n_555),
.Y(n_568)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_503),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_540),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_506),
.B(n_468),
.C(n_477),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_542),
.B(n_552),
.C(n_530),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_513),
.A2(n_483),
.B1(n_475),
.B2(n_477),
.Y(n_543)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_517),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_545),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_501),
.A2(n_493),
.B1(n_490),
.B2(n_460),
.Y(n_547)
);

A2O1A1Ixp33_ASAP7_75t_SL g567 ( 
.A1(n_548),
.A2(n_554),
.B(n_557),
.C(n_549),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_505),
.A2(n_468),
.B1(n_464),
.B2(n_473),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_499),
.Y(n_550)
);

CKINVDCx14_ASAP7_75t_R g563 ( 
.A(n_550),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_502),
.A2(n_484),
.B1(n_468),
.B2(n_428),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_514),
.B(n_444),
.C(n_448),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_496),
.A2(n_428),
.B1(n_456),
.B2(n_444),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_553),
.A2(n_526),
.B1(n_510),
.B2(n_503),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_512),
.A2(n_448),
.B(n_456),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g556 ( 
.A(n_500),
.B(n_385),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_556),
.B(n_558),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_507),
.A2(n_516),
.B(n_520),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_559),
.B(n_567),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_560),
.B(n_570),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_552),
.B(n_525),
.C(n_515),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_562),
.B(n_565),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_550),
.A2(n_502),
.B1(n_496),
.B2(n_523),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_541),
.B(n_542),
.C(n_537),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_569),
.B(n_571),
.C(n_580),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_537),
.B(n_522),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_541),
.B(n_524),
.C(n_511),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_556),
.B(n_511),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_573),
.B(n_575),
.Y(n_597)
);

NOR3xp33_ASAP7_75t_SL g574 ( 
.A(n_546),
.B(n_499),
.C(n_517),
.Y(n_574)
);

CKINVDCx14_ASAP7_75t_R g589 ( 
.A(n_574),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_534),
.B(n_528),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_534),
.B(n_529),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_576),
.B(n_578),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_539),
.B(n_529),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_558),
.B(n_526),
.C(n_504),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_581),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_561),
.A2(n_531),
.B1(n_548),
.B2(n_532),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_585),
.A2(n_596),
.B1(n_599),
.B2(n_259),
.Y(n_613)
);

BUFx24_ASAP7_75t_SL g586 ( 
.A(n_563),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_586),
.B(n_577),
.Y(n_604)
);

AO221x1_ASAP7_75t_L g587 ( 
.A1(n_567),
.A2(n_546),
.B1(n_544),
.B2(n_533),
.C(n_532),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_587),
.B(n_588),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_560),
.B(n_543),
.C(n_553),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_569),
.B(n_555),
.C(n_533),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_591),
.B(n_592),
.C(n_594),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_562),
.B(n_545),
.C(n_554),
.Y(n_592)
);

INVx13_ASAP7_75t_L g593 ( 
.A(n_566),
.Y(n_593)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_593),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_540),
.C(n_538),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g595 ( 
.A1(n_567),
.A2(n_580),
.B(n_572),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_595),
.B(n_385),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_567),
.A2(n_544),
.B(n_536),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g599 ( 
.A1(n_573),
.A2(n_510),
.B1(n_508),
.B2(n_497),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_590),
.A2(n_572),
.B1(n_577),
.B2(n_568),
.Y(n_602)
);

XNOR2x1_ASAP7_75t_L g626 ( 
.A(n_602),
.B(n_612),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g603 ( 
.A(n_597),
.B(n_571),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_603),
.B(n_607),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_604),
.B(n_606),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_583),
.B(n_568),
.C(n_579),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_597),
.B(n_564),
.Y(n_607)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_591),
.B(n_574),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_609),
.B(n_616),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_589),
.A2(n_508),
.B1(n_497),
.B2(n_480),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_610),
.B(n_611),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_584),
.A2(n_480),
.B1(n_366),
.B2(n_319),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_613),
.A2(n_596),
.B(n_595),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_583),
.B(n_249),
.C(n_253),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_614),
.B(n_615),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_253),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_582),
.B(n_259),
.Y(n_616)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_617),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_582),
.C(n_606),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_620),
.B(n_588),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_609),
.A2(n_598),
.B(n_605),
.Y(n_621)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_621),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_601),
.A2(n_590),
.B(n_587),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_623),
.B(n_627),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g627 ( 
.A(n_607),
.B(n_592),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_623),
.A2(n_584),
.B1(n_602),
.B2(n_608),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_628),
.A2(n_633),
.B1(n_585),
.B2(n_599),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_619),
.B(n_616),
.Y(n_629)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_629),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_620),
.B(n_603),
.Y(n_631)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_631),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_627),
.B(n_584),
.Y(n_634)
);

AOI31xp67_ASAP7_75t_L g638 ( 
.A1(n_634),
.A2(n_618),
.A3(n_622),
.B(n_626),
.Y(n_638)
);

AOI31xp67_ASAP7_75t_SL g636 ( 
.A1(n_632),
.A2(n_617),
.A3(n_614),
.B(n_622),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_636),
.B(n_638),
.C(n_630),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_637),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_641),
.A2(n_642),
.B(n_635),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_640),
.B(n_635),
.C(n_628),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_644),
.B(n_645),
.C(n_625),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_643),
.B(n_639),
.C(n_618),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_624),
.C(n_626),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_647),
.A2(n_600),
.B(n_612),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_648),
.A2(n_600),
.B1(n_593),
.B2(n_230),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_649),
.A2(n_304),
.B(n_375),
.Y(n_650)
);


endmodule