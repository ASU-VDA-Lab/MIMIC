module fake_jpeg_28030_n_178 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_36),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_SL g40 ( 
.A1(n_17),
.A2(n_1),
.B(n_2),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_2),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_48),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_54),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_25),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_18),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_18),
.Y(n_57)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_70),
.C(n_76),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_20),
.Y(n_64)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_77),
.C(n_47),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_74),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_16),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_10),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_10),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_83),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_45),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_95),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_57),
.B1(n_45),
.B2(n_42),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_18),
.B(n_33),
.C(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_70),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_77),
.A3(n_80),
.B1(n_21),
.B2(n_19),
.C1(n_15),
.C2(n_8),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_28),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_21),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_62),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_81),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_104),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_76),
.C(n_61),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_83),
.C(n_84),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_37),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_109),
.B(n_114),
.Y(n_124)
);

AOI322xp5_ASAP7_75t_SL g121 ( 
.A1(n_108),
.A2(n_97),
.A3(n_14),
.B1(n_9),
.B2(n_12),
.C1(n_13),
.C2(n_15),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_78),
.B(n_75),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_111),
.B(n_94),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_56),
.B(n_66),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_56),
.B(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_131),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_132),
.C(n_3),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_123),
.C(n_107),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_128),
.B(n_110),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_130),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_91),
.B(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_98),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_90),
.Y(n_131)
);

NOR3xp33_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_19),
.C(n_87),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_106),
.B1(n_109),
.B2(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_102),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_142),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_118),
.Y(n_142)
);

AOI321xp33_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_128),
.A3(n_122),
.B1(n_131),
.B2(n_123),
.C(n_110),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_110),
.B(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_117),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_146),
.A2(n_126),
.B(n_124),
.Y(n_148)
);

OAI21x1_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_150),
.B(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_132),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_155),
.C(n_135),
.Y(n_158)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_90),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_3),
.C(n_4),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_155),
.B(n_137),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_141),
.B1(n_145),
.B2(n_100),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_157),
.A2(n_158),
.B(n_30),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_161),
.Y(n_168)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_160),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_163),
.A2(n_165),
.B(n_167),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_143),
.C(n_136),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_166),
.C(n_27),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_137),
.C(n_30),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_170),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_23),
.B1(n_27),
.B2(n_5),
.C(n_3),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_4),
.A3(n_5),
.B1(n_46),
.B2(n_49),
.C1(n_43),
.C2(n_44),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_4),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_174),
.C(n_53),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_46),
.B(n_43),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_177),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_175),
.Y(n_177)
);


endmodule