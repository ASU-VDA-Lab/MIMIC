module fake_jpeg_18113_n_212 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx11_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_26),
.Y(n_37)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_29),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_17),
.B1(n_12),
.B2(n_24),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_40),
.B1(n_42),
.B2(n_28),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_17),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_32),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_24),
.B(n_18),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_12),
.B1(n_22),
.B2(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_25),
.B(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_29),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_51),
.B1(n_62),
.B2(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_63),
.B(n_39),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_27),
.B1(n_26),
.B2(n_30),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_12),
.B1(n_33),
.B2(n_13),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_38),
.B(n_45),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_30),
.B1(n_29),
.B2(n_32),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_67),
.B(n_71),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_32),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_78),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_40),
.B(n_41),
.C(n_37),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_75),
.B(n_76),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_41),
.B(n_36),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_43),
.B(n_45),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_38),
.B(n_42),
.C(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_62),
.B1(n_44),
.B2(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_57),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_21),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_50),
.C(n_60),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_97),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_96),
.B1(n_78),
.B2(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_73),
.B(n_35),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_63),
.B1(n_59),
.B2(n_58),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_60),
.C(n_55),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_99),
.A2(n_111),
.B1(n_84),
.B2(n_96),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_75),
.B(n_68),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_101),
.B(n_104),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_76),
.B1(n_87),
.B2(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_85),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_102),
.B(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_81),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_69),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_71),
.B(n_64),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_90),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_69),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_113),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_49),
.B1(n_53),
.B2(n_44),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_114),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_65),
.B1(n_66),
.B2(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_0),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_87),
.C(n_91),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_117),
.C(n_120),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_91),
.C(n_88),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_88),
.C(n_97),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_122),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_112),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_104),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_97),
.C(n_86),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_98),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_89),
.B1(n_114),
.B2(n_95),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_108),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_96),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_133),
.Y(n_136)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_130),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_135),
.A2(n_131),
.B1(n_133),
.B2(n_127),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_99),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_138),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_95),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_149),
.C(n_20),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_108),
.B(n_113),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_119),
.B(n_129),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_102),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_21),
.C(n_20),
.Y(n_162)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_145),
.B(n_146),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_92),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_98),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_157),
.B1(n_142),
.B2(n_35),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_127),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_120),
.B1(n_118),
.B2(n_125),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_1),
.C(n_2),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_123),
.B1(n_132),
.B2(n_77),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_159),
.A2(n_150),
.B1(n_149),
.B2(n_145),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_138),
.A2(n_66),
.B(n_2),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_161),
.A2(n_134),
.B(n_135),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_164),
.C(n_20),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_172),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_141),
.B1(n_150),
.B2(n_137),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_168),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_176),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_170),
.A2(n_155),
.B1(n_163),
.B2(n_161),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_170),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_16),
.C(n_14),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_175),
.C(n_2),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_16),
.C(n_14),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_157),
.B(n_159),
.Y(n_176)
);

OAI321xp33_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_160),
.A3(n_153),
.B1(n_152),
.B2(n_155),
.C(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_181),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_172),
.B1(n_4),
.B2(n_5),
.Y(n_194)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_16),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_173),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_165),
.B1(n_167),
.B2(n_171),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_188),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_182),
.C(n_181),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_192),
.C(n_194),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_174),
.Y(n_192)
);

NOR2xp67_ASAP7_75t_SL g196 ( 
.A(n_189),
.B(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_198),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_199),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_191),
.A2(n_3),
.B(n_4),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_187),
.A2(n_4),
.B(n_5),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_195),
.C(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_204),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_190),
.C(n_193),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_201),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_206),
.B(n_8),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_6),
.C(n_7),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_209),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_199),
.Y(n_210)
);

AOI321xp33_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C(n_206),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_8),
.C(n_9),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_11),
.Y(n_212)
);


endmodule