module real_aes_15448_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_23;
wire n_20;
wire n_18;
wire n_21;
wire n_10;
INVx2_ASAP7_75t_L g21 ( .A(n_0), .Y(n_21) );
OAI221xp5_ASAP7_75t_L g18 ( .A1(n_1), .A2(n_4), .B1(n_19), .B2(n_22), .C(n_25), .Y(n_18) );
INVx1_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_3), .Y(n_14) );
OAI21xp33_ASAP7_75t_L g13 ( .A1(n_5), .A2(n_14), .B(n_15), .Y(n_13) );
AOI321xp33_ASAP7_75t_L g9 ( .A1(n_6), .A2(n_7), .A3(n_10), .B1(n_12), .B2(n_13), .C(n_17), .Y(n_9) );
HB1xp67_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
CKINVDCx16_ASAP7_75t_R g16 ( .A(n_10), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_10), .B(n_18), .Y(n_17) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_12), .B(n_16), .Y(n_15) );
CKINVDCx16_ASAP7_75t_R g25 ( .A(n_12), .Y(n_25) );
INVx2_ASAP7_75t_SL g19 ( .A(n_20), .Y(n_19) );
INVx1_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
INVx2_ASAP7_75t_L g20 ( .A(n_21), .Y(n_20) );
INVx2_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
BUFx2_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
endmodule