module fake_jpeg_27753_n_189 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_12),
.B(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_28),
.Y(n_47)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_1),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_16),
.B1(n_32),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_52),
.B1(n_55),
.B2(n_19),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_16),
.B1(n_32),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_25),
.B1(n_18),
.B2(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_21),
.B1(n_23),
.B2(n_30),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_23),
.B1(n_19),
.B2(n_30),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_57),
.Y(n_87)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_29),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_17),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_74),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_35),
.B1(n_41),
.B2(n_23),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_72),
.B1(n_73),
.B2(n_79),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_29),
.B(n_26),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_47),
.B(n_20),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_23),
.B1(n_27),
.B2(n_20),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_19),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_77),
.Y(n_92)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

XNOR2x1_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_17),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_86),
.Y(n_97)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_18),
.C(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_78),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_105),
.B(n_68),
.Y(n_110)
);

OAI32xp33_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_20),
.A3(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_62),
.B(n_71),
.C(n_77),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_100),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_62),
.B(n_58),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_76),
.B(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_85),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_58),
.C(n_75),
.Y(n_125)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_111),
.B(n_115),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_79),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_91),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_73),
.B(n_68),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_120),
.B(n_124),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_68),
.B1(n_75),
.B2(n_77),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_104),
.B1(n_105),
.B2(n_90),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_81),
.B(n_67),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_127),
.C(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_67),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_67),
.C(n_75),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_90),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_136),
.B1(n_113),
.B2(n_2),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_97),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_116),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_140),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_89),
.C(n_98),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_101),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_94),
.B1(n_93),
.B2(n_103),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_118),
.B1(n_122),
.B2(n_126),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_94),
.B1(n_95),
.B2(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_95),
.C(n_88),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_143),
.C(n_123),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_103),
.C(n_107),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_115),
.A3(n_121),
.B1(n_114),
.B2(n_117),
.C1(n_111),
.C2(n_112),
.Y(n_147)
);

AOI322xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_140),
.A3(n_138),
.B1(n_142),
.B2(n_129),
.C1(n_15),
.C2(n_14),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_156),
.B1(n_139),
.B2(n_144),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_1),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_153),
.C(n_155),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_119),
.C(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_113),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_159),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_138),
.B1(n_135),
.B2(n_136),
.Y(n_159)
);

NOR4xp25_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_163),
.C(n_169),
.D(n_165),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_14),
.C(n_2),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_153),
.Y(n_170)
);

AOI31xp33_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_1),
.A3(n_3),
.B(n_4),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_151),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_3),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_4),
.B(n_5),
.Y(n_166)
);

AOI21x1_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_6),
.B(n_7),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

OAI31xp33_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_176),
.A3(n_8),
.B(n_10),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_172),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_175),
.A2(n_157),
.B(n_159),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_174),
.B(n_160),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_167),
.B1(n_158),
.B2(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_179),
.B(n_181),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_180),
.B(n_172),
.C(n_10),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_12),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_184),
.B(n_183),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_187),
.Y(n_189)
);


endmodule