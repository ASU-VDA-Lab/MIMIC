module fake_jpeg_30946_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_63),
.Y(n_65)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_0),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_48),
.B1(n_56),
.B2(n_51),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_46),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_79),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_53),
.B1(n_52),
.B2(n_56),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_36),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_47),
.Y(n_84)
);

OR2x2_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_5),
.Y(n_97)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_43),
.B1(n_37),
.B2(n_24),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_20),
.B1(n_35),
.B2(n_34),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_90),
.B(n_6),
.Y(n_98)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_91),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_30),
.B(n_31),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_12),
.B1(n_13),
.B2(n_17),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_18),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_112),
.Y(n_116)
);

XNOR2x1_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_102),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_114),
.Y(n_117)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_94),
.B(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_118),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_105),
.C(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_119),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_117),
.B(n_115),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_110),
.B(n_121),
.C(n_112),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_96),
.Y(n_127)
);


endmodule