module fake_jpeg_25612_n_273 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_13;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_29),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_22),
.B1(n_26),
.B2(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_22),
.B1(n_36),
.B2(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_50),
.B(n_19),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_27),
.B(n_30),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NAND2x1_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_56),
.B1(n_41),
.B2(n_38),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_46),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_67),
.Y(n_90)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_65),
.B1(n_59),
.B2(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_22),
.B1(n_38),
.B2(n_41),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_97),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_51),
.B(n_58),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_92),
.B(n_27),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_58),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_39),
.CI(n_33),
.CON(n_93),
.SN(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_37),
.B1(n_44),
.B2(n_47),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_105),
.B1(n_98),
.B2(n_102),
.Y(n_112)
);

OAI22x1_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_59),
.B1(n_52),
.B2(n_41),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_64),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_102),
.Y(n_123)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_68),
.B(n_83),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_124),
.B(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_120),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_83),
.B1(n_81),
.B2(n_70),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_115),
.B1(n_120),
.B2(n_107),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_117),
.B1(n_98),
.B2(n_102),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_84),
.B1(n_101),
.B2(n_73),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_74),
.B1(n_82),
.B2(n_37),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_39),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_71),
.B1(n_57),
.B2(n_60),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_35),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_121),
.C(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_78),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_33),
.C(n_38),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_35),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_111),
.B(n_119),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_135),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_125),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_131),
.B(n_137),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_133),
.Y(n_166)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_104),
.B1(n_89),
.B2(n_100),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_139),
.B1(n_146),
.B2(n_149),
.Y(n_170)
);

AND2x6_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_84),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_144),
.B(n_111),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_104),
.B1(n_89),
.B2(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_99),
.C(n_54),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_32),
.C(n_31),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_115),
.A2(n_101),
.B1(n_37),
.B2(n_44),
.Y(n_146)
);

BUFx24_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_110),
.B(n_78),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_63),
.B1(n_47),
.B2(n_76),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_126),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_152),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_127),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_143),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_153),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_154),
.A2(n_163),
.B(n_77),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_158),
.B(n_164),
.Y(n_177)
);

AO22x1_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_47),
.B1(n_118),
.B2(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_121),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_171),
.C(n_144),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_52),
.C(n_46),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_182),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

XNOR2x2_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_138),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_183),
.B(n_160),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_186),
.Y(n_195)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_133),
.B1(n_142),
.B2(n_147),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_170),
.B1(n_151),
.B2(n_165),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_88),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_165),
.B(n_173),
.Y(n_206)
);

XOR2x2_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_161),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_190),
.A2(n_160),
.B(n_173),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_157),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_198),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_205),
.C(n_191),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_203),
.C(n_207),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_183),
.A2(n_170),
.B1(n_156),
.B2(n_162),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_200),
.A2(n_201),
.B1(n_181),
.B2(n_184),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_169),
.C(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_77),
.C(n_46),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_10),
.C(n_9),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_210),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_45),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_194),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_200),
.A2(n_181),
.B1(n_177),
.B2(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_191),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_23),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_221),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_206),
.A3(n_190),
.B1(n_199),
.B2(n_179),
.C1(n_203),
.C2(n_207),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_225),
.B(n_226),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_198),
.A2(n_13),
.B1(n_19),
.B2(n_25),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_223),
.A2(n_11),
.B1(n_9),
.B2(n_8),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_45),
.C(n_32),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_45),
.C(n_16),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_11),
.C(n_7),
.Y(n_225)
);

AOI221xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_13),
.B1(n_25),
.B2(n_7),
.C(n_8),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_16),
.B1(n_20),
.B2(n_45),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_228),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_229),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_223),
.B1(n_219),
.B2(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_233),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_234),
.C(n_18),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_16),
.C(n_18),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_18),
.C(n_42),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_0),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_213),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_238),
.C(n_237),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_246),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_225),
.B(n_9),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_234),
.B(n_228),
.Y(n_252)
);

NOR2xp67_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_23),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_248),
.A2(n_42),
.B1(n_24),
.B2(n_20),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_235),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_242),
.Y(n_250)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_252),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_232),
.C(n_20),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_249),
.C(n_1),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_257),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_1),
.B(n_3),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_24),
.Y(n_261)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_262),
.B(n_0),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_0),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_265),
.A3(n_14),
.B1(n_260),
.B2(n_259),
.C1(n_5),
.C2(n_1),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_263),
.A2(n_256),
.B(n_28),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_3),
.C(n_4),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_268),
.C(n_3),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_4),
.B(n_5),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_4),
.B1(n_6),
.B2(n_14),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_4),
.C(n_6),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_272),
.A2(n_6),
.B(n_259),
.Y(n_273)
);


endmodule