module fake_jpeg_28139_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_14),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_18),
.B1(n_20),
.B2(n_16),
.Y(n_55)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_30),
.B1(n_23),
.B2(n_29),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_55),
.B1(n_18),
.B2(n_20),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_21),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_40),
.C(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_19),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_67),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_61),
.B(n_62),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_15),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_30),
.B1(n_23),
.B2(n_29),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_30),
.B1(n_31),
.B2(n_15),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NAND2x1p5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_34),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_28),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_80),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_27),
.B1(n_28),
.B2(n_18),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_79),
.B(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_24),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_82),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_20),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_37),
.Y(n_98)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_57),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_72),
.B1(n_61),
.B2(n_85),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_41),
.B1(n_60),
.B2(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_99),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_36),
.Y(n_143)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_109),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_73),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_65),
.C(n_34),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_122),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_52),
.B1(n_82),
.B2(n_41),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_117),
.A2(n_131),
.B1(n_105),
.B2(n_107),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_52),
.B1(n_53),
.B2(n_75),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_118),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_52),
.B1(n_78),
.B2(n_77),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_60),
.B1(n_32),
.B2(n_25),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_89),
.B1(n_111),
.B2(n_88),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_1),
.B(n_32),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_142),
.B(n_144),
.Y(n_155)
);

OAI22x1_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_19),
.B1(n_26),
.B2(n_35),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_88),
.A2(n_108),
.B1(n_98),
.B2(n_112),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_92),
.A2(n_40),
.B1(n_81),
.B2(n_86),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_16),
.B1(n_46),
.B2(n_36),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_36),
.C(n_46),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_123),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_93),
.B1(n_16),
.B2(n_102),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_141),
.A2(n_131),
.B(n_118),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_93),
.A2(n_25),
.B(n_24),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_94),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_95),
.A2(n_19),
.B(n_26),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_17),
.C(n_21),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_145),
.B(n_153),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_99),
.B(n_109),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_100),
.B(n_1),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_150),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_104),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_156),
.B(n_169),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_157),
.Y(n_184)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_159),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_121),
.B(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_168),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_177),
.B1(n_168),
.B2(n_172),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_119),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_162),
.B(n_165),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_101),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_163),
.B(n_164),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_130),
.A2(n_101),
.B(n_3),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_124),
.B(n_121),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_129),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_174),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_143),
.A3(n_122),
.B1(n_125),
.B2(n_139),
.C1(n_134),
.C2(n_127),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_180),
.B(n_158),
.CI(n_150),
.CON(n_216),
.SN(n_216)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_163),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_8),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_183),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_221)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_192),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_120),
.B1(n_107),
.B2(n_21),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_191),
.A2(n_148),
.B1(n_173),
.B2(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_21),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_206),
.Y(n_229)
);

XNOR2x2_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_17),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_164),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_57),
.C(n_17),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_197),
.C(n_170),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_145),
.B(n_57),
.C(n_17),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_201),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_148),
.B1(n_152),
.B2(n_160),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_14),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_146),
.B(n_174),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_217),
.B(n_179),
.Y(n_246)
);

INVxp33_ASAP7_75t_SL g210 ( 
.A(n_186),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_215),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_155),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_224),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_188),
.B(n_2),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_222),
.B(n_230),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_195),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_223),
.Y(n_233)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_226),
.C(n_207),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_8),
.C(n_9),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_225),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_198),
.B1(n_200),
.B2(n_185),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_245),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_234),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_209),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_239),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_208),
.A2(n_198),
.B(n_200),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_240),
.A2(n_246),
.B(n_229),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_226),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_196),
.C(n_207),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_247),
.C(n_212),
.Y(n_259)
);

OA22x2_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_183),
.B1(n_184),
.B2(n_186),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_197),
.C(n_193),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_253),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_258),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_241),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_263),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_208),
.B(n_218),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_240),
.B(n_254),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_257),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_261),
.C(n_244),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_260),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_216),
.C(n_190),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_248),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_249),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_264),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_223),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_273),
.C(n_265),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_236),
.C(n_242),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_261),
.C(n_258),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_275),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_236),
.B1(n_242),
.B2(n_233),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_276),
.A2(n_256),
.B1(n_238),
.B2(n_245),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_285),
.C(n_267),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_SL g281 ( 
.A(n_270),
.B(n_231),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_250),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_283),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_269),
.B(n_254),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_232),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_287),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_271),
.B1(n_266),
.B2(n_277),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_280),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_273),
.C(n_267),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_276),
.C(n_252),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_295),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_238),
.C(n_245),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_292),
.B(n_294),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_299),
.B(n_301),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_296),
.B(n_280),
.C(n_245),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_186),
.B(n_9),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_303),
.A2(n_298),
.B(n_9),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_304),
.A2(n_302),
.B(n_10),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_305),
.Y(n_306)
);

NOR3xp33_ASAP7_75t_SL g307 ( 
.A(n_306),
.B(n_8),
.C(n_10),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_10),
.B(n_11),
.C(n_305),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_11),
.Y(n_309)
);


endmodule