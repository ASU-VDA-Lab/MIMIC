module real_aes_8064_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_0), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g443 ( .A(n_0), .Y(n_443) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_1), .A2(n_148), .B(n_151), .C(n_231), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_2), .A2(n_177), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g508 ( .A(n_3), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_4), .B(n_207), .Y(n_206) );
AOI21xp33_ASAP7_75t_L g491 ( .A1(n_5), .A2(n_177), .B(n_492), .Y(n_491) );
AND2x6_ASAP7_75t_L g148 ( .A(n_6), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g244 ( .A(n_7), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_8), .B(n_43), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_9), .A2(n_176), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_10), .B(n_160), .Y(n_233) );
INVx1_ASAP7_75t_L g496 ( .A(n_11), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_12), .B(n_201), .Y(n_531) );
OAI22xp5_ASAP7_75t_SL g450 ( .A1(n_13), .A2(n_451), .B1(n_452), .B2(n_458), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_13), .Y(n_458) );
INVx1_ASAP7_75t_L g140 ( .A(n_14), .Y(n_140) );
INVx1_ASAP7_75t_L g543 ( .A(n_15), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_16), .A2(n_81), .B1(n_456), .B2(n_457), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_16), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_17), .A2(n_185), .B(n_266), .C(n_268), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_18), .B(n_207), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_19), .B(n_474), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_20), .B(n_177), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_21), .B(n_191), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_22), .A2(n_201), .B(n_252), .C(n_254), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_23), .B(n_207), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_24), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_25), .A2(n_187), .B(n_268), .C(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_26), .B(n_160), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g142 ( .A(n_27), .Y(n_142) );
INVx1_ASAP7_75t_L g214 ( .A(n_28), .Y(n_214) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_29), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_30), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_31), .B(n_160), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_32), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g183 ( .A(n_33), .Y(n_183) );
INVx1_ASAP7_75t_L g486 ( .A(n_34), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_35), .A2(n_453), .B1(n_454), .B2(n_455), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_35), .Y(n_453) );
INVx2_ASAP7_75t_L g146 ( .A(n_36), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_37), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_38), .A2(n_201), .B(n_202), .C(n_204), .Y(n_200) );
INVxp67_ASAP7_75t_L g186 ( .A(n_39), .Y(n_186) );
CKINVDCx14_ASAP7_75t_R g199 ( .A(n_40), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_41), .A2(n_151), .B(n_213), .C(n_217), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_42), .A2(n_148), .B(n_151), .C(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g485 ( .A(n_44), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_45), .A2(n_162), .B(n_242), .C(n_243), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_46), .B(n_160), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_47), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_48), .Y(n_179) );
INVx1_ASAP7_75t_L g250 ( .A(n_49), .Y(n_250) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_50), .A2(n_105), .B1(n_114), .B2(n_752), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_51), .Y(n_487) );
AOI222xp33_ASAP7_75t_SL g448 ( .A1(n_52), .A2(n_449), .B1(n_450), .B2(n_459), .C1(n_745), .C2(n_748), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g431 ( .A1(n_53), .A2(n_62), .B1(n_432), .B2(n_433), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_53), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_54), .B(n_177), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_55), .A2(n_151), .B1(n_254), .B2(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_56), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_57), .Y(n_505) );
CKINVDCx14_ASAP7_75t_R g240 ( .A(n_58), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_59), .A2(n_204), .B(n_242), .C(n_495), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_60), .A2(n_122), .B1(n_123), .B2(n_436), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_60), .Y(n_436) );
INVx1_ASAP7_75t_L g493 ( .A(n_61), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_62), .Y(n_433) );
INVx1_ASAP7_75t_L g149 ( .A(n_63), .Y(n_149) );
INVx1_ASAP7_75t_L g139 ( .A(n_64), .Y(n_139) );
INVx1_ASAP7_75t_SL g203 ( .A(n_65), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_66), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g430 ( .A1(n_67), .A2(n_431), .B1(n_434), .B2(n_435), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_67), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_68), .B(n_207), .Y(n_256) );
INVx1_ASAP7_75t_L g155 ( .A(n_69), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_SL g473 ( .A1(n_70), .A2(n_204), .B(n_474), .C(n_475), .Y(n_473) );
INVxp67_ASAP7_75t_L g476 ( .A(n_71), .Y(n_476) );
INVx1_ASAP7_75t_L g111 ( .A(n_72), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_73), .A2(n_177), .B(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_74), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_75), .A2(n_177), .B(n_263), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_76), .Y(n_489) );
INVx1_ASAP7_75t_L g549 ( .A(n_77), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_78), .A2(n_176), .B(n_178), .Y(n_175) );
CKINVDCx16_ASAP7_75t_R g211 ( .A(n_79), .Y(n_211) );
INVx1_ASAP7_75t_L g264 ( .A(n_80), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_81), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_82), .A2(n_148), .B(n_151), .C(n_551), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_83), .A2(n_177), .B(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g267 ( .A(n_84), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_85), .B(n_184), .Y(n_520) );
INVx2_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx1_ASAP7_75t_L g232 ( .A(n_87), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_88), .B(n_474), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_89), .A2(n_148), .B(n_151), .C(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g108 ( .A(n_90), .Y(n_108) );
OR2x2_ASAP7_75t_L g440 ( .A(n_90), .B(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g460 ( .A(n_90), .B(n_442), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_91), .A2(n_151), .B(n_154), .C(n_164), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_92), .B(n_169), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_93), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_94), .A2(n_148), .B(n_151), .C(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_95), .Y(n_535) );
INVx1_ASAP7_75t_L g472 ( .A(n_96), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_97), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_98), .B(n_184), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_99), .B(n_135), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_100), .B(n_135), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_101), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g253 ( .A(n_102), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_103), .A2(n_177), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_106), .Y(n_754) );
OR2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_112), .Y(n_106) );
OR2x2_ASAP7_75t_L g744 ( .A(n_108), .B(n_442), .Y(n_744) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_108), .B(n_441), .Y(n_747) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g442 ( .A(n_113), .B(n_443), .Y(n_442) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_447), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g751 ( .A(n_118), .Y(n_751) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_437), .B(n_444), .Y(n_120) );
INVxp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
XOR2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_430), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g459 ( .A1(n_124), .A2(n_460), .B1(n_461), .B2(n_742), .Y(n_459) );
INVx2_ASAP7_75t_L g749 ( .A(n_124), .Y(n_749) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_364), .Y(n_124) );
NAND5xp2_ASAP7_75t_L g125 ( .A(n_126), .B(n_293), .C(n_323), .D(n_344), .E(n_350), .Y(n_125) );
AOI221xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_223), .B1(n_257), .B2(n_259), .C(n_270), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_220), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_192), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_SL g344 ( .A1(n_131), .A2(n_208), .B(n_345), .C(n_348), .Y(n_344) );
AND2x2_ASAP7_75t_L g414 ( .A(n_131), .B(n_209), .Y(n_414) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_170), .Y(n_131) );
AND2x2_ASAP7_75t_L g272 ( .A(n_132), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g276 ( .A(n_132), .B(n_273), .Y(n_276) );
OR2x2_ASAP7_75t_L g302 ( .A(n_132), .B(n_209), .Y(n_302) );
AND2x2_ASAP7_75t_L g304 ( .A(n_132), .B(n_195), .Y(n_304) );
AND2x2_ASAP7_75t_L g322 ( .A(n_132), .B(n_194), .Y(n_322) );
INVx1_ASAP7_75t_L g355 ( .A(n_132), .Y(n_355) );
INVx2_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
BUFx2_ASAP7_75t_L g222 ( .A(n_133), .Y(n_222) );
AND2x2_ASAP7_75t_L g258 ( .A(n_133), .B(n_195), .Y(n_258) );
AND2x2_ASAP7_75t_L g411 ( .A(n_133), .B(n_209), .Y(n_411) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_166), .Y(n_133) );
INVx3_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_134), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_134), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_SL g522 ( .A(n_134), .B(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_135), .Y(n_196) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_135), .A2(n_470), .B(n_477), .Y(n_469) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_137), .B(n_138), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_150), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_143), .A2(n_169), .B(n_211), .C(n_212), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_143), .A2(n_229), .B(n_230), .Y(n_228) );
OAI22xp33_ASAP7_75t_L g482 ( .A1(n_143), .A2(n_165), .B1(n_483), .B2(n_487), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_143), .A2(n_505), .B(n_506), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_143), .A2(n_549), .B(n_550), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
AND2x4_ASAP7_75t_L g177 ( .A(n_144), .B(n_148), .Y(n_177) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
INVx1_ASAP7_75t_L g255 ( .A(n_146), .Y(n_255) );
INVx1_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_147), .Y(n_160) );
INVx3_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
INVx1_ASAP7_75t_L g474 ( .A(n_147), .Y(n_474) );
INVx4_ASAP7_75t_SL g165 ( .A(n_148), .Y(n_165) );
BUFx3_ASAP7_75t_L g217 ( .A(n_148), .Y(n_217) );
INVx5_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx3_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_152), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_159), .C(n_161), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_L g231 ( .A1(n_156), .A2(n_161), .B(n_232), .C(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g484 ( .A1(n_157), .A2(n_158), .B1(n_485), .B2(n_486), .Y(n_484) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx4_ASAP7_75t_L g187 ( .A(n_158), .Y(n_187) );
INVx4_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
INVx2_ASAP7_75t_L g242 ( .A(n_160), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_161), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_161), .A2(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g268 ( .A(n_163), .Y(n_268) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_SL g178 ( .A1(n_165), .A2(n_179), .B(n_180), .C(n_181), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_165), .A2(n_180), .B(n_199), .C(n_200), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_SL g239 ( .A1(n_165), .A2(n_180), .B(n_240), .C(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_165), .A2(n_180), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_SL g263 ( .A1(n_165), .A2(n_180), .B(n_264), .C(n_265), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_165), .A2(n_180), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_165), .A2(n_180), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_165), .A2(n_180), .B(n_540), .C(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx1_ASAP7_75t_L g191 ( .A(n_168), .Y(n_191) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_168), .A2(n_527), .B(n_534), .Y(n_526) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_169), .A2(n_238), .B(n_245), .Y(n_237) );
OA21x2_ASAP7_75t_L g537 ( .A1(n_169), .A2(n_538), .B(n_544), .Y(n_537) );
AND2x2_ASAP7_75t_L g292 ( .A(n_170), .B(n_193), .Y(n_292) );
OR2x2_ASAP7_75t_L g296 ( .A(n_170), .B(n_209), .Y(n_296) );
AND2x2_ASAP7_75t_L g321 ( .A(n_170), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g368 ( .A(n_170), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_170), .B(n_330), .Y(n_416) );
AO21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_174), .B(n_189), .Y(n_170) );
INVx1_ASAP7_75t_L g274 ( .A(n_171), .Y(n_274) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_171), .A2(n_548), .B(n_554), .Y(n_547) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_SL g516 ( .A1(n_172), .A2(n_517), .B(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_173), .A2(n_482), .B(n_488), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_173), .B(n_489), .Y(n_488) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_173), .A2(n_504), .B(n_511), .Y(n_503) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_175), .A2(n_190), .B(n_274), .Y(n_273) );
BUFx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_182), .B(n_188), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B1(n_186), .B2(n_187), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_184), .A2(n_214), .B(n_215), .C(n_216), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_184), .A2(n_508), .B(n_509), .C(n_510), .Y(n_507) );
INVx5_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_185), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_185), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_185), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_187), .B(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_187), .B(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_187), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g216 ( .A(n_188), .Y(n_216) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI322xp33_ASAP7_75t_L g417 ( .A1(n_192), .A2(n_353), .A3(n_376), .B1(n_397), .B2(n_418), .C1(n_420), .C2(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_193), .B(n_273), .Y(n_420) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_208), .Y(n_193) );
AND2x2_ASAP7_75t_L g221 ( .A(n_194), .B(n_222), .Y(n_221) );
AND2x4_ASAP7_75t_L g289 ( .A(n_194), .B(n_209), .Y(n_289) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g330 ( .A(n_195), .B(n_209), .Y(n_330) );
AND2x2_ASAP7_75t_L g374 ( .A(n_195), .B(n_208), .Y(n_374) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_206), .Y(n_195) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_196), .A2(n_248), .B(n_256), .Y(n_247) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_196), .A2(n_262), .B(n_269), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_201), .B(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_205), .Y(n_532) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_207), .A2(n_491), .B(n_497), .Y(n_490) );
AND2x2_ASAP7_75t_L g257 ( .A(n_208), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g275 ( .A(n_208), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_208), .B(n_304), .Y(n_428) );
INVx3_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g220 ( .A(n_209), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_209), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g342 ( .A(n_209), .B(n_273), .Y(n_342) );
AND2x2_ASAP7_75t_L g369 ( .A(n_209), .B(n_304), .Y(n_369) );
OR2x2_ASAP7_75t_L g425 ( .A(n_209), .B(n_276), .Y(n_425) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_218), .Y(n_209) );
INVx1_ASAP7_75t_SL g311 ( .A(n_220), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_221), .B(n_342), .Y(n_343) );
AND2x2_ASAP7_75t_L g377 ( .A(n_221), .B(n_367), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_221), .B(n_300), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_221), .B(n_422), .Y(n_421) );
OAI31xp33_ASAP7_75t_L g395 ( .A1(n_223), .A2(n_257), .A3(n_396), .B(n_398), .Y(n_395) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_236), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g362 ( .A(n_224), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g378 ( .A(n_224), .B(n_313), .Y(n_378) );
OR2x2_ASAP7_75t_L g385 ( .A(n_224), .B(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g397 ( .A(n_224), .B(n_286), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g331 ( .A(n_225), .B(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g259 ( .A(n_226), .B(n_260), .Y(n_259) );
INVx4_ASAP7_75t_L g280 ( .A(n_226), .Y(n_280) );
AND2x2_ASAP7_75t_L g317 ( .A(n_226), .B(n_261), .Y(n_317) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_234), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_227), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_227), .B(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_227), .B(n_436), .Y(n_554) );
AND2x2_ASAP7_75t_L g316 ( .A(n_236), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g386 ( .A(n_236), .Y(n_386) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_246), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_237), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g286 ( .A(n_237), .B(n_247), .Y(n_286) );
INVx2_ASAP7_75t_L g306 ( .A(n_237), .Y(n_306) );
AND2x2_ASAP7_75t_L g320 ( .A(n_237), .B(n_247), .Y(n_320) );
AND2x2_ASAP7_75t_L g327 ( .A(n_237), .B(n_283), .Y(n_327) );
BUFx3_ASAP7_75t_L g337 ( .A(n_237), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_237), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g282 ( .A(n_246), .Y(n_282) );
AND2x2_ASAP7_75t_L g290 ( .A(n_246), .B(n_280), .Y(n_290) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g260 ( .A(n_247), .B(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_247), .Y(n_314) );
INVx2_ASAP7_75t_L g510 ( .A(n_254), .Y(n_510) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_SL g297 ( .A(n_258), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_258), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_258), .B(n_367), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_259), .B(n_337), .Y(n_390) );
INVx1_ASAP7_75t_SL g424 ( .A(n_259), .Y(n_424) );
INVx1_ASAP7_75t_SL g332 ( .A(n_260), .Y(n_332) );
INVx1_ASAP7_75t_SL g283 ( .A(n_261), .Y(n_283) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_261), .Y(n_294) );
OR2x2_ASAP7_75t_L g305 ( .A(n_261), .B(n_280), .Y(n_305) );
AND2x2_ASAP7_75t_L g319 ( .A(n_261), .B(n_280), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_261), .B(n_309), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_275), .B(n_277), .C(n_288), .Y(n_270) );
AOI31xp33_ASAP7_75t_L g387 ( .A1(n_271), .A2(n_388), .A3(n_389), .B(n_390), .Y(n_387) );
AND2x2_ASAP7_75t_L g360 ( .A(n_272), .B(n_289), .Y(n_360) );
BUFx3_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_273), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g336 ( .A(n_273), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_273), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g291 ( .A(n_276), .Y(n_291) );
OAI222xp33_ASAP7_75t_L g400 ( .A1(n_276), .A2(n_401), .B1(n_404), .B2(n_405), .C1(n_406), .C2(n_407), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_284), .Y(n_277) );
INVx1_ASAP7_75t_L g406 ( .A(n_278), .Y(n_406) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_280), .B(n_283), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_280), .B(n_306), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_280), .B(n_281), .Y(n_376) );
INVx1_ASAP7_75t_L g427 ( .A(n_280), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_281), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g429 ( .A(n_281), .Y(n_429) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx2_ASAP7_75t_L g309 ( .A(n_282), .Y(n_309) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_283), .Y(n_352) );
AOI32xp33_ASAP7_75t_L g288 ( .A1(n_284), .A2(n_289), .A3(n_290), .B1(n_291), .B2(n_292), .Y(n_288) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_286), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g363 ( .A(n_286), .Y(n_363) );
OR2x2_ASAP7_75t_L g404 ( .A(n_286), .B(n_305), .Y(n_404) );
INVx1_ASAP7_75t_L g340 ( .A(n_287), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_289), .B(n_300), .Y(n_325) );
INVx3_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
AOI322xp5_ASAP7_75t_L g350 ( .A1(n_289), .A2(n_334), .A3(n_351), .B1(n_353), .B2(n_356), .C1(n_360), .C2(n_361), .Y(n_350) );
AND2x2_ASAP7_75t_L g326 ( .A(n_290), .B(n_327), .Y(n_326) );
INVxp67_ASAP7_75t_L g403 ( .A(n_290), .Y(n_403) );
A2O1A1O1Ixp25_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B(n_298), .C(n_306), .D(n_307), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_294), .B(n_337), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
OAI221xp5_ASAP7_75t_L g307 ( .A1(n_296), .A2(n_308), .B1(n_311), .B2(n_312), .C(n_315), .Y(n_307) );
INVx1_ASAP7_75t_SL g422 ( .A(n_296), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_303), .B(n_305), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_300), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI221xp5_ASAP7_75t_SL g392 ( .A1(n_302), .A2(n_386), .B1(n_393), .B2(n_394), .C(n_395), .Y(n_392) );
OAI222xp33_ASAP7_75t_L g423 ( .A1(n_303), .A2(n_424), .B1(n_425), .B2(n_426), .C1(n_428), .C2(n_429), .Y(n_423) );
AND2x2_ASAP7_75t_L g381 ( .A(n_304), .B(n_367), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_304), .A2(n_319), .B(n_366), .Y(n_393) );
INVx1_ASAP7_75t_L g407 ( .A(n_304), .Y(n_407) );
INVx2_ASAP7_75t_SL g310 ( .A(n_305), .Y(n_310) );
AND2x2_ASAP7_75t_L g313 ( .A(n_306), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_SL g347 ( .A(n_309), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_309), .B(n_319), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_310), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_310), .B(n_320), .Y(n_349) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI21xp5_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_318), .B(n_321), .Y(n_315) );
INVx1_ASAP7_75t_SL g333 ( .A(n_317), .Y(n_333) );
AND2x2_ASAP7_75t_L g380 ( .A(n_317), .B(n_363), .Y(n_380) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x2_ASAP7_75t_L g419 ( .A(n_319), .B(n_337), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_320), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g405 ( .A(n_321), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_326), .B1(n_328), .B2(n_335), .C(n_338), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B1(n_333), .B2(n_334), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_332), .A2(n_339), .B1(n_341), .B2(n_343), .Y(n_338) );
OR2x2_ASAP7_75t_L g409 ( .A(n_333), .B(n_337), .Y(n_409) );
OR2x2_ASAP7_75t_L g412 ( .A(n_333), .B(n_347), .Y(n_412) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_354), .A2(n_409), .B1(n_410), .B2(n_412), .C(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND3xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_379), .C(n_391), .Y(n_364) );
AOI222xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_370), .B1(n_372), .B2(n_375), .C1(n_377), .C2(n_378), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_367), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g389 ( .A(n_369), .Y(n_389) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_382), .B2(n_384), .C(n_387), .Y(n_379) );
INVx1_ASAP7_75t_L g394 ( .A(n_380), .Y(n_394) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI21xp33_ASAP7_75t_L g413 ( .A1(n_384), .A2(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
NOR5xp2_ASAP7_75t_L g391 ( .A(n_392), .B(n_400), .C(n_408), .D(n_417), .E(n_423), .Y(n_391) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_431), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g446 ( .A(n_440), .Y(n_446) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_444), .B(n_448), .C(n_750), .Y(n_447) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_460), .A2(n_462), .B1(n_742), .B2(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_SL g462 ( .A(n_463), .B(n_679), .Y(n_462) );
NOR4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_609), .C(n_640), .D(n_659), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_465), .B(n_567), .C(n_582), .D(n_600), .Y(n_464) );
AOI222xp33_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_513), .B1(n_545), .B2(n_555), .C1(n_560), .C2(n_562), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_498), .Y(n_466) );
INVx1_ASAP7_75t_L g623 ( .A(n_467), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
AND2x2_ASAP7_75t_L g499 ( .A(n_468), .B(n_490), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_468), .B(n_502), .Y(n_652) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g559 ( .A(n_469), .B(n_480), .Y(n_559) );
AND2x2_ASAP7_75t_L g568 ( .A(n_469), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g594 ( .A(n_469), .Y(n_594) );
AND2x2_ASAP7_75t_L g615 ( .A(n_469), .B(n_480), .Y(n_615) );
BUFx2_ASAP7_75t_L g638 ( .A(n_469), .Y(n_638) );
AND2x2_ASAP7_75t_L g662 ( .A(n_469), .B(n_481), .Y(n_662) );
AND2x2_ASAP7_75t_L g726 ( .A(n_469), .B(n_490), .Y(n_726) );
AND2x2_ASAP7_75t_L g627 ( .A(n_478), .B(n_558), .Y(n_627) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_479), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_490), .Y(n_479) );
OR2x2_ASAP7_75t_L g587 ( .A(n_480), .B(n_503), .Y(n_587) );
AND2x2_ASAP7_75t_L g599 ( .A(n_480), .B(n_558), .Y(n_599) );
BUFx2_ASAP7_75t_L g731 ( .A(n_480), .Y(n_731) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g501 ( .A(n_481), .B(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g581 ( .A(n_481), .B(n_503), .Y(n_581) );
AND2x2_ASAP7_75t_L g634 ( .A(n_481), .B(n_490), .Y(n_634) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_481), .Y(n_670) );
AND2x2_ASAP7_75t_L g557 ( .A(n_490), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_SL g569 ( .A(n_490), .Y(n_569) );
INVx2_ASAP7_75t_L g580 ( .A(n_490), .Y(n_580) );
BUFx2_ASAP7_75t_L g604 ( .A(n_490), .Y(n_604) );
AND2x2_ASAP7_75t_SL g661 ( .A(n_490), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
AOI332xp33_ASAP7_75t_L g582 ( .A1(n_499), .A2(n_583), .A3(n_587), .B1(n_588), .B2(n_592), .B3(n_595), .C1(n_596), .C2(n_598), .Y(n_582) );
NAND2x1_ASAP7_75t_L g667 ( .A(n_499), .B(n_558), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_499), .B(n_572), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_SL g600 ( .A1(n_500), .A2(n_601), .B(n_604), .C(n_605), .Y(n_600) );
AND2x2_ASAP7_75t_L g739 ( .A(n_500), .B(n_580), .Y(n_739) );
INVx3_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g636 ( .A(n_501), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g641 ( .A(n_501), .B(n_638), .Y(n_641) );
INVx1_ASAP7_75t_L g572 ( .A(n_502), .Y(n_572) );
AND2x2_ASAP7_75t_L g675 ( .A(n_502), .B(n_634), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_502), .B(n_615), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_502), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_502), .B(n_593), .Y(n_701) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g558 ( .A(n_503), .Y(n_558) );
OAI31xp33_ASAP7_75t_L g740 ( .A1(n_513), .A2(n_661), .A3(n_668), .B(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_524), .Y(n_513) );
AND2x2_ASAP7_75t_L g545 ( .A(n_514), .B(n_546), .Y(n_545) );
NAND2x1_ASAP7_75t_SL g563 ( .A(n_514), .B(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_514), .Y(n_650) );
AND2x2_ASAP7_75t_L g655 ( .A(n_514), .B(n_566), .Y(n_655) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_515), .A2(n_568), .B(n_570), .C(n_573), .Y(n_567) );
OR2x2_ASAP7_75t_L g584 ( .A(n_515), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g597 ( .A(n_515), .Y(n_597) );
AND2x2_ASAP7_75t_L g603 ( .A(n_515), .B(n_547), .Y(n_603) );
INVx2_ASAP7_75t_L g621 ( .A(n_515), .Y(n_621) );
AND2x2_ASAP7_75t_L g632 ( .A(n_515), .B(n_586), .Y(n_632) );
AND2x2_ASAP7_75t_L g664 ( .A(n_515), .B(n_622), .Y(n_664) );
AND2x2_ASAP7_75t_L g668 ( .A(n_515), .B(n_591), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_515), .B(n_524), .Y(n_673) );
AND2x2_ASAP7_75t_L g707 ( .A(n_515), .B(n_708), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_515), .B(n_610), .Y(n_741) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_522), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_524), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g649 ( .A(n_524), .Y(n_649) );
AND2x2_ASAP7_75t_L g711 ( .A(n_524), .B(n_632), .Y(n_711) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_536), .Y(n_524) );
OR2x2_ASAP7_75t_L g565 ( .A(n_525), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g575 ( .A(n_525), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_525), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g683 ( .A(n_525), .Y(n_683) );
AND2x2_ASAP7_75t_L g700 ( .A(n_525), .B(n_547), .Y(n_700) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g591 ( .A(n_526), .B(n_536), .Y(n_591) );
AND2x2_ASAP7_75t_L g620 ( .A(n_526), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g631 ( .A(n_526), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_526), .B(n_586), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_533), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_532), .Y(n_529) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g546 ( .A(n_537), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g566 ( .A(n_537), .Y(n_566) );
AND2x2_ASAP7_75t_L g622 ( .A(n_537), .B(n_586), .Y(n_622) );
INVx1_ASAP7_75t_L g724 ( .A(n_545), .Y(n_724) );
INVx1_ASAP7_75t_L g728 ( .A(n_546), .Y(n_728) );
INVx2_ASAP7_75t_L g586 ( .A(n_547), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_557), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_557), .B(n_662), .Y(n_720) );
OR2x2_ASAP7_75t_L g561 ( .A(n_558), .B(n_559), .Y(n_561) );
INVx1_ASAP7_75t_SL g613 ( .A(n_558), .Y(n_613) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_564), .A2(n_617), .B1(n_619), .B2(n_623), .C(n_624), .Y(n_616) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g644 ( .A(n_565), .B(n_608), .Y(n_644) );
INVx2_ASAP7_75t_L g576 ( .A(n_566), .Y(n_576) );
INVx1_ASAP7_75t_L g602 ( .A(n_566), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_566), .B(n_586), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_566), .B(n_589), .Y(n_696) );
INVx1_ASAP7_75t_L g704 ( .A(n_566), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_568), .B(n_572), .Y(n_618) );
AND2x4_ASAP7_75t_L g593 ( .A(n_569), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g706 ( .A(n_572), .B(n_662), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_575), .B(n_607), .Y(n_606) );
INVxp67_ASAP7_75t_L g714 ( .A(n_576), .Y(n_714) );
INVxp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g614 ( .A(n_580), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g686 ( .A(n_580), .B(n_662), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_580), .B(n_599), .Y(n_692) );
AOI322xp5_ASAP7_75t_L g646 ( .A1(n_581), .A2(n_615), .A3(n_622), .B1(n_647), .B2(n_650), .C1(n_651), .C2(n_653), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_581), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g712 ( .A(n_584), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g658 ( .A(n_585), .Y(n_658) );
INVx2_ASAP7_75t_L g589 ( .A(n_586), .Y(n_589) );
INVx1_ASAP7_75t_L g648 ( .A(n_586), .Y(n_648) );
CKINVDCx16_ASAP7_75t_R g595 ( .A(n_587), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x2_ASAP7_75t_L g684 ( .A(n_589), .B(n_597), .Y(n_684) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g596 ( .A(n_591), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g639 ( .A(n_591), .B(n_632), .Y(n_639) );
AND2x2_ASAP7_75t_L g643 ( .A(n_591), .B(n_603), .Y(n_643) );
OAI21xp33_ASAP7_75t_SL g653 ( .A1(n_592), .A2(n_654), .B(n_656), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g723 ( .A1(n_592), .A2(n_724), .B1(n_725), .B2(n_727), .Y(n_723) );
INVx3_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g598 ( .A(n_593), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_593), .B(n_613), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_595), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g735 ( .A(n_602), .Y(n_735) );
INVx4_ASAP7_75t_L g608 ( .A(n_603), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_603), .B(n_630), .Y(n_678) );
INVx1_ASAP7_75t_SL g690 ( .A(n_604), .Y(n_690) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g703 ( .A(n_608), .B(n_704), .Y(n_703) );
OAI211xp5_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_611), .B(n_616), .C(n_633), .Y(n_609) );
OAI221xp5_ASAP7_75t_SL g729 ( .A1(n_611), .A2(n_649), .B1(n_728), .B2(n_730), .C(n_732), .Y(n_729) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_613), .B(n_726), .Y(n_725) );
OAI31xp33_ASAP7_75t_L g705 ( .A1(n_614), .A2(n_691), .A3(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g645 ( .A(n_615), .Y(n_645) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx1_ASAP7_75t_L g695 ( .A(n_620), .Y(n_695) );
AND2x2_ASAP7_75t_L g708 ( .A(n_622), .B(n_631), .Y(n_708) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_628), .Y(n_624) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_632), .B(n_735), .Y(n_734) );
OAI21xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B(n_639), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI221xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_642), .B1(n_644), .B2(n_645), .C(n_646), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_L g709 ( .A1(n_641), .A2(n_710), .B(n_712), .C(n_715), .Y(n_709) );
CKINVDCx16_ASAP7_75t_R g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_644), .B(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g671 ( .A(n_652), .Y(n_671) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g657 ( .A(n_655), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g699 ( .A(n_655), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI211xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_665), .C(n_674), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_663), .A2(n_673), .B1(n_737), .B2(n_738), .C(n_740), .Y(n_736) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B1(n_669), .B2(n_672), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI21xp5_ASAP7_75t_SL g674 ( .A1(n_675), .A2(n_676), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_SL g737 ( .A(n_676), .Y(n_737) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR4xp25_ASAP7_75t_L g679 ( .A(n_680), .B(n_709), .C(n_729), .D(n_736), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_685), .B(n_687), .C(n_705), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_691), .B(n_693), .C(n_697), .Y(n_687) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g716 ( .A(n_694), .Y(n_716) );
OR2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
OR2x2_ASAP7_75t_L g727 ( .A(n_695), .B(n_728), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_701), .B(n_702), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_719), .B2(n_721), .C(n_723), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_726), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
endmodule