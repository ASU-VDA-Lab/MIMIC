module fake_jpeg_26186_n_105 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_1),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_62),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_42),
.Y(n_73)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_56),
.B1(n_47),
.B2(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_74),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_56),
.B1(n_54),
.B2(n_46),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_69),
.A2(n_72),
.B1(n_3),
.B2(n_4),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_43),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_1),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_2),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_78),
.A2(n_83),
.B1(n_4),
.B2(n_5),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_81),
.B1(n_67),
.B2(n_76),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_25),
.C(n_38),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_81),
.A2(n_69),
.B1(n_72),
.B2(n_70),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_85),
.B1(n_79),
.B2(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_82),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_6),
.Y(n_92)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_89),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_27),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_6),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_92),
.B(n_9),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_7),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_95),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_97),
.A2(n_91),
.B(n_13),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_12),
.B(n_14),
.C(n_16),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_17),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_23),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_30),
.B(n_32),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_33),
.B(n_34),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_37),
.B(n_39),
.Y(n_105)
);


endmodule