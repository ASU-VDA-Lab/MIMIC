module fake_jpeg_31631_n_152 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_0),
.B(n_6),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_62),
.Y(n_77)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_53),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_77),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_52),
.B1(n_54),
.B2(n_49),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_57),
.B1(n_55),
.B2(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_60),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_64),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_64),
.B(n_56),
.C(n_61),
.Y(n_86)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_50),
.B1(n_49),
.B2(n_51),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_16),
.B(n_17),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_96),
.Y(n_100)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_51),
.B(n_45),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_5),
.B(n_7),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_0),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_8),
.B1(n_9),
.B2(n_44),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_79),
.B1(n_74),
.B2(n_76),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_12),
.B(n_13),
.C(n_15),
.Y(n_115)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_103),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_107),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_92),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_108),
.B1(n_114),
.B2(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_4),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_116),
.B(n_18),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_24),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_43),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_31),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_118),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_100),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_20),
.B(n_22),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_130),
.B(n_37),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_115),
.A2(n_23),
.B1(n_27),
.B2(n_29),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_127),
.B(n_128),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_34),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_32),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_42),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_137),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_142),
.B1(n_129),
.B2(n_131),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_121),
.C(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_141),
.Y(n_144)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_141),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_144),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_139),
.B(n_123),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_138),
.B(n_124),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_150),
.A2(n_136),
.B(n_135),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_40),
.Y(n_152)
);


endmodule