module fake_jpeg_25150_n_202 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_13),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_39),
.Y(n_51)
);

CKINVDCx12_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_13),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_25),
.B(n_33),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_13),
.B1(n_20),
.B2(n_16),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_52),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_27),
.B1(n_29),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_27),
.B1(n_29),
.B2(n_24),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_20),
.B1(n_16),
.B2(n_11),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_10),
.B1(n_19),
.B2(n_11),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_10),
.B(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_31),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_39),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_68),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_70),
.B1(n_73),
.B2(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_72),
.B(n_22),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_38),
.B1(n_30),
.B2(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_78),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_49),
.Y(n_76)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_84),
.B(n_88),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_51),
.C(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_56),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_49),
.B1(n_10),
.B2(n_19),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_90),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_61),
.A2(n_49),
.B1(n_31),
.B2(n_43),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_73),
.B1(n_71),
.B2(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_52),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_23),
.B1(n_24),
.B2(n_57),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_18),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_12),
.B1(n_28),
.B2(n_22),
.Y(n_114)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_55),
.B(n_27),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_67),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_87),
.B1(n_85),
.B2(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_97),
.B(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_59),
.C(n_28),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_115),
.C(n_89),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

AO22x1_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_23),
.B1(n_50),
.B2(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_112),
.Y(n_132)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_110),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_80),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_12),
.B1(n_50),
.B2(n_28),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_22),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_18),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_117),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_22),
.C(n_14),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_18),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_18),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_118),
.A2(n_122),
.B1(n_125),
.B2(n_94),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_114),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_79),
.B1(n_75),
.B2(n_84),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_74),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_81),
.B1(n_76),
.B2(n_14),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_107),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_15),
.B(n_14),
.C(n_6),
.D(n_8),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_134),
.B(n_111),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_14),
.C(n_15),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_138),
.C(n_139),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_0),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_95),
.A2(n_0),
.B(n_1),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_15),
.C(n_6),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_7),
.C(n_9),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_96),
.B(n_101),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_141),
.A2(n_134),
.B(n_137),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_115),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_150),
.C(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_105),
.C(n_111),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_153),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_135),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_121),
.B1(n_128),
.B2(n_133),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_150),
.B1(n_144),
.B2(n_147),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_142),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_121),
.C(n_139),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_161),
.C(n_142),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_128),
.C(n_105),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_131),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_164),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_174),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_171),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_156),
.B(n_162),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_158),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_175),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_157),
.B1(n_147),
.B2(n_160),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_167),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_159),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_179),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_171),
.C(n_168),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_186),
.C(n_109),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_181),
.B(n_119),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_180),
.B(n_136),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_188),
.B(n_184),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_176),
.A2(n_163),
.B(n_110),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_192),
.B(n_7),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_182),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_193),
.C(n_111),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_188),
.A2(n_177),
.B(n_129),
.Y(n_192)
);

NOR2x1_ASAP7_75t_R g198 ( 
.A(n_194),
.B(n_196),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_195),
.A2(n_189),
.B(n_4),
.Y(n_197)
);

OAI221xp5_ASAP7_75t_SL g196 ( 
.A1(n_192),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.C(n_5),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_198),
.B(n_4),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_1),
.B(n_4),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_5),
.Y(n_202)
);


endmodule