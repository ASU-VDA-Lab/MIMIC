module fake_jpeg_15527_n_352 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_352);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_352;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_44),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_19),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_18),
.B(n_27),
.C(n_29),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_53),
.A2(n_30),
.B(n_1),
.C(n_2),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_59),
.B1(n_74),
.B2(n_28),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_22),
.B1(n_33),
.B2(n_24),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_57),
.A2(n_67),
.B1(n_73),
.B2(n_35),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_22),
.B1(n_24),
.B2(n_20),
.Y(n_59)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_36),
.C(n_25),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_30),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_35),
.B1(n_23),
.B2(n_28),
.Y(n_67)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_39),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_29),
.B1(n_27),
.B2(n_18),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_29),
.B1(n_27),
.B2(n_18),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_26),
.B1(n_20),
.B2(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_76),
.A2(n_86),
.B1(n_95),
.B2(n_63),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_82),
.Y(n_113)
);

OR2x4_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx2_ASAP7_75t_SL g110 ( 
.A(n_87),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_46),
.B1(n_45),
.B2(n_42),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_90),
.B1(n_102),
.B2(n_71),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_26),
.B1(n_20),
.B2(n_32),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_89),
.A2(n_92),
.B1(n_97),
.B2(n_71),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_45),
.B1(n_33),
.B2(n_26),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_94),
.B(n_73),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_92)
);

NAND3xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_41),
.C(n_16),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_25),
.B1(n_36),
.B2(n_30),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_30),
.B1(n_15),
.B2(n_14),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_41),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_25),
.B1(n_36),
.B2(n_30),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_58),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_104),
.B(n_69),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_113),
.B1(n_129),
.B2(n_101),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_55),
.C(n_68),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_83),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_112),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_131),
.Y(n_137)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_70),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_124),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_122),
.B(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_62),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_62),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

AO22x2_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_68),
.B1(n_71),
.B2(n_63),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_51),
.B1(n_93),
.B2(n_85),
.Y(n_155)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_100),
.Y(n_142)
);

AOI22x1_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_94),
.B1(n_103),
.B2(n_91),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_135),
.A2(n_141),
.B(n_151),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_80),
.C(n_77),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_153),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_150),
.B1(n_161),
.B2(n_162),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_113),
.B(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_142),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_103),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_148),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_81),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_91),
.B1(n_90),
.B2(n_88),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_102),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_93),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_160),
.B(n_114),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_133),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_125),
.B1(n_112),
.B2(n_134),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_106),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_110),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_15),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_118),
.A2(n_104),
.B(n_99),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_51),
.B1(n_85),
.B2(n_69),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_118),
.A2(n_51),
.B1(n_65),
.B2(n_79),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_98),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_164),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_123),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_168),
.B(n_180),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_167),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_108),
.B(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_109),
.Y(n_172)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_179),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_128),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_185),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_139),
.A2(n_150),
.B1(n_135),
.B2(n_151),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_177),
.B1(n_158),
.B2(n_65),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_161),
.B1(n_152),
.B2(n_154),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_186),
.C(n_145),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_105),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_58),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_146),
.B(n_125),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_162),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_193),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_130),
.B1(n_116),
.B2(n_131),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_0),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_127),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_192),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_127),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_196),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_65),
.B1(n_96),
.B2(n_83),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_144),
.B1(n_154),
.B2(n_137),
.Y(n_198)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_198),
.A2(n_200),
.B1(n_205),
.B2(n_215),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_145),
.B1(n_155),
.B2(n_136),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_224),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_164),
.C(n_83),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_179),
.A2(n_156),
.B1(n_83),
.B2(n_55),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_48),
.CI(n_55),
.CON(n_206),
.SN(n_206)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_206),
.B(n_219),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_106),
.C(n_96),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_48),
.C(n_14),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_213),
.Y(n_253)
);

NOR3xp33_ASAP7_75t_SL g210 ( 
.A(n_169),
.B(n_12),
.C(n_11),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_173),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_48),
.C(n_12),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_220),
.B(n_191),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_48),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_223),
.B1(n_166),
.B2(n_6),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_192),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_12),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_173),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_183),
.Y(n_227)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_228),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_230),
.B(n_235),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_197),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_236),
.B(n_251),
.Y(n_263)
);

NAND2x1p5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_167),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_214),
.B1(n_187),
.B2(n_206),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_166),
.Y(n_238)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_245),
.Y(n_262)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_166),
.B1(n_177),
.B2(n_176),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_185),
.B1(n_187),
.B2(n_180),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_252),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_204),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_171),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_189),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_254),
.A2(n_223),
.B1(n_215),
.B2(n_221),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_202),
.C(n_208),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_257),
.C(n_258),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_201),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_212),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_259),
.A2(n_184),
.B1(n_196),
.B2(n_188),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_214),
.B1(n_198),
.B2(n_203),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_261),
.A2(n_233),
.B1(n_241),
.B2(n_229),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_212),
.C(n_206),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_270),
.C(n_273),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_209),
.C(n_213),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_237),
.B(n_224),
.C(n_168),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_253),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_231),
.B(n_174),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_210),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_253),
.C(n_229),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_266),
.B(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_240),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_281),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_250),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_284),
.C(n_291),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_250),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_288),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_262),
.A2(n_237),
.B(n_245),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_287),
.A2(n_269),
.B(n_259),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_292),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_260),
.A2(n_239),
.B1(n_238),
.B2(n_252),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_243),
.B1(n_242),
.B2(n_228),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_184),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_258),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_293),
.B(n_264),
.Y(n_297)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_311),
.B(n_287),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_257),
.C(n_267),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_7),
.C(n_8),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_290),
.A2(n_276),
.B1(n_274),
.B2(n_272),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_308),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_303),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_285),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_307),
.B(n_7),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_261),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_270),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_308),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_284),
.A2(n_283),
.B(n_288),
.Y(n_311)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_313),
.B(n_319),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_292),
.B(n_295),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_315),
.B(n_318),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_298),
.A2(n_277),
.B(n_291),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_316),
.A2(n_309),
.B(n_304),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_285),
.B(n_7),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_5),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_7),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_314),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_330),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_301),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_300),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_333),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_302),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_334),
.A2(n_312),
.B(n_316),
.Y(n_337)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_337),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_317),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_338),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_334),
.A2(n_328),
.B(n_332),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_339),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_320),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_SL g344 ( 
.A1(n_340),
.A2(n_341),
.B(n_342),
.C(n_8),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_325),
.A2(n_310),
.B(n_9),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_344),
.A2(n_8),
.B(n_9),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_347),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_343),
.A2(n_336),
.B(n_335),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_348),
.B(n_346),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_345),
.C(n_10),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_10),
.Y(n_352)
);


endmodule