module fake_jpeg_19604_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_0),
.B(n_2),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

AND2x2_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_4),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_7),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_14),
.A2(n_9),
.B1(n_11),
.B2(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_8),
.B(n_6),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_15),
.A2(n_16),
.B(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_20),
.B(n_9),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_12),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_17),
.Y(n_28)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_21),
.B(n_15),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_28),
.B(n_29),
.Y(n_30)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_22),
.C(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_27),
.B1(n_29),
.B2(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_34),
.Y(n_37)
);


endmodule