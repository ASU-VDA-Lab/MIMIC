module fake_netlist_6_307_n_881 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_881);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_881;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_624;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_652;
wire n_553;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_612;
wire n_453;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_197),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_99),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_65),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_140),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_86),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_121),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_16),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_164),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_186),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_194),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_16),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_73),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_34),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_184),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_69),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_17),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_0),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_179),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_115),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_84),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_3),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_134),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_93),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_75),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_12),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_9),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_29),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_57),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_37),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_128),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_27),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_32),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_49),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_141),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_48),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_74),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_45),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_162),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_132),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_183),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_25),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_189),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_147),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_108),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_163),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_91),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_2),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_110),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_78),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_28),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_10),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_10),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_85),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_169),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_19),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_160),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_152),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_68),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_178),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_193),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_216),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_213),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_0),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_213),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_232),
.B(n_1),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_1),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g279 ( 
.A(n_201),
.B(n_33),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_201),
.B(n_2),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_199),
.B(n_3),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_221),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_205),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_205),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_227),
.B(n_35),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_199),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_4),
.Y(n_289)
);

AND2x6_ASAP7_75t_L g290 ( 
.A(n_219),
.B(n_36),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g291 ( 
.A(n_222),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_219),
.B(n_38),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_227),
.B(n_4),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_219),
.Y(n_296)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_259),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_203),
.B(n_5),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_252),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_5),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

BUFx8_ASAP7_75t_SL g305 ( 
.A(n_209),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_208),
.B(n_6),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_207),
.Y(n_307)
);

AND2x4_ASAP7_75t_L g308 ( 
.A(n_217),
.B(n_225),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_229),
.Y(n_309)
);

BUFx8_ASAP7_75t_SL g310 ( 
.A(n_220),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_236),
.B(n_6),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_244),
.B(n_7),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_226),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_208),
.B(n_7),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_238),
.B(n_8),
.Y(n_315)
);

CKINVDCx11_ASAP7_75t_R g316 ( 
.A(n_224),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_228),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_230),
.B(n_8),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_208),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_208),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_239),
.B(n_39),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_245),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_208),
.B(n_9),
.Y(n_324)
);

AO22x2_ASAP7_75t_L g325 ( 
.A1(n_275),
.A2(n_263),
.B1(n_262),
.B2(n_267),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_L g327 ( 
.A1(n_280),
.A2(n_300),
.B1(n_273),
.B2(n_276),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_313),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g329 ( 
.A1(n_273),
.A2(n_272),
.B1(n_248),
.B2(n_255),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_198),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_277),
.B(n_269),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_300),
.A2(n_271),
.B1(n_270),
.B2(n_268),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_283),
.B(n_200),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_202),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_281),
.Y(n_337)
);

OR2x6_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_254),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_312),
.A2(n_282),
.B1(n_292),
.B2(n_291),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_274),
.B(n_11),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

AO22x2_ASAP7_75t_L g344 ( 
.A1(n_275),
.A2(n_256),
.B1(n_265),
.B2(n_208),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_312),
.A2(n_266),
.B1(n_264),
.B2(n_260),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_292),
.A2(n_233),
.B1(n_251),
.B2(n_250),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_299),
.A2(n_257),
.B1(n_249),
.B2(n_247),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_286),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_274),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_299),
.A2(n_289),
.B1(n_301),
.B2(n_288),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_204),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_294),
.B(n_206),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_278),
.A2(n_246),
.B1(n_243),
.B2(n_240),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_276),
.B(n_210),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_306),
.A2(n_235),
.B1(n_234),
.B2(n_231),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_295),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_311),
.B(n_211),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_314),
.A2(n_223),
.B1(n_218),
.B2(n_215),
.Y(n_363)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_305),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_324),
.A2(n_214),
.B1(n_212),
.B2(n_13),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_288),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_315),
.B(n_40),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_295),
.Y(n_368)
);

AO22x2_ASAP7_75t_L g369 ( 
.A1(n_279),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_284),
.B(n_41),
.Y(n_370)
);

AO22x2_ASAP7_75t_L g371 ( 
.A1(n_279),
.A2(n_287),
.B1(n_318),
.B2(n_298),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_298),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_372)
);

AO22x2_ASAP7_75t_L g373 ( 
.A1(n_279),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_284),
.B(n_42),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_321),
.Y(n_375)
);

AND2x2_ASAP7_75t_SL g376 ( 
.A(n_287),
.B(n_20),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_321),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_318),
.B(n_22),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_328),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_329),
.B(n_310),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_343),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_356),
.Y(n_385)
);

OR2x6_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_287),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_321),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_359),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_354),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_351),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_313),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_355),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_326),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_326),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_332),
.B(n_317),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_337),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_337),
.Y(n_401)
);

INVxp33_ASAP7_75t_L g402 ( 
.A(n_378),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_340),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_340),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_346),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_349),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_361),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_361),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_362),
.B(n_307),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_341),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_329),
.B(n_310),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_364),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_335),
.B(n_309),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_338),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_364),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g420 ( 
.A(n_375),
.B(n_367),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_319),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_375),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_336),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

NAND2x1p5_ASAP7_75t_L g425 ( 
.A(n_376),
.B(n_284),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_353),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_347),
.B(n_316),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_325),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_348),
.B(n_316),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_357),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_357),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_325),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_339),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_334),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_338),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_344),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

INVxp33_ASAP7_75t_L g441 ( 
.A(n_345),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_SL g442 ( 
.A(n_372),
.B(n_369),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_344),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_377),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_374),
.B(n_319),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_R g447 ( 
.A(n_439),
.B(n_342),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_376),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_391),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_327),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_411),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_394),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_389),
.B(n_360),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_395),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_391),
.B(n_305),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_426),
.B(n_363),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_369),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_396),
.B(n_327),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_396),
.B(n_433),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_342),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_358),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_417),
.B(n_373),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_373),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_397),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_400),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_401),
.Y(n_468)
);

BUFx4f_ASAP7_75t_L g469 ( 
.A(n_425),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_366),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_365),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_317),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_412),
.B(n_373),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_429),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_422),
.B(n_338),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_317),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_435),
.B(n_444),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_317),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_388),
.B(n_322),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_388),
.B(n_322),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_414),
.B(n_369),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_437),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_399),
.B(n_352),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_399),
.B(n_322),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_427),
.B(n_421),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_421),
.B(n_322),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_420),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_425),
.B(n_420),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_404),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_441),
.B(n_284),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_406),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_434),
.B(n_445),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_416),
.Y(n_496)
);

INVx4_ASAP7_75t_L g497 ( 
.A(n_420),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_407),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_420),
.B(n_323),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_379),
.B(n_323),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_410),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_419),
.Y(n_503)
);

AND2x2_ASAP7_75t_SL g504 ( 
.A(n_398),
.B(n_323),
.Y(n_504)
);

AND2x2_ASAP7_75t_SL g505 ( 
.A(n_398),
.B(n_323),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_442),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_413),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_442),
.A2(n_290),
.B1(n_293),
.B2(n_304),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_380),
.B(n_290),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_381),
.B(n_382),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_423),
.B(n_296),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_390),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_403),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_398),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_384),
.B(n_290),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_438),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_461),
.B(n_441),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_448),
.B(n_488),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_466),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_466),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_514),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_466),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_488),
.B(n_385),
.Y(n_523)
);

CKINVDCx6p67_ASAP7_75t_R g524 ( 
.A(n_449),
.Y(n_524)
);

BUFx4f_ASAP7_75t_L g525 ( 
.A(n_495),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_477),
.B(n_386),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_456),
.Y(n_527)
);

OR2x6_ASAP7_75t_L g528 ( 
.A(n_482),
.B(n_489),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_487),
.B(n_403),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_497),
.B(n_403),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_477),
.B(n_386),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_487),
.B(n_409),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_474),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_450),
.B(n_409),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_452),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_482),
.B(n_393),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_514),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_459),
.B(n_402),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_477),
.B(n_386),
.Y(n_539)
);

BUFx2_ASAP7_75t_SL g540 ( 
.A(n_485),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_467),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_460),
.B(n_409),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_467),
.Y(n_543)
);

NAND2x1p5_ASAP7_75t_L g544 ( 
.A(n_497),
.B(n_387),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_485),
.B(n_290),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_506),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_514),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_467),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_497),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_456),
.B(n_293),
.Y(n_550)
);

NAND2x1_ASAP7_75t_SL g551 ( 
.A(n_508),
.B(n_383),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_483),
.B(n_402),
.Y(n_552)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_513),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_468),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_456),
.B(n_436),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_479),
.B(n_293),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_464),
.B(n_418),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_511),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_480),
.B(n_293),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_486),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_471),
.B(n_293),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_464),
.B(n_473),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_468),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_506),
.B(n_415),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_504),
.B(n_505),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_482),
.Y(n_566)
);

BUFx12f_ASAP7_75t_L g567 ( 
.A(n_475),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_452),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_504),
.B(n_296),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_491),
.Y(n_570)
);

NOR2x1_ASAP7_75t_L g571 ( 
.A(n_463),
.B(n_428),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_504),
.B(n_296),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_524),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_519),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_519),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_535),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_524),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_546),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_564),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_517),
.B(n_458),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_568),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_567),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_557),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

BUFx12f_ASAP7_75t_L g585 ( 
.A(n_555),
.Y(n_585)
);

AO22x2_ASAP7_75t_L g586 ( 
.A1(n_565),
.A2(n_518),
.B1(n_458),
.B2(n_465),
.Y(n_586)
);

CKINVDCx11_ASAP7_75t_R g587 ( 
.A(n_564),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_566),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_520),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_527),
.Y(n_590)
);

BUFx12f_ASAP7_75t_L g591 ( 
.A(n_555),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_534),
.B(n_473),
.Y(n_592)
);

INVx5_ASAP7_75t_SL g593 ( 
.A(n_528),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_527),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_540),
.B(n_562),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_538),
.A2(n_457),
.B1(n_495),
.B2(n_470),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_570),
.Y(n_597)
);

CKINVDCx6p67_ASAP7_75t_R g598 ( 
.A(n_567),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_558),
.B(n_529),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_522),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_555),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_522),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_541),
.Y(n_603)
);

INVx3_ASAP7_75t_SL g604 ( 
.A(n_564),
.Y(n_604)
);

BUFx2_ASAP7_75t_SL g605 ( 
.A(n_516),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_566),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_558),
.B(n_495),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_541),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_543),
.Y(n_609)
);

INVx8_ASAP7_75t_L g610 ( 
.A(n_528),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_528),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_516),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_543),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_566),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_532),
.B(n_495),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_552),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_548),
.Y(n_617)
);

NAND2x1p5_ASAP7_75t_L g618 ( 
.A(n_525),
.B(n_489),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_548),
.B(n_465),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_566),
.Y(n_620)
);

BUFx2_ASAP7_75t_L g621 ( 
.A(n_578),
.Y(n_621)
);

INVx6_ASAP7_75t_L g622 ( 
.A(n_585),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_619),
.B(n_495),
.Y(n_623)
);

CKINVDCx11_ASAP7_75t_R g624 ( 
.A(n_587),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_576),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_581),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_SL g627 ( 
.A1(n_616),
.A2(n_455),
.B1(n_484),
.B2(n_470),
.Y(n_627)
);

BUFx6f_ASAP7_75t_SL g628 ( 
.A(n_573),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_616),
.A2(n_484),
.B1(n_552),
.B2(n_470),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_596),
.A2(n_580),
.B1(n_525),
.B2(n_611),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_582),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_597),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_583),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_619),
.Y(n_634)
);

INVx6_ASAP7_75t_L g635 ( 
.A(n_585),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_574),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_592),
.A2(n_571),
.B1(n_470),
.B2(n_495),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_574),
.Y(n_638)
);

CKINVDCx11_ASAP7_75t_R g639 ( 
.A(n_587),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_583),
.A2(n_495),
.B1(n_470),
.B2(n_601),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_586),
.A2(n_470),
.B1(n_531),
.B2(n_526),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_603),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_608),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_588),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_586),
.A2(n_470),
.B1(n_526),
.B2(n_531),
.Y(n_645)
);

CKINVDCx8_ASAP7_75t_R g646 ( 
.A(n_582),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_611),
.A2(n_525),
.B1(n_469),
.B2(n_528),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_SL g648 ( 
.A1(n_579),
.A2(n_481),
.B1(n_469),
.B2(n_489),
.Y(n_648)
);

INVx6_ASAP7_75t_L g649 ( 
.A(n_591),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_579),
.Y(n_650)
);

INVx6_ASAP7_75t_L g651 ( 
.A(n_591),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_613),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_595),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_575),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_611),
.A2(n_469),
.B1(n_527),
.B2(n_531),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_573),
.A2(n_475),
.B1(n_496),
.B2(n_503),
.Y(n_656)
);

INVx6_ASAP7_75t_L g657 ( 
.A(n_577),
.Y(n_657)
);

INVx3_ASAP7_75t_SL g658 ( 
.A(n_598),
.Y(n_658)
);

BUFx4_ASAP7_75t_R g659 ( 
.A(n_577),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_612),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_612),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_586),
.A2(n_539),
.B1(n_526),
.B2(n_516),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_588),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_598),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_617),
.Y(n_665)
);

OAI222xp33_ASAP7_75t_L g666 ( 
.A1(n_629),
.A2(n_431),
.B1(n_599),
.B2(n_615),
.C1(n_607),
.C2(n_508),
.Y(n_666)
);

OAI222xp33_ASAP7_75t_L g667 ( 
.A1(n_627),
.A2(n_453),
.B1(n_542),
.B2(n_493),
.C1(n_523),
.C2(n_481),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_627),
.A2(n_586),
.B1(n_604),
.B2(n_539),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_653),
.A2(n_604),
.B1(n_539),
.B2(n_512),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_625),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_653),
.B(n_533),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_655),
.B(n_610),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_626),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_636),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_621),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_634),
.A2(n_512),
.B1(n_475),
.B2(n_563),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_SL g677 ( 
.A1(n_622),
.A2(n_610),
.B1(n_611),
.B2(n_593),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_648),
.A2(n_475),
.B1(n_563),
.B2(n_554),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_648),
.A2(n_611),
.B1(n_527),
.B2(n_593),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_638),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_637),
.A2(n_593),
.B1(n_605),
.B2(n_618),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_633),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_644),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_654),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_660),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_661),
.B(n_511),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_637),
.A2(n_593),
.B1(n_618),
.B2(n_490),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_632),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_642),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_643),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_641),
.A2(n_554),
.B1(n_610),
.B2(n_589),
.Y(n_691)
);

AOI222xp33_ASAP7_75t_L g692 ( 
.A1(n_624),
.A2(n_551),
.B1(n_561),
.B2(n_510),
.C1(n_498),
.C2(n_491),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_652),
.Y(n_693)
);

OAI22xp33_ASAP7_75t_L g694 ( 
.A1(n_622),
.A2(n_610),
.B1(n_497),
.B2(n_545),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_645),
.A2(n_600),
.B1(n_589),
.B2(n_609),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_665),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_SL g697 ( 
.A1(n_635),
.A2(n_649),
.B1(n_651),
.B2(n_650),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_635),
.A2(n_550),
.B1(n_590),
.B2(n_594),
.Y(n_698)
);

NAND2x1_ASAP7_75t_L g699 ( 
.A(n_655),
.B(n_588),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_639),
.Y(n_700)
);

BUFx12f_ASAP7_75t_L g701 ( 
.A(n_631),
.Y(n_701)
);

AOI222xp33_ASAP7_75t_L g702 ( 
.A1(n_623),
.A2(n_492),
.B1(n_498),
.B2(n_499),
.C1(n_584),
.C2(n_575),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_623),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_SL g704 ( 
.A1(n_649),
.A2(n_536),
.B1(n_614),
.B2(n_588),
.Y(n_704)
);

OAI222xp33_ASAP7_75t_L g705 ( 
.A1(n_640),
.A2(n_569),
.B1(n_572),
.B2(n_590),
.C1(n_594),
.C2(n_584),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_662),
.A2(n_609),
.B1(n_602),
.B2(n_600),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_656),
.A2(n_553),
.B1(n_549),
.B2(n_500),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_630),
.A2(n_549),
.B1(n_505),
.B2(n_620),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_630),
.A2(n_549),
.B1(n_505),
.B2(n_620),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_651),
.B(n_602),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_657),
.A2(n_620),
.B1(n_614),
.B2(n_588),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_628),
.A2(n_499),
.B1(n_492),
.B2(n_454),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_663),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_628),
.A2(n_647),
.B1(n_664),
.B2(n_454),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_669),
.A2(n_646),
.B1(n_657),
.B2(n_658),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_692),
.A2(n_647),
.B1(n_507),
.B2(n_502),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_668),
.A2(n_502),
.B1(n_507),
.B2(n_494),
.Y(n_717)
);

OAI222xp33_ASAP7_75t_L g718 ( 
.A1(n_668),
.A2(n_669),
.B1(n_678),
.B2(n_712),
.C1(n_714),
.C2(n_697),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_689),
.B(n_606),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_689),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_690),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_SL g722 ( 
.A1(n_679),
.A2(n_644),
.B1(n_659),
.B2(n_620),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_703),
.A2(n_502),
.B1(n_494),
.B2(n_507),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_703),
.A2(n_468),
.B1(n_494),
.B2(n_606),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_SL g725 ( 
.A1(n_681),
.A2(n_644),
.B1(n_620),
.B2(n_614),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_712),
.A2(n_714),
.B1(n_678),
.B2(n_691),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_675),
.A2(n_672),
.B1(n_686),
.B2(n_685),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_672),
.A2(n_606),
.B1(n_536),
.B2(n_614),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_672),
.A2(n_536),
.B1(n_614),
.B2(n_472),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_676),
.B(n_501),
.C(n_478),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_671),
.A2(n_559),
.B1(n_556),
.B2(n_544),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_691),
.A2(n_462),
.B1(n_544),
.B2(n_530),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_702),
.A2(n_536),
.B1(n_451),
.B2(n_476),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_676),
.A2(n_530),
.B1(n_560),
.B2(n_537),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_687),
.A2(n_682),
.B1(n_707),
.B2(n_713),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_SL g736 ( 
.A1(n_708),
.A2(n_536),
.B1(n_547),
.B2(n_537),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_701),
.A2(n_451),
.B1(n_509),
.B2(n_513),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_677),
.A2(n_513),
.B1(n_560),
.B2(n_537),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_690),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_SL g740 ( 
.A1(n_709),
.A2(n_547),
.B1(n_521),
.B2(n_560),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_710),
.A2(n_547),
.B1(n_521),
.B2(n_486),
.Y(n_741)
);

OAI222xp33_ASAP7_75t_L g742 ( 
.A1(n_704),
.A2(n_521),
.B1(n_320),
.B2(n_25),
.C1(n_26),
.C2(n_27),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_696),
.A2(n_486),
.B1(n_515),
.B2(n_320),
.Y(n_743)
);

OAI221xp5_ASAP7_75t_SL g744 ( 
.A1(n_698),
.A2(n_706),
.B1(n_673),
.B2(n_670),
.C(n_695),
.Y(n_744)
);

AOI222xp33_ASAP7_75t_L g745 ( 
.A1(n_666),
.A2(n_320),
.B1(n_447),
.B2(n_26),
.C1(n_28),
.C2(n_23),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_L g746 ( 
.A(n_667),
.B(n_486),
.C(n_447),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_706),
.A2(n_320),
.B1(n_303),
.B2(n_302),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_695),
.A2(n_303),
.B1(n_302),
.B2(n_297),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_SL g749 ( 
.A1(n_683),
.A2(n_304),
.B1(n_296),
.B2(n_30),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_694),
.A2(n_303),
.B(n_297),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_683),
.A2(n_304),
.B1(n_29),
.B2(n_30),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_696),
.A2(n_304),
.B1(n_303),
.B2(n_302),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_745),
.B(n_693),
.C(n_688),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_739),
.B(n_720),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_744),
.A2(n_699),
.B1(n_683),
.B2(n_680),
.Y(n_755)
);

OAI221xp5_ASAP7_75t_L g756 ( 
.A1(n_751),
.A2(n_700),
.B1(n_711),
.B2(n_684),
.C(n_674),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_735),
.B(n_674),
.C(n_683),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_739),
.B(n_24),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_720),
.B(n_24),
.Y(n_759)
);

OAI221xp5_ASAP7_75t_SL g760 ( 
.A1(n_749),
.A2(n_31),
.B1(n_705),
.B2(n_44),
.C(n_46),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_742),
.B(n_31),
.C(n_43),
.Y(n_761)
);

OA21x2_ASAP7_75t_L g762 ( 
.A1(n_750),
.A2(n_47),
.B(n_50),
.Y(n_762)
);

AOI221xp5_ASAP7_75t_L g763 ( 
.A1(n_718),
.A2(n_302),
.B1(n_297),
.B2(n_285),
.C(n_54),
.Y(n_763)
);

NAND3xp33_ASAP7_75t_L g764 ( 
.A(n_727),
.B(n_297),
.C(n_285),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_721),
.B(n_51),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_721),
.B(n_52),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_719),
.B(n_53),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_716),
.B(n_285),
.C(n_56),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_719),
.B(n_55),
.Y(n_769)
);

OA211x2_ASAP7_75t_L g770 ( 
.A1(n_729),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_715),
.B(n_61),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_722),
.B(n_285),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_726),
.B(n_62),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_725),
.B(n_63),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_728),
.B(n_64),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_717),
.B(n_740),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_746),
.B(n_196),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_731),
.B(n_66),
.Y(n_778)
);

OAI221xp5_ASAP7_75t_L g779 ( 
.A1(n_737),
.A2(n_67),
.B1(n_71),
.B2(n_72),
.C(n_76),
.Y(n_779)
);

OAI21xp33_ASAP7_75t_L g780 ( 
.A1(n_733),
.A2(n_77),
.B(n_79),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_730),
.B(n_80),
.Y(n_781)
);

OAI221xp5_ASAP7_75t_L g782 ( 
.A1(n_736),
.A2(n_738),
.B1(n_730),
.B2(n_724),
.C(n_741),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_763),
.B(n_747),
.C(n_748),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_761),
.A2(n_732),
.B1(n_723),
.B2(n_734),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_754),
.B(n_743),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_754),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_758),
.B(n_752),
.Y(n_787)
);

NAND3xp33_ASAP7_75t_L g788 ( 
.A(n_781),
.B(n_81),
.C(n_82),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_759),
.Y(n_789)
);

NAND4xp75_ASAP7_75t_L g790 ( 
.A(n_770),
.B(n_83),
.C(n_87),
.D(n_88),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_773),
.B(n_89),
.C(n_90),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_765),
.B(n_92),
.Y(n_792)
);

OAI21xp33_ASAP7_75t_SL g793 ( 
.A1(n_772),
.A2(n_94),
.B(n_95),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_766),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_777),
.B(n_96),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_777),
.B(n_97),
.Y(n_796)
);

NOR2x1_ASAP7_75t_L g797 ( 
.A(n_757),
.B(n_98),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_753),
.B(n_100),
.C(n_101),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_771),
.B(n_102),
.C(n_103),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_789),
.B(n_756),
.Y(n_800)
);

NAND4xp75_ASAP7_75t_SL g801 ( 
.A(n_795),
.B(n_762),
.C(n_775),
.D(n_760),
.Y(n_801)
);

XNOR2x2_ASAP7_75t_L g802 ( 
.A(n_798),
.B(n_764),
.Y(n_802)
);

NAND4xp75_ASAP7_75t_L g803 ( 
.A(n_797),
.B(n_793),
.C(n_762),
.D(n_796),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_786),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_789),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_SL g806 ( 
.A(n_790),
.B(n_799),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_794),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_794),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_785),
.B(n_788),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_787),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_805),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_806),
.A2(n_755),
.B1(n_791),
.B2(n_783),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_804),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_810),
.B(n_792),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_807),
.Y(n_815)
);

XOR2x2_ASAP7_75t_L g816 ( 
.A(n_812),
.B(n_800),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_813),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_811),
.Y(n_818)
);

OA22x2_ASAP7_75t_L g819 ( 
.A1(n_814),
.A2(n_809),
.B1(n_808),
.B2(n_784),
.Y(n_819)
);

INVx3_ASAP7_75t_SL g820 ( 
.A(n_814),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_817),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_820),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_817),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_818),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_822),
.A2(n_816),
.B1(n_819),
.B2(n_809),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_824),
.Y(n_826)
);

OAI322xp33_ASAP7_75t_L g827 ( 
.A1(n_821),
.A2(n_802),
.A3(n_815),
.B1(n_755),
.B2(n_774),
.C1(n_778),
.C2(n_801),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_827),
.A2(n_824),
.B(n_823),
.C(n_783),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_825),
.A2(n_803),
.B1(n_780),
.B2(n_779),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_826),
.A2(n_803),
.B1(n_769),
.B2(n_767),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_826),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_831),
.Y(n_832)
);

AO22x2_ASAP7_75t_L g833 ( 
.A1(n_828),
.A2(n_802),
.B1(n_768),
.B2(n_776),
.Y(n_833)
);

AO22x2_ASAP7_75t_L g834 ( 
.A1(n_829),
.A2(n_782),
.B1(n_105),
.B2(n_106),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_830),
.B(n_104),
.Y(n_835)
);

AOI22xp5_ASAP7_75t_L g836 ( 
.A1(n_829),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_831),
.B(n_112),
.Y(n_837)
);

NAND4xp25_ASAP7_75t_L g838 ( 
.A(n_828),
.B(n_113),
.C(n_114),
.D(n_116),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_832),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_833),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_837),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_835),
.Y(n_842)
);

NOR3xp33_ASAP7_75t_L g843 ( 
.A(n_838),
.B(n_122),
.C(n_123),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_836),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_834),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_832),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_839),
.Y(n_847)
);

NAND5xp2_ASAP7_75t_L g848 ( 
.A(n_845),
.B(n_124),
.C(n_125),
.D(n_126),
.E(n_127),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_L g849 ( 
.A(n_842),
.B(n_129),
.C(n_130),
.Y(n_849)
);

NOR2x1_ASAP7_75t_L g850 ( 
.A(n_846),
.B(n_131),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_841),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_844),
.Y(n_852)
);

NOR2xp67_ASAP7_75t_L g853 ( 
.A(n_840),
.B(n_191),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_843),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_854)
);

AND4x1_ASAP7_75t_L g855 ( 
.A(n_843),
.B(n_138),
.C(n_142),
.D(n_143),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_847),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_852),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_850),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_851),
.Y(n_859)
);

INVxp67_ASAP7_75t_SL g860 ( 
.A(n_853),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_854),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_848),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_855),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_863),
.A2(n_862),
.B1(n_861),
.B2(n_857),
.Y(n_864)
);

BUFx8_ASAP7_75t_L g865 ( 
.A(n_859),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_860),
.A2(n_858),
.B1(n_856),
.B2(n_849),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_856),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_867)
);

AO22x2_ASAP7_75t_L g868 ( 
.A1(n_856),
.A2(n_190),
.B1(n_149),
.B2(n_150),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_862),
.A2(n_148),
.B1(n_151),
.B2(n_153),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_862),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_865),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_866),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_868),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_871),
.A2(n_864),
.B1(n_869),
.B2(n_870),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_872),
.A2(n_867),
.B1(n_158),
.B2(n_159),
.Y(n_875)
);

AOI221xp5_ASAP7_75t_L g876 ( 
.A1(n_873),
.A2(n_157),
.B1(n_161),
.B2(n_165),
.C(n_170),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_875),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_877),
.A2(n_874),
.B1(n_876),
.B2(n_173),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_878),
.Y(n_879)
);

AOI221xp5_ASAP7_75t_L g880 ( 
.A1(n_879),
.A2(n_171),
.B1(n_172),
.B2(n_175),
.C(n_176),
.Y(n_880)
);

AOI211xp5_ASAP7_75t_L g881 ( 
.A1(n_880),
.A2(n_180),
.B(n_181),
.C(n_185),
.Y(n_881)
);


endmodule