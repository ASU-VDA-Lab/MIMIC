module real_aes_294_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_668;
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_0), .A2(n_148), .B1(n_426), .B2(n_427), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_1), .A2(n_48), .B1(n_371), .B2(n_555), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_2), .B(n_288), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_3), .A2(n_108), .B1(n_434), .B2(n_454), .Y(n_562) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_4), .A2(n_9), .B1(n_548), .B2(n_584), .Y(n_583) );
AO22x2_ASAP7_75t_L g304 ( .A1(n_5), .A2(n_206), .B1(n_294), .B2(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g740 ( .A(n_5), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_6), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_7), .A2(n_173), .B1(n_336), .B2(n_352), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_8), .A2(n_19), .B1(n_660), .B2(n_661), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_10), .A2(n_52), .B1(n_375), .B2(n_377), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_11), .A2(n_132), .B1(n_359), .B2(n_379), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_12), .A2(n_75), .B1(n_391), .B2(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_13), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_14), .A2(n_254), .B1(n_370), .B2(n_371), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_15), .A2(n_142), .B1(n_436), .B2(n_437), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g417 ( .A1(n_16), .A2(n_248), .B1(n_418), .B2(n_419), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_17), .A2(n_157), .B1(n_339), .B2(n_344), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_18), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_20), .A2(n_47), .B1(n_494), .B2(n_661), .Y(n_783) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_21), .A2(n_73), .B1(n_294), .B2(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_21), .B(n_739), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_22), .A2(n_135), .B1(n_390), .B2(n_586), .Y(n_585) );
AO222x2_ASAP7_75t_L g701 ( .A1(n_23), .A2(n_72), .B1(n_224), .B2(n_413), .C1(n_419), .C2(n_527), .Y(n_701) );
XOR2x2_ASAP7_75t_L g767 ( .A(n_24), .B(n_768), .Y(n_767) );
INVxp67_ASAP7_75t_L g792 ( .A(n_24), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_25), .A2(n_158), .B1(n_317), .B2(n_321), .Y(n_316) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_26), .A2(n_225), .B1(n_426), .B2(n_427), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_27), .A2(n_251), .B1(n_429), .B2(n_430), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_28), .A2(n_152), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_29), .A2(n_197), .B1(n_359), .B2(n_558), .Y(n_557) );
AOI222xp33_ASAP7_75t_L g685 ( .A1(n_30), .A2(n_65), .B1(n_162), .B2(n_413), .C1(n_414), .C2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_31), .A2(n_59), .B1(n_330), .B2(n_475), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_32), .A2(n_231), .B1(n_478), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_33), .A2(n_37), .B1(n_436), .B2(n_437), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_34), .A2(n_50), .B1(n_344), .B2(n_347), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_35), .A2(n_223), .B1(n_350), .B2(n_352), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_36), .A2(n_221), .B1(n_383), .B2(n_384), .Y(n_382) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_38), .A2(n_235), .B1(n_415), .B2(n_523), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_39), .A2(n_262), .B1(n_669), .B2(n_771), .Y(n_770) );
AOI222xp33_ASAP7_75t_L g479 ( .A1(n_40), .A2(n_171), .B1(n_237), .B2(n_321), .C1(n_480), .C2(n_481), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_41), .A2(n_130), .B1(n_436), .B2(n_437), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_42), .A2(n_220), .B1(n_475), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_43), .A2(n_116), .B1(n_434), .B2(n_454), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_44), .Y(n_636) );
OA22x2_ASAP7_75t_L g605 ( .A1(n_45), .A2(n_606), .B1(n_607), .B2(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_45), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_46), .A2(n_242), .B1(n_348), .B2(n_350), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_49), .A2(n_193), .B1(n_418), .B2(n_419), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_51), .A2(n_136), .B1(n_326), .B2(n_548), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_53), .A2(n_138), .B1(n_355), .B2(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_54), .A2(n_177), .B1(n_355), .B2(n_357), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_55), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_56), .A2(n_166), .B1(n_307), .B2(n_312), .Y(n_306) );
AOI22xp33_ASAP7_75t_SL g703 ( .A1(n_57), .A2(n_118), .B1(n_418), .B2(n_421), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_58), .A2(n_99), .B1(n_497), .B2(n_727), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_60), .A2(n_263), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_61), .A2(n_154), .B1(n_399), .B2(n_402), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_62), .A2(n_264), .B1(n_399), .B2(n_402), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_63), .A2(n_255), .B1(n_321), .B2(n_544), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_64), .A2(n_284), .B1(n_285), .B2(n_361), .Y(n_283) );
INVxp67_ASAP7_75t_L g361 ( .A(n_64), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_66), .A2(n_194), .B1(n_580), .B2(n_752), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_67), .A2(n_258), .B1(n_379), .B2(n_591), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_68), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_69), .B(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_70), .A2(n_187), .B1(n_352), .B2(n_561), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_71), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_74), .A2(n_145), .B1(n_336), .B2(n_465), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_76), .A2(n_128), .B1(n_493), .B2(n_494), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_77), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_78), .A2(n_180), .B1(n_429), .B2(n_436), .Y(n_708) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_79), .A2(n_236), .B1(n_426), .B2(n_427), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_80), .A2(n_243), .B1(n_430), .B2(n_434), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_81), .A2(n_200), .B1(n_497), .B2(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g596 ( .A(n_82), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_83), .A2(n_131), .B1(n_421), .B2(n_422), .Y(n_445) );
OAI22x1_ASAP7_75t_L g671 ( .A1(n_84), .A2(n_672), .B1(n_687), .B2(n_688), .Y(n_671) );
CKINVDCx16_ASAP7_75t_R g688 ( .A(n_84), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_85), .A2(n_149), .B1(n_384), .B2(n_773), .Y(n_772) );
INVx3_ASAP7_75t_L g294 ( .A(n_86), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_87), .A2(n_164), .B1(n_433), .B2(n_437), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_88), .A2(n_170), .B1(n_307), .B2(n_586), .Y(n_656) );
AO21x2_ASAP7_75t_L g364 ( .A1(n_89), .A2(n_365), .B(n_404), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_89), .B(n_367), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_90), .A2(n_94), .B1(n_393), .B2(n_395), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_91), .A2(n_133), .B1(n_433), .B2(n_434), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_92), .A2(n_210), .B1(n_465), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_93), .A2(n_244), .B1(n_781), .B2(n_782), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_95), .A2(n_199), .B1(n_476), .B2(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_96), .A2(n_189), .B1(n_475), .B2(n_548), .Y(n_674) );
OA22x2_ASAP7_75t_L g485 ( .A1(n_97), .A2(n_486), .B1(n_487), .B2(n_508), .Y(n_485) );
INVxp67_ASAP7_75t_L g508 ( .A(n_97), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_98), .A2(n_253), .B1(n_755), .B2(n_756), .Y(n_754) );
XOR2x2_ASAP7_75t_L g714 ( .A(n_100), .B(n_715), .Y(n_714) );
AO222x2_ASAP7_75t_L g412 ( .A1(n_101), .A2(n_155), .B1(n_179), .B2(n_413), .C1(n_414), .C2(n_415), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_102), .A2(n_122), .B1(n_777), .B2(n_778), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_103), .A2(n_208), .B1(n_376), .B2(n_491), .Y(n_589) );
INVx1_ASAP7_75t_L g483 ( .A(n_104), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_105), .A2(n_190), .B1(n_427), .B2(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_106), .A2(n_159), .B1(n_421), .B2(n_422), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_107), .Y(n_619) );
INVx1_ASAP7_75t_SL g295 ( .A(n_109), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_109), .B(n_143), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_110), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g784 ( .A1(n_111), .A2(n_123), .B1(n_239), .B2(n_393), .C1(n_395), .C2(n_480), .Y(n_784) );
INVx2_ASAP7_75t_L g276 ( .A(n_112), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_113), .A2(n_192), .B1(n_339), .B2(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_114), .A2(n_184), .B1(n_494), .B2(n_679), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_115), .A2(n_249), .B1(n_433), .B2(n_434), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_117), .A2(n_234), .B1(n_663), .B2(n_664), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_119), .A2(n_181), .B1(n_336), .B2(n_339), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_120), .A2(n_245), .B1(n_504), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_121), .A2(n_265), .B1(n_627), .B2(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_124), .A2(n_202), .B1(n_470), .B2(n_472), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_125), .A2(n_156), .B1(n_393), .B2(n_395), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_126), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_127), .B(n_288), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_129), .A2(n_172), .B1(n_348), .B2(n_497), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_134), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_137), .A2(n_151), .B1(n_336), .B2(n_664), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_139), .A2(n_744), .B1(n_745), .B2(n_763), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_139), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_140), .A2(n_268), .B1(n_529), .B2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_141), .A2(n_146), .B1(n_344), .B2(n_491), .Y(n_490) );
AO22x2_ASAP7_75t_L g297 ( .A1(n_143), .A2(n_214), .B1(n_294), .B2(n_298), .Y(n_297) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_144), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_147), .A2(n_163), .B1(n_330), .B2(n_475), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_150), .A2(n_247), .B1(n_344), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_153), .A2(n_174), .B1(n_491), .B2(n_623), .Y(n_758) );
INVx1_ASAP7_75t_L g296 ( .A(n_160), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_161), .A2(n_230), .B1(n_414), .B2(n_415), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_165), .A2(n_169), .B1(n_357), .B2(n_760), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_167), .A2(n_185), .B1(n_429), .B2(n_430), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_168), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_175), .A2(n_211), .B1(n_355), .B2(n_357), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_176), .A2(n_218), .B1(n_307), .B2(n_504), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_178), .A2(n_238), .B1(n_389), .B2(n_391), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_182), .A2(n_196), .B1(n_317), .B2(n_506), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_183), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_186), .A2(n_209), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_188), .A2(n_256), .B1(n_307), .B2(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_191), .A2(n_232), .B1(n_373), .B2(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_195), .B(n_387), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_198), .A2(n_219), .B1(n_419), .B2(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_201), .A2(n_217), .B1(n_326), .B2(n_330), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_203), .B(n_288), .Y(n_287) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_204), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_205), .A2(n_266), .B1(n_383), .B2(n_727), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_207), .A2(n_226), .B1(n_534), .B2(n_594), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_212), .A2(n_267), .B1(n_352), .B2(n_561), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_213), .A2(n_698), .B1(n_699), .B2(n_712), .Y(n_697) );
INVx1_ASAP7_75t_L g712 ( .A(n_213), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_215), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_216), .A2(n_260), .B1(n_415), .B2(n_523), .Y(n_522) );
AND2x4_ASAP7_75t_L g278 ( .A(n_222), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g736 ( .A(n_222), .Y(n_736) );
AO21x1_ASAP7_75t_L g790 ( .A1(n_222), .A2(n_274), .B(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_227), .A2(n_259), .B1(n_389), .B2(n_391), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_228), .A2(n_271), .B(n_280), .C(n_742), .Y(n_270) );
INVx1_ASAP7_75t_L g279 ( .A(n_229), .Y(n_279) );
AND2x2_ASAP7_75t_R g765 ( .A(n_229), .B(n_736), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_233), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_240), .A2(n_257), .B1(n_317), .B2(n_321), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_241), .A2(n_269), .B1(n_317), .B2(n_321), .Y(n_719) );
INVxp67_ASAP7_75t_L g275 ( .A(n_246), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_250), .B(n_413), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_252), .B(n_387), .Y(n_386) );
AOI22x1_ASAP7_75t_L g646 ( .A1(n_261), .A2(n_647), .B1(n_648), .B2(n_670), .Y(n_646) );
INVx1_ASAP7_75t_L g670 ( .A(n_261), .Y(n_670) );
XNOR2x1_ASAP7_75t_L g691 ( .A(n_261), .B(n_648), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_279), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g791 ( .A(n_279), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_511), .B1(n_731), .B2(n_732), .C(n_733), .Y(n_280) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_281), .Y(n_731) );
XNOR2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_362), .Y(n_281) );
HB1xp67_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp67_ASAP7_75t_L g285 ( .A(n_286), .B(n_334), .Y(n_285) );
NAND4xp25_ASAP7_75t_L g286 ( .A(n_287), .B(n_306), .C(n_316), .D(n_325), .Y(n_286) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_288), .Y(n_748) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g387 ( .A(n_289), .Y(n_387) );
INVx4_ASAP7_75t_SL g480 ( .A(n_289), .Y(n_480) );
INVx4_ASAP7_75t_SL g521 ( .A(n_289), .Y(n_521) );
INVx3_ASAP7_75t_SL g577 ( .A(n_289), .Y(n_577) );
INVx6_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_299), .Y(n_290) );
AND2x4_ASAP7_75t_L g314 ( .A(n_291), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g331 ( .A(n_291), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g413 ( .A(n_291), .B(n_299), .Y(n_413) );
AND2x2_ASAP7_75t_L g419 ( .A(n_291), .B(n_315), .Y(n_419) );
AND2x2_ASAP7_75t_L g422 ( .A(n_291), .B(n_332), .Y(n_422) );
AND2x2_ASAP7_75t_L g527 ( .A(n_291), .B(n_332), .Y(n_527) );
AND2x2_ASAP7_75t_L g676 ( .A(n_291), .B(n_315), .Y(n_676) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_297), .Y(n_291) );
INVx2_ASAP7_75t_L g311 ( .A(n_292), .Y(n_311) );
AND2x2_ASAP7_75t_L g319 ( .A(n_292), .B(n_320), .Y(n_319) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_292), .Y(n_324) );
OAI22x1_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B1(n_295), .B2(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g298 ( .A(n_294), .Y(n_298) );
INVx2_ASAP7_75t_L g302 ( .A(n_294), .Y(n_302) );
INVx1_ASAP7_75t_L g305 ( .A(n_294), .Y(n_305) );
AND2x2_ASAP7_75t_L g310 ( .A(n_297), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g320 ( .A(n_297), .Y(n_320) );
BUFx2_ASAP7_75t_L g360 ( .A(n_297), .Y(n_360) );
AND2x2_ASAP7_75t_L g338 ( .A(n_299), .B(n_310), .Y(n_338) );
AND2x4_ASAP7_75t_L g346 ( .A(n_299), .B(n_342), .Y(n_346) );
AND2x4_ASAP7_75t_L g351 ( .A(n_299), .B(n_319), .Y(n_351) );
AND2x2_ASAP7_75t_L g429 ( .A(n_299), .B(n_342), .Y(n_429) );
AND2x2_ASAP7_75t_L g433 ( .A(n_299), .B(n_319), .Y(n_433) );
AND2x6_ASAP7_75t_L g436 ( .A(n_299), .B(n_310), .Y(n_436) );
AND2x2_ASAP7_75t_L g454 ( .A(n_299), .B(n_319), .Y(n_454) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x4_ASAP7_75t_L g309 ( .A(n_301), .B(n_303), .Y(n_309) );
AND2x2_ASAP7_75t_L g323 ( .A(n_301), .B(n_304), .Y(n_323) );
INVx1_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
INVxp67_ASAP7_75t_L g315 ( .A(n_303), .Y(n_315) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g328 ( .A(n_304), .B(n_329), .Y(n_328) );
BUFx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_308), .Y(n_390) );
BUFx2_ASAP7_75t_L g478 ( .A(n_308), .Y(n_478) );
BUFx2_ASAP7_75t_L g750 ( .A(n_308), .Y(n_750) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g318 ( .A(n_309), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g353 ( .A(n_309), .B(n_342), .Y(n_353) );
AND2x4_ASAP7_75t_L g415 ( .A(n_309), .B(n_319), .Y(n_415) );
AND2x2_ASAP7_75t_L g418 ( .A(n_309), .B(n_310), .Y(n_418) );
AND2x2_ASAP7_75t_L g430 ( .A(n_309), .B(n_342), .Y(n_430) );
AND2x2_ASAP7_75t_L g529 ( .A(n_309), .B(n_310), .Y(n_529) );
AND2x2_ASAP7_75t_L g356 ( .A(n_310), .B(n_328), .Y(n_356) );
AND2x2_ASAP7_75t_SL g426 ( .A(n_310), .B(n_328), .Y(n_426) );
AND2x2_ASAP7_75t_L g450 ( .A(n_310), .B(n_328), .Y(n_450) );
AND2x4_ASAP7_75t_L g342 ( .A(n_311), .B(n_320), .Y(n_342) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g391 ( .A(n_313), .Y(n_391) );
INVx1_ASAP7_75t_L g504 ( .A(n_313), .Y(n_504) );
INVx2_ASAP7_75t_L g551 ( .A(n_313), .Y(n_551) );
INVx2_ASAP7_75t_SL g586 ( .A(n_313), .Y(n_586) );
INVx2_ASAP7_75t_SL g778 ( .A(n_313), .Y(n_778) );
INVx6_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx5_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx3_ASAP7_75t_L g394 ( .A(n_318), .Y(n_394) );
INVx2_ASAP7_75t_L g482 ( .A(n_318), .Y(n_482) );
BUFx3_ASAP7_75t_L g753 ( .A(n_318), .Y(n_753) );
AND2x2_ASAP7_75t_L g327 ( .A(n_319), .B(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g421 ( .A(n_319), .B(n_328), .Y(n_421) );
BUFx3_ASAP7_75t_L g580 ( .A(n_321), .Y(n_580) );
BUFx12f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx3_ASAP7_75t_L g397 ( .A(n_322), .Y(n_397) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x4_ASAP7_75t_L g348 ( .A(n_323), .B(n_342), .Y(n_348) );
AND2x4_ASAP7_75t_L g359 ( .A(n_323), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_SL g414 ( .A(n_323), .B(n_324), .Y(n_414) );
AND2x4_ASAP7_75t_L g427 ( .A(n_323), .B(n_360), .Y(n_427) );
AND2x4_ASAP7_75t_L g434 ( .A(n_323), .B(n_342), .Y(n_434) );
AND2x2_ASAP7_75t_SL g523 ( .A(n_323), .B(n_324), .Y(n_523) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_326), .Y(n_755) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx3_ASAP7_75t_L g401 ( .A(n_327), .Y(n_401) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_327), .Y(n_475) );
AND2x4_ASAP7_75t_L g341 ( .A(n_328), .B(n_342), .Y(n_341) );
AND2x6_ASAP7_75t_L g437 ( .A(n_328), .B(n_342), .Y(n_437) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_329), .Y(n_333) );
BUFx4f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx3_ASAP7_75t_L g403 ( .A(n_331), .Y(n_403) );
BUFx6f_ASAP7_75t_SL g476 ( .A(n_331), .Y(n_476) );
INVx2_ASAP7_75t_L g549 ( .A(n_331), .Y(n_549) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND4xp25_ASAP7_75t_L g334 ( .A(n_335), .B(n_343), .C(n_349), .D(n_354), .Y(n_334) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx3_ASAP7_75t_L g555 ( .A(n_337), .Y(n_555) );
INVx2_ASAP7_75t_L g632 ( .A(n_337), .Y(n_632) );
INVx2_ASAP7_75t_SL g663 ( .A(n_337), .Y(n_663) );
INVx2_ASAP7_75t_SL g781 ( .A(n_337), .Y(n_781) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g376 ( .A(n_338), .Y(n_376) );
BUFx2_ASAP7_75t_L g681 ( .A(n_338), .Y(n_681) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g377 ( .A(n_340), .Y(n_377) );
INVx2_ASAP7_75t_L g491 ( .A(n_340), .Y(n_491) );
INVx2_ASAP7_75t_SL g556 ( .A(n_340), .Y(n_556) );
INVx2_ASAP7_75t_L g635 ( .A(n_340), .Y(n_635) );
INVx2_ASAP7_75t_SL g664 ( .A(n_340), .Y(n_664) );
INVx1_ASAP7_75t_SL g782 ( .A(n_340), .Y(n_782) );
INVx8_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx4_ASAP7_75t_L g370 ( .A(n_345), .Y(n_370) );
INVx3_ASAP7_75t_SL g534 ( .A(n_345), .Y(n_534) );
INVx2_ASAP7_75t_L g561 ( .A(n_345), .Y(n_561) );
INVx2_ASAP7_75t_SL g624 ( .A(n_345), .Y(n_624) );
INVx8_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_SL g384 ( .A(n_348), .Y(n_384) );
BUFx3_ASAP7_75t_L g472 ( .A(n_348), .Y(n_472) );
INVx2_ASAP7_75t_L g499 ( .A(n_348), .Y(n_499) );
BUFx2_ASAP7_75t_SL g627 ( .A(n_348), .Y(n_627) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g383 ( .A(n_351), .Y(n_383) );
INVx6_ASAP7_75t_L g471 ( .A(n_351), .Y(n_471) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_352), .Y(n_594) );
INVx1_ASAP7_75t_L g725 ( .A(n_352), .Y(n_725) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_353), .Y(n_373) );
BUFx3_ASAP7_75t_L g465 ( .A(n_353), .Y(n_465) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
BUFx3_ASAP7_75t_L g558 ( .A(n_356), .Y(n_558) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI22xp33_ASAP7_75t_SL g637 ( .A1(n_358), .A2(n_638), .B1(n_641), .B2(n_642), .Y(n_637) );
INVx3_ASAP7_75t_L g661 ( .A(n_358), .Y(n_661) );
INVx5_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g493 ( .A(n_359), .Y(n_493) );
BUFx3_ASAP7_75t_L g591 ( .A(n_359), .Y(n_591) );
BUFx2_ASAP7_75t_L g679 ( .A(n_359), .Y(n_679) );
XNOR2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_405), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_385), .Y(n_367) );
NAND4xp25_ASAP7_75t_SL g368 ( .A(n_369), .B(n_374), .C(n_378), .D(n_382), .Y(n_368) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_370), .Y(n_669) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g617 ( .A1(n_372), .A2(n_471), .B1(n_618), .B2(n_619), .Y(n_617) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_373), .Y(n_771) );
BUFx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g495 ( .A(n_381), .Y(n_495) );
NAND4xp25_ASAP7_75t_SL g385 ( .A(n_386), .B(n_388), .C(n_392), .D(n_398), .Y(n_385) );
BUFx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx4f_ASAP7_75t_SL g777 ( .A(n_390), .Y(n_777) );
BUFx6f_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g506 ( .A(n_397), .Y(n_506) );
BUFx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g502 ( .A(n_401), .Y(n_502) );
INVx4_ASAP7_75t_L g526 ( .A(n_401), .Y(n_526) );
BUFx6f_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_459), .B1(n_509), .B2(n_510), .Y(n_405) );
INVx1_ASAP7_75t_L g509 ( .A(n_406), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_438), .B1(n_457), .B2(n_458), .Y(n_406) );
INVx1_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
XNOR2x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_423), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .Y(n_411) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_415), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_431), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g458 ( .A(n_438), .Y(n_458) );
XOR2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_456), .Y(n_438) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_440), .B(n_447), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_444), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_451), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
INVx2_ASAP7_75t_SL g510 ( .A(n_459), .Y(n_510) );
OA22x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_484), .B2(n_485), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
XOR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_483), .Y(n_461) );
NAND4xp75_ASAP7_75t_L g462 ( .A(n_463), .B(n_467), .C(n_473), .D(n_479), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx3_ASAP7_75t_L g497 ( .A(n_471), .Y(n_497) );
INVx2_ASAP7_75t_L g667 ( .A(n_471), .Y(n_667) );
INVx2_ASAP7_75t_L g773 ( .A(n_471), .Y(n_773) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_477), .Y(n_473) );
BUFx6f_ASAP7_75t_SL g584 ( .A(n_475), .Y(n_584) );
BUFx2_ASAP7_75t_SL g756 ( .A(n_476), .Y(n_756) );
INVx1_ASAP7_75t_L g651 ( .A(n_480), .Y(n_651) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g544 ( .A(n_482), .Y(n_544) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
NOR2x1_ASAP7_75t_L g487 ( .A(n_488), .B(n_500), .Y(n_487) );
NAND4xp25_ASAP7_75t_SL g488 ( .A(n_489), .B(n_490), .C(n_492), .D(n_496), .Y(n_488) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g640 ( .A(n_495), .Y(n_640) );
INVx2_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g727 ( .A(n_499), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .C(n_505), .D(n_507), .Y(n_500) );
INVx1_ASAP7_75t_L g732 ( .A(n_511), .Y(n_732) );
XNOR2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_600), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OAI22xp33_ASAP7_75t_R g513 ( .A1(n_514), .A2(n_515), .B1(n_566), .B2(n_567), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AO22x2_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_539), .B1(n_564), .B2(n_565), .Y(n_515) );
INVx1_ASAP7_75t_SL g565 ( .A(n_516), .Y(n_565) );
INVx1_ASAP7_75t_L g598 ( .A(n_516), .Y(n_598) );
XOR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_538), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_518), .B(n_530), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_524), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g564 ( .A(n_539), .Y(n_564) );
XOR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_563), .Y(n_539) );
NAND2x1p5_ASAP7_75t_L g540 ( .A(n_541), .B(n_552), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_544), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .Y(n_546) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NOR2x1_ASAP7_75t_L g552 ( .A(n_553), .B(n_559), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
BUFx2_ASAP7_75t_L g760 ( .A(n_558), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_597), .B1(n_598), .B2(n_599), .Y(n_567) );
INVx3_ASAP7_75t_L g599 ( .A(n_568), .Y(n_599) );
XOR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_596), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_570), .B(n_587), .Y(n_569) );
NOR2x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_582), .Y(n_570) );
OAI222xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B1(n_575), .B2(n_578), .C1(n_579), .C2(n_581), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g610 ( .A1(n_575), .A2(n_611), .B(n_612), .Y(n_610) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_592), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_694), .B2(n_730), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_643), .B1(n_644), .B2(n_692), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_605), .Y(n_693) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND3x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_616), .C(n_628), .Y(n_608) );
NOR2xp67_ASAP7_75t_SL g609 ( .A(n_610), .B(n_613), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_614), .B(n_615), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_625), .B2(n_626), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_637), .Y(n_628) );
OAI22xp33_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_633), .B1(n_634), .B2(n_636), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g660 ( .A(n_640), .Y(n_660) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AO22x2_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_671), .B1(n_689), .B2(n_690), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_657), .Y(n_648) );
NOR2xp67_ASAP7_75t_L g649 ( .A(n_650), .B(n_654), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B(n_653), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
NOR2x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_665), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVx2_ASAP7_75t_L g689 ( .A(n_671), .Y(n_689) );
NAND4xp25_ASAP7_75t_SL g672 ( .A(n_673), .B(n_677), .C(n_682), .D(n_685), .Y(n_672) );
AND4x1_ASAP7_75t_L g687 ( .A(n_673), .B(n_677), .C(n_682), .D(n_685), .Y(n_687) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g730 ( .A(n_695), .Y(n_730) );
AO22x2_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_713), .B1(n_714), .B2(n_729), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
BUFx2_ASAP7_75t_L g729 ( .A(n_697), .Y(n_729) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_700), .B(n_705), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_709), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR2xp67_ASAP7_75t_L g715 ( .A(n_716), .B(n_721), .Y(n_715) );
NAND4xp25_ASAP7_75t_SL g716 ( .A(n_717), .B(n_718), .C(n_719), .D(n_720), .Y(n_716) );
NAND4xp25_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .C(n_726), .D(n_728), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_737), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_735), .B(n_738), .Y(n_787) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
OAI222xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_764), .B1(n_766), .B2(n_785), .C1(n_788), .C2(n_792), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_757), .Y(n_745) );
NAND4xp25_ASAP7_75t_SL g746 ( .A(n_747), .B(n_749), .C(n_751), .D(n_754), .Y(n_746) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
NAND4xp25_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .C(n_761), .D(n_762), .Y(n_757) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
NAND4xp75_ASAP7_75t_SL g768 ( .A(n_769), .B(n_774), .C(n_779), .D(n_784), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
AND2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_783), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
CKINVDCx6p67_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
endmodule