module fake_jpeg_28541_n_377 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_377);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_377;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_27),
.Y(n_45)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_9),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_63),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_9),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx4f_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_8),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_35),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_39),
.B1(n_29),
.B2(n_36),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_83),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_74),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_107),
.B1(n_65),
.B2(n_51),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_36),
.B(n_35),
.C(n_43),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_87),
.B(n_0),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_93),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_96),
.B1(n_118),
.B2(n_52),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_44),
.A2(n_27),
.B1(n_29),
.B2(n_39),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_109),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_23),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_48),
.A2(n_34),
.B1(n_36),
.B2(n_43),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_58),
.A2(n_34),
.B1(n_18),
.B2(n_28),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_122),
.B1(n_95),
.B2(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_30),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_19),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_46),
.A2(n_69),
.B1(n_56),
.B2(n_62),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_21),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_124),
.B(n_128),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_30),
.B(n_23),
.C(n_26),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_126),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_127),
.A2(n_136),
.B1(n_146),
.B2(n_161),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_21),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_82),
.A2(n_57),
.B1(n_60),
.B2(n_112),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_129),
.A2(n_132),
.B1(n_158),
.B2(n_98),
.Y(n_172)
);

AOI32xp33_ASAP7_75t_L g130 ( 
.A1(n_85),
.A2(n_111),
.A3(n_89),
.B1(n_114),
.B2(n_102),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_130),
.A2(n_6),
.B(n_7),
.C(n_128),
.Y(n_195)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_81),
.B(n_28),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_135),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_55),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_91),
.A2(n_26),
.B1(n_19),
.B2(n_55),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_137),
.A2(n_152),
.B1(n_157),
.B2(n_99),
.Y(n_191)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_89),
.A2(n_86),
.B1(n_106),
.B2(n_94),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_144),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_147),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_16),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_86),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_106),
.A2(n_14),
.B1(n_12),
.B2(n_11),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_0),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_153),
.B(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_105),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_96),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_97),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_1),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_100),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_103),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_162),
.B(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_113),
.B(n_5),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_6),
.Y(n_192)
);

CKINVDCx11_ASAP7_75t_R g167 ( 
.A(n_126),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_167),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_80),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_186),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_190),
.B1(n_191),
.B2(n_194),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_136),
.B(n_153),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_195),
.B(n_175),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_124),
.B(n_110),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_142),
.B(n_80),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_197),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_154),
.A2(n_99),
.B1(n_117),
.B2(n_83),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_132),
.A2(n_117),
.B1(n_83),
.B2(n_7),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_155),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_141),
.B(n_7),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_141),
.A2(n_158),
.B1(n_146),
.B2(n_137),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_203),
.B1(n_194),
.B2(n_172),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_134),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_166),
.B1(n_165),
.B2(n_134),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_135),
.C(n_147),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_210),
.C(n_173),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_153),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_167),
.A2(n_138),
.B1(n_133),
.B2(n_163),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_158),
.B1(n_164),
.B2(n_160),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_221),
.B1(n_232),
.B2(n_182),
.Y(n_243)
);

OAI32xp33_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_161),
.A3(n_156),
.B1(n_131),
.B2(n_125),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_215),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_216),
.A2(n_233),
.B(n_189),
.Y(n_261)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_176),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_184),
.A2(n_204),
.B1(n_193),
.B2(n_202),
.Y(n_221)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_230),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_227),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_180),
.B(n_185),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_229),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_190),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_193),
.A2(n_198),
.B1(n_197),
.B2(n_183),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_168),
.A2(n_196),
.B(n_195),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_168),
.A2(n_196),
.B(n_191),
.C(n_177),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_189),
.Y(n_259)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_236),
.Y(n_256)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_174),
.B(n_192),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_169),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

INVx13_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_178),
.B(n_177),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_205),
.A2(n_169),
.B1(n_173),
.B2(n_188),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_241),
.A2(n_266),
.B1(n_227),
.B2(n_235),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_243),
.A2(n_245),
.B1(n_244),
.B2(n_259),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_251),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_225),
.B(n_232),
.CI(n_216),
.CON(n_252),
.SN(n_252)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_253),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_226),
.Y(n_253)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_254),
.Y(n_285)
);

OAI32xp33_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_207),
.A3(n_213),
.B1(n_221),
.B2(n_212),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_265),
.Y(n_275)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_233),
.A2(n_234),
.B(n_222),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_205),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_210),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_209),
.C(n_214),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_219),
.B1(n_231),
.B2(n_222),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_268),
.Y(n_294)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_270),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_234),
.B1(n_206),
.B2(n_215),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_280),
.B(n_284),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_239),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_286),
.C(n_251),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_256),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_277),
.Y(n_298)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_279),
.B(n_249),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_266),
.A2(n_237),
.B1(n_218),
.B2(n_217),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_284),
.Y(n_295)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_283),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_236),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_288),
.B1(n_246),
.B2(n_248),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_244),
.A2(n_246),
.B1(n_243),
.B2(n_245),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_255),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_293),
.A2(n_310),
.B1(n_272),
.B2(n_269),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_275),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_252),
.C(n_248),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_303),
.C(n_247),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_287),
.B(n_289),
.Y(n_301)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_265),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_302),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_252),
.C(n_261),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_309),
.B(n_302),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_273),
.B(n_252),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_311),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_285),
.B(n_263),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_290),
.A2(n_241),
.B1(n_249),
.B2(n_258),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_275),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_297),
.C(n_292),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_280),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_318),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_314),
.A2(n_295),
.B1(n_305),
.B2(n_297),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_240),
.CI(n_271),
.CON(n_315),
.SN(n_315)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_271),
.B1(n_281),
.B2(n_291),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_317),
.A2(n_324),
.B1(n_325),
.B2(n_298),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_240),
.Y(n_318)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_319),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_320),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_247),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_325),
.Y(n_338)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_293),
.CI(n_310),
.CON(n_322),
.SN(n_322)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_306),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_294),
.A2(n_258),
.B1(n_285),
.B2(n_263),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_326),
.B(n_309),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_308),
.A2(n_282),
.B(n_264),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_328),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_339),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_334),
.A2(n_336),
.B1(n_340),
.B2(n_315),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_320),
.A2(n_298),
.B1(n_304),
.B2(n_295),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_323),
.A2(n_316),
.B1(n_322),
.B2(n_313),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_318),
.C(n_327),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_326),
.B(n_316),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_343),
.A2(n_348),
.B(n_336),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_317),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_344),
.B(n_347),
.Y(n_359)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_321),
.C(n_322),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_346),
.Y(n_357)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_312),
.C(n_327),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_332),
.A2(n_315),
.B(n_282),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_349),
.B(n_338),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_340),
.C(n_330),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_352),
.C(n_247),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_292),
.C(n_264),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_351),
.A2(n_331),
.B(n_338),
.Y(n_353)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_353),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_342),
.B(n_299),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_356),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_355),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_344),
.A2(n_262),
.B1(n_254),
.B2(n_242),
.Y(n_358)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_352),
.A2(n_262),
.B(n_254),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_345),
.Y(n_362)
);

NAND2x1_ASAP7_75t_L g363 ( 
.A(n_361),
.B(n_346),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_362),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_357),
.Y(n_368)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_368),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_357),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_369),
.B(n_371),
.C(n_364),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_359),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_370),
.B(n_367),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_374),
.A2(n_372),
.B1(n_358),
.B2(n_363),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_375),
.B(n_242),
.C(n_371),
.Y(n_376)
);

BUFx24_ASAP7_75t_SL g377 ( 
.A(n_376),
.Y(n_377)
);


endmodule