module fake_jpeg_4466_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_42),
.Y(n_60)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_43),
.B1(n_48),
.B2(n_29),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_0),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_18),
.C(n_19),
.Y(n_74)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_20),
.B1(n_29),
.B2(n_27),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_48),
.B1(n_17),
.B2(n_28),
.Y(n_90)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_53),
.Y(n_100)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_67),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_27),
.B(n_17),
.C(n_24),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_64),
.B(n_48),
.Y(n_94)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_68),
.B(n_32),
.Y(n_98)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_74),
.B(n_42),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_78),
.B1(n_83),
.B2(n_31),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_20),
.B1(n_42),
.B2(n_29),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_41),
.B1(n_48),
.B2(n_17),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_48),
.B1(n_18),
.B2(n_19),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_39),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_93),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_61),
.B1(n_21),
.B2(n_28),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_39),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_72),
.B(n_61),
.C(n_49),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_19),
.B1(n_34),
.B2(n_31),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_44),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_98),
.Y(n_128)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_63),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_44),
.C(n_39),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_51),
.C(n_33),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_104),
.B1(n_117),
.B2(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_62),
.Y(n_103)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_57),
.B1(n_55),
.B2(n_21),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_122),
.B1(n_129),
.B2(n_130),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_44),
.C(n_39),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_127),
.C(n_77),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_107),
.A2(n_108),
.B1(n_32),
.B2(n_33),
.Y(n_156)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_124),
.Y(n_143)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_30),
.B1(n_28),
.B2(n_33),
.Y(n_117)
);

NAND2xp67_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_25),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_30),
.B(n_76),
.C(n_25),
.Y(n_144)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_44),
.B1(n_39),
.B2(n_37),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_83),
.B1(n_92),
.B2(n_81),
.Y(n_131)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_100),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_91),
.Y(n_136)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_104),
.B1(n_119),
.B2(n_115),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_157),
.B1(n_129),
.B2(n_23),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_96),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_90),
.B1(n_82),
.B2(n_81),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_148),
.B1(n_123),
.B2(n_116),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_99),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_107),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_144),
.A2(n_153),
.B(n_152),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_87),
.B1(n_92),
.B2(n_91),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_158),
.C(n_37),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_87),
.B(n_77),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_154),
.B(n_126),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_44),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_51),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_44),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_119),
.A2(n_121),
.B(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_11),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_79),
.B1(n_23),
.B2(n_26),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_79),
.C(n_39),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_160),
.A2(n_166),
.B1(n_167),
.B2(n_181),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_163),
.C(n_165),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_164),
.B(n_174),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_51),
.C(n_37),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_142),
.B1(n_149),
.B2(n_141),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_113),
.B1(n_105),
.B2(n_122),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_168),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_SL g211 ( 
.A1(n_169),
.A2(n_150),
.B(n_147),
.C(n_155),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_171),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_37),
.C(n_109),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_178),
.C(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_23),
.B1(n_26),
.B2(n_22),
.Y(n_175)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_138),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_22),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_26),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_130),
.B1(n_26),
.B2(n_22),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_184),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_26),
.B1(n_22),
.B2(n_125),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_183),
.Y(n_188)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_26),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_133),
.B(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_22),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_146),
.C(n_155),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_176),
.Y(n_226)
);

AOI22x1_ASAP7_75t_SL g195 ( 
.A1(n_162),
.A2(n_138),
.B1(n_137),
.B2(n_133),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g238 ( 
.A1(n_195),
.A2(n_16),
.B(n_15),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_199),
.B(n_200),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_177),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_145),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_212),
.C(n_214),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_145),
.B1(n_139),
.B2(n_147),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_25),
.B1(n_2),
.B2(n_4),
.Y(n_237)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_207),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_211),
.A2(n_184),
.B1(n_160),
.B2(n_161),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_146),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_150),
.Y(n_214)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_178),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_226),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_220),
.B1(n_242),
.B2(n_203),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_210),
.A2(n_163),
.B1(n_165),
.B2(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_223),
.B(n_235),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_206),
.A2(n_180),
.B(n_185),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_227),
.A2(n_240),
.B1(n_232),
.B2(n_202),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_187),
.C(n_171),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_234),
.C(n_218),
.Y(n_246)
);

XNOR2x2_ASAP7_75t_SL g232 ( 
.A(n_206),
.B(n_25),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_198),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_208),
.A2(n_159),
.B(n_25),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_237),
.B1(n_202),
.B2(n_204),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_201),
.C(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_194),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_211),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_241),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_248),
.C(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_191),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_250),
.Y(n_266)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_251),
.B(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_254),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_217),
.A2(n_197),
.B1(n_196),
.B2(n_192),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_263),
.B1(n_216),
.B2(n_225),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_205),
.B1(n_212),
.B2(n_188),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_256),
.A2(n_259),
.B1(n_228),
.B2(n_238),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_10),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_209),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_221),
.B(n_228),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_198),
.B1(n_209),
.B2(n_190),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_189),
.C(n_2),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_225),
.A2(n_189),
.B1(n_5),
.B2(n_6),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_0),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_220),
.B1(n_230),
.B2(n_227),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_283),
.B1(n_282),
.B2(n_270),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_233),
.B1(n_259),
.B2(n_265),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_272),
.B(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_280),
.Y(n_292)
);

AOI211xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_264),
.B(n_257),
.C(n_255),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_281),
.B(n_261),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_284),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_5),
.C(n_6),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_262),
.C(n_252),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_10),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_256),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_286),
.B(n_284),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_299),
.B1(n_279),
.B2(n_12),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_291),
.A2(n_294),
.B(n_297),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_252),
.Y(n_294)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_274),
.A2(n_245),
.B(n_7),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_8),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_276),
.A2(n_245),
.B1(n_7),
.B2(n_8),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_6),
.C(n_7),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_269),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_285),
.C(n_300),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_278),
.Y(n_304)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_304),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_306),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_295),
.B(n_273),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_311),
.Y(n_321)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_292),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_310),
.B(n_313),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_13),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_288),
.B(n_13),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_13),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_8),
.Y(n_315)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_294),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_314),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_285),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_320),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_289),
.Y(n_320)
);

FAx1_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_296),
.CI(n_307),
.CON(n_331),
.SN(n_331)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_289),
.C(n_298),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_291),
.Y(n_326)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_326),
.A2(n_330),
.B(n_317),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_312),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_331),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_319),
.B(n_308),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_321),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_332),
.B(n_315),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_336),
.C(n_14),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_335),
.B(n_327),
.Y(n_338)
);

A2O1A1Ixp33_ASAP7_75t_SL g336 ( 
.A1(n_328),
.A2(n_15),
.B(n_14),
.C(n_9),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_338),
.B(n_339),
.C(n_325),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_337),
.B(n_334),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_341),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_14),
.B(n_9),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_9),
.Y(n_344)
);


endmodule