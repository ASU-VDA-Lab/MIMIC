module fake_jpeg_20164_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_1),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_1),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_1),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_16),
.B1(n_33),
.B2(n_22),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_48),
.Y(n_84)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_33),
.B1(n_39),
.B2(n_37),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_79),
.B1(n_86),
.B2(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_44),
.B1(n_42),
.B2(n_40),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_85),
.B1(n_96),
.B2(n_65),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_69),
.B(n_81),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_33),
.B1(n_39),
.B2(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_42),
.B(n_30),
.C(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_43),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_40),
.B1(n_35),
.B2(n_37),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_39),
.B1(n_35),
.B2(n_20),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_40),
.B1(n_35),
.B2(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_24),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_21),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_64),
.B1(n_65),
.B2(n_29),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_21),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_78),
.B1(n_93),
.B2(n_81),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_63),
.B1(n_65),
.B2(n_29),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_120),
.Y(n_153)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_28),
.B1(n_23),
.B2(n_19),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_32),
.B1(n_63),
.B2(n_70),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_28),
.B1(n_23),
.B2(n_19),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_70),
.B1(n_90),
.B2(n_82),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_119),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_21),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_73),
.A2(n_26),
.B1(n_32),
.B2(n_34),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_85),
.B1(n_90),
.B2(n_74),
.Y(n_140)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_94),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_24),
.Y(n_124)
);

XNOR2x1_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_68),
.Y(n_127)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_36),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_83),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_148),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_130),
.A2(n_145),
.B1(n_155),
.B2(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_69),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_132),
.B(n_136),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_80),
.B(n_76),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_133),
.A2(n_147),
.B(n_113),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_154),
.B(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_99),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_100),
.B1(n_123),
.B2(n_106),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_143),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_75),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_43),
.B1(n_36),
.B2(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_2),
.B(n_3),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_114),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_99),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_152),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_100),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_94),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_125),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_156),
.B(n_160),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_169),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_98),
.B(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_165),
.Y(n_198)
);

HAxp5_ASAP7_75t_SL g191 ( 
.A(n_164),
.B(n_186),
.CON(n_191),
.SN(n_191)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_125),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_174),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_21),
.C(n_24),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_133),
.A2(n_21),
.B(n_24),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_187),
.B(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_155),
.A2(n_110),
.B1(n_116),
.B2(n_97),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_175),
.A2(n_177),
.B1(n_145),
.B2(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_134),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_178),
.B(n_183),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_134),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_180),
.Y(n_192)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_116),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_137),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_126),
.B(n_97),
.C(n_113),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_130),
.C(n_148),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_126),
.A2(n_2),
.B(n_3),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_25),
.Y(n_190)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_200),
.B1(n_214),
.B2(n_177),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_199),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_144),
.B1(n_149),
.B2(n_152),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_179),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_201),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_185),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_131),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_197),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_136),
.C(n_135),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_207),
.C(n_216),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_141),
.C(n_34),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_209),
.A2(n_190),
.B(n_161),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_157),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_158),
.A2(n_34),
.B1(n_31),
.B2(n_25),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_34),
.C(n_25),
.Y(n_216)
);

AO32x1_ASAP7_75t_L g219 ( 
.A1(n_178),
.A2(n_10),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_219),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_198),
.B(n_186),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_222),
.B1(n_209),
.B2(n_192),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_164),
.B(n_183),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_171),
.B1(n_188),
.B2(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_188),
.B1(n_159),
.B2(n_162),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_174),
.B(n_165),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_234),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_187),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_233),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_169),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_193),
.A2(n_211),
.B1(n_218),
.B2(n_199),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_239),
.B1(n_244),
.B2(n_214),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_161),
.B(n_170),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_240),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_173),
.C(n_189),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_217),
.C(n_203),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_193),
.A2(n_176),
.B1(n_157),
.B2(n_17),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_212),
.B(n_195),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_207),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_216),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_218),
.A2(n_17),
.B1(n_31),
.B2(n_5),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_203),
.Y(n_248)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_235),
.C(n_202),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_255),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_225),
.A2(n_215),
.B1(n_205),
.B2(n_208),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_244),
.B1(n_221),
.B2(n_226),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_228),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_262),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_215),
.C(n_205),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_230),
.C(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_208),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_219),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_236),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_238),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_266),
.A2(n_255),
.B1(n_11),
.B2(n_12),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_220),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_230),
.C(n_232),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_274),
.C(n_275),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_264),
.A2(n_241),
.B(n_237),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_276),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_273),
.A2(n_245),
.B1(n_246),
.B2(n_249),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_222),
.C(n_233),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_228),
.C(n_241),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_248),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_9),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_9),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g281 ( 
.A(n_266),
.B(n_254),
.CI(n_256),
.CON(n_281),
.SN(n_281)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_284),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_261),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_263),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_289),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_270),
.A2(n_250),
.B1(n_246),
.B2(n_258),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_247),
.B1(n_257),
.B2(n_259),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_247),
.B1(n_272),
.B2(n_274),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_8),
.B(n_13),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_8),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_265),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_11),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_8),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_268),
.C(n_269),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_300),
.C(n_291),
.Y(n_310)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_283),
.B(n_281),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_267),
.C(n_31),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_290),
.B(n_288),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_295),
.B(n_7),
.C(n_12),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_285),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_15),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_312),
.B(n_313),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_15),
.B1(n_7),
.B2(n_11),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_308),
.A2(n_297),
.B(n_301),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_310),
.B(n_309),
.Y(n_320)
);

NOR2x1_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_307),
.Y(n_319)
);

OAI311xp33_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_320),
.A3(n_314),
.B1(n_315),
.C1(n_12),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_321),
.C(n_4),
.Y(n_323)
);

OAI31xp33_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_3),
.A3(n_6),
.B(n_322),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_3),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_6),
.B(n_195),
.Y(n_326)
);


endmodule