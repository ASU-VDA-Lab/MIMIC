module fake_jpeg_29666_n_112 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_112);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_8),
.B(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_23),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_20),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_26),
.A2(n_33),
.B1(n_12),
.B2(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_20),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.Y(n_38)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_44),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_15),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_21),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_33),
.B1(n_12),
.B2(n_19),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_17),
.B1(n_22),
.B2(n_19),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_27),
.B1(n_22),
.B2(n_36),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_31),
.B1(n_28),
.B2(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_69),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_37),
.A2(n_22),
.B1(n_29),
.B2(n_36),
.Y(n_61)
);

BUFx12f_ASAP7_75t_SL g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_34),
.B1(n_29),
.B2(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_67),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_34),
.B(n_23),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_68),
.B(n_23),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_14),
.B1(n_24),
.B2(n_18),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_24),
.B1(n_18),
.B2(n_16),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_43),
.B(n_39),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_66),
.C(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_7),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_54),
.Y(n_96)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_57),
.Y(n_86)
);

AOI322xp5_ASAP7_75t_SL g94 ( 
.A1(n_86),
.A2(n_46),
.A3(n_67),
.B1(n_74),
.B2(n_40),
.C1(n_9),
.C2(n_8),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_59),
.B1(n_65),
.B2(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_89),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_70),
.C(n_79),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_92),
.Y(n_98)
);

A2O1A1O1Ixp25_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_78),
.B(n_74),
.C(n_72),
.D(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_89),
.B(n_83),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_9),
.B1(n_86),
.B2(n_4),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_96),
.A2(n_81),
.B1(n_95),
.B2(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_101),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_90),
.A2(n_87),
.B1(n_51),
.B2(n_46),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_90),
.C(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_95),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_106),
.A2(n_100),
.B(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_101),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_108),
.B1(n_103),
.B2(n_102),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_110),
.B(n_4),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_23),
.Y(n_112)
);


endmodule