module real_aes_17836_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1835;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1784;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_1779;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1800;
wire n_1435;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1802;
wire n_727;
wire n_397;
wire n_1056;
wire n_1083;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1790;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_1826;
wire n_1836;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1823;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1280;
wire n_729;
wire n_394;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_0), .A2(n_284), .B1(n_720), .B2(n_721), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_0), .A2(n_177), .B1(n_619), .B2(n_768), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_1), .A2(n_61), .B1(n_587), .B2(n_590), .Y(n_1115) );
INVxp67_ASAP7_75t_SL g1135 ( .A(n_1), .Y(n_1135) );
INVx1_ASAP7_75t_L g1291 ( .A(n_2), .Y(n_1291) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_3), .A2(n_276), .B1(n_507), .B2(n_512), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_3), .A2(n_355), .B1(n_549), .B2(n_551), .Y(n_548) );
INVx1_ASAP7_75t_L g389 ( .A(n_4), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_4), .B(n_399), .Y(n_505) );
INVx1_ASAP7_75t_L g745 ( .A(n_5), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_5), .A2(n_201), .B1(n_568), .B2(n_756), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g1160 ( .A(n_6), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1253 ( .A1(n_7), .A2(n_271), .B1(n_512), .B2(n_1254), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_7), .A2(n_208), .B1(n_1271), .B2(n_1272), .Y(n_1270) );
INVx1_ASAP7_75t_L g1815 ( .A(n_8), .Y(n_1815) );
INVx1_ASAP7_75t_L g1752 ( .A(n_9), .Y(n_1752) );
OAI22xp33_ASAP7_75t_SL g1173 ( .A1(n_10), .A2(n_361), .B1(n_580), .B2(n_1120), .Y(n_1173) );
OAI22xp33_ASAP7_75t_L g1184 ( .A1(n_10), .A2(n_192), .B1(n_485), .B2(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g947 ( .A(n_11), .Y(n_947) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_12), .A2(n_56), .B1(n_1526), .B2(n_1534), .Y(n_1580) );
INVx1_ASAP7_75t_L g1246 ( .A(n_13), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_13), .A2(n_271), .B1(n_1272), .B2(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g751 ( .A(n_14), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g1067 ( .A(n_15), .Y(n_1067) );
INVx1_ASAP7_75t_L g1097 ( .A(n_16), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1478 ( .A1(n_17), .A2(n_46), .B1(n_841), .B2(n_1479), .Y(n_1478) );
OAI22xp33_ASAP7_75t_L g1494 ( .A1(n_17), .A2(n_46), .B1(n_391), .B2(n_662), .Y(n_1494) );
INVx1_ASAP7_75t_L g1775 ( .A(n_18), .Y(n_1775) );
OAI211xp5_ASAP7_75t_L g1783 ( .A1(n_18), .A2(n_642), .B(n_1784), .C(n_1785), .Y(n_1783) );
INVx1_ASAP7_75t_L g1331 ( .A(n_19), .Y(n_1331) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_19), .A2(n_319), .B1(n_569), .B2(n_641), .C(n_1339), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_20), .A2(n_124), .B1(n_720), .B2(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g766 ( .A(n_20), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g1192 ( .A(n_21), .Y(n_1192) );
XOR2x2_ASAP7_75t_L g558 ( .A(n_22), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g1756 ( .A(n_23), .Y(n_1756) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_24), .A2(n_338), .B1(n_833), .B2(n_834), .Y(n_1039) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_24), .A2(n_338), .B1(n_636), .B2(n_847), .Y(n_1042) );
INVx2_ASAP7_75t_L g457 ( .A(n_25), .Y(n_457) );
XNOR2xp5_ASAP7_75t_L g1086 ( .A(n_26), .B(n_1087), .Y(n_1086) );
OAI22xp33_ASAP7_75t_SL g1386 ( .A1(n_27), .A2(n_282), .B1(n_485), .B2(n_1185), .Y(n_1386) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_27), .A2(n_282), .B1(n_580), .B2(n_921), .Y(n_1393) );
INVx1_ASAP7_75t_L g940 ( .A(n_28), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g1346 ( .A1(n_29), .A2(n_298), .B1(n_1347), .B2(n_1349), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_29), .A2(n_165), .B1(n_617), .B2(n_1356), .Y(n_1355) );
INVx1_ASAP7_75t_L g874 ( .A(n_30), .Y(n_874) );
INVx1_ASAP7_75t_L g987 ( .A(n_31), .Y(n_987) );
INVx1_ASAP7_75t_L g1401 ( .A(n_32), .Y(n_1401) );
AOI22xp5_ASAP7_75t_L g1562 ( .A1(n_32), .A2(n_232), .B1(n_1538), .B2(n_1541), .Y(n_1562) );
INVx1_ASAP7_75t_L g1763 ( .A(n_33), .Y(n_1763) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_34), .A2(n_340), .B1(n_440), .B2(n_441), .Y(n_919) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_34), .A2(n_340), .B1(n_454), .B2(n_462), .Y(n_930) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_35), .A2(n_94), .B1(n_454), .B2(n_1185), .C(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1315 ( .A(n_35), .Y(n_1315) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_36), .Y(n_384) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_36), .B(n_382), .Y(n_1527) );
AOI22xp5_ASAP7_75t_L g1579 ( .A1(n_37), .A2(n_206), .B1(n_1538), .B2(n_1541), .Y(n_1579) );
OAI22xp33_ASAP7_75t_SL g1804 ( .A1(n_38), .A2(n_178), .B1(n_833), .B2(n_834), .Y(n_1804) );
OAI22xp5_ASAP7_75t_L g1806 ( .A1(n_38), .A2(n_178), .B1(n_847), .B2(n_848), .Y(n_1806) );
AOI22xp5_ASAP7_75t_L g1554 ( .A1(n_39), .A2(n_297), .B1(n_1538), .B2(n_1541), .Y(n_1554) );
CKINVDCx5p33_ASAP7_75t_R g1450 ( .A(n_40), .Y(n_1450) );
AOI22xp33_ASAP7_75t_SL g613 ( .A1(n_41), .A2(n_280), .B1(n_512), .B2(n_604), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_41), .A2(n_164), .B1(n_616), .B2(n_617), .Y(n_621) );
INVx1_ASAP7_75t_L g804 ( .A(n_42), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g1572 ( .A1(n_43), .A2(n_125), .B1(n_1538), .B2(n_1541), .Y(n_1572) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_44), .A2(n_197), .B1(n_885), .B2(n_886), .Y(n_884) );
OAI22xp33_ASAP7_75t_L g898 ( .A1(n_44), .A2(n_197), .B1(n_391), .B2(n_899), .Y(n_898) );
INVxp67_ASAP7_75t_SL g1114 ( .A(n_45), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_45), .A2(n_61), .B1(n_472), .B2(n_1137), .Y(n_1136) );
AOI22xp5_ASAP7_75t_L g1570 ( .A1(n_47), .A2(n_179), .B1(n_1534), .B2(n_1571), .Y(n_1570) );
OAI22xp33_ASAP7_75t_L g920 ( .A1(n_48), .A2(n_289), .B1(n_580), .B2(n_921), .Y(n_920) );
OAI22xp33_ASAP7_75t_SL g923 ( .A1(n_48), .A2(n_289), .B1(n_485), .B2(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g1012 ( .A(n_49), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_49), .A2(n_366), .B1(n_907), .B2(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1498 ( .A(n_50), .Y(n_1498) );
INVx1_ASAP7_75t_L g895 ( .A(n_51), .Y(n_895) );
OAI211xp5_ASAP7_75t_L g900 ( .A1(n_51), .A2(n_828), .B(n_901), .C(n_904), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_52), .A2(n_309), .B1(n_440), .B2(n_441), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_52), .A2(n_309), .B1(n_454), .B2(n_462), .Y(n_453) );
XNOR2x1_ASAP7_75t_L g1363 ( .A(n_53), .B(n_1364), .Y(n_1363) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_54), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g1244 ( .A(n_55), .Y(n_1244) );
INVx1_ASAP7_75t_L g695 ( .A(n_57), .Y(n_695) );
INVx1_ASAP7_75t_L g1294 ( .A(n_58), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_59), .A2(n_279), .B1(n_515), .B2(n_518), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_59), .A2(n_100), .B1(n_545), .B2(n_547), .Y(n_544) );
INVx1_ASAP7_75t_L g979 ( .A(n_60), .Y(n_979) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_62), .B(n_475), .Y(n_1304) );
INVxp67_ASAP7_75t_SL g1312 ( .A(n_62), .Y(n_1312) );
OAI211xp5_ASAP7_75t_SL g1480 ( .A1(n_63), .A2(n_808), .B(n_889), .C(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1491 ( .A(n_63), .Y(n_1491) );
AOI22xp33_ASAP7_75t_L g1533 ( .A1(n_64), .A2(n_252), .B1(n_1526), .B2(n_1534), .Y(n_1533) );
OAI211xp5_ASAP7_75t_L g1168 ( .A1(n_65), .A2(n_914), .B(n_1169), .C(n_1170), .Y(n_1168) );
INVx1_ASAP7_75t_L g1183 ( .A(n_65), .Y(n_1183) );
INVx1_ASAP7_75t_L g872 ( .A(n_66), .Y(n_872) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_67), .A2(n_250), .B1(n_454), .B2(n_636), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_67), .A2(n_250), .B1(n_659), .B2(n_660), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g1484 ( .A1(n_68), .A2(n_187), .B1(n_636), .B2(n_847), .Y(n_1484) );
OAI22xp5_ASAP7_75t_L g1492 ( .A1(n_68), .A2(n_187), .B1(n_833), .B2(n_1493), .Y(n_1492) );
CKINVDCx5p33_ASAP7_75t_R g1152 ( .A(n_69), .Y(n_1152) );
INVx1_ASAP7_75t_L g1117 ( .A(n_70), .Y(n_1117) );
INVx1_ASAP7_75t_L g692 ( .A(n_71), .Y(n_692) );
OAI222xp33_ASAP7_75t_L g1233 ( .A1(n_72), .A2(n_195), .B1(n_434), .B2(n_581), .C1(n_1234), .C2(n_1235), .Y(n_1233) );
OAI222xp33_ASAP7_75t_L g1260 ( .A1(n_72), .A2(n_195), .B1(n_237), .B2(n_568), .C1(n_1261), .C2(n_1262), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1334 ( .A1(n_73), .A2(n_130), .B1(n_440), .B2(n_441), .Y(n_1334) );
OAI22xp5_ASAP7_75t_L g1340 ( .A1(n_73), .A2(n_130), .B1(n_454), .B2(n_462), .Y(n_1340) );
INVx1_ASAP7_75t_L g946 ( .A(n_74), .Y(n_946) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_75), .A2(n_324), .B1(n_391), .B2(n_662), .Y(n_835) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_75), .A2(n_324), .B1(n_839), .B2(n_841), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g1307 ( .A1(n_76), .A2(n_198), .B1(n_485), .B2(n_1308), .Y(n_1307) );
INVxp67_ASAP7_75t_SL g1314 ( .A(n_76), .Y(n_1314) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_77), .Y(n_1203) );
OAI22xp33_ASAP7_75t_L g896 ( .A1(n_78), .A2(n_184), .B1(n_847), .B2(n_848), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_78), .A2(n_184), .B1(n_834), .B2(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g1118 ( .A(n_79), .Y(n_1118) );
INVx1_ASAP7_75t_L g1508 ( .A(n_80), .Y(n_1508) );
CKINVDCx5p33_ASAP7_75t_R g1414 ( .A(n_81), .Y(n_1414) );
INVx1_ASAP7_75t_L g1378 ( .A(n_82), .Y(n_1378) );
OAI211xp5_ASAP7_75t_L g912 ( .A1(n_83), .A2(n_913), .B(n_914), .C(n_915), .Y(n_912) );
INVx1_ASAP7_75t_L g927 ( .A(n_83), .Y(n_927) );
INVx1_ASAP7_75t_L g1110 ( .A(n_84), .Y(n_1110) );
INVx1_ASAP7_75t_L g717 ( .A(n_85), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g418 ( .A1(n_86), .A2(n_419), .B(n_423), .C(n_429), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g466 ( .A1(n_86), .A2(n_215), .B1(n_467), .B2(n_472), .C(n_477), .Y(n_466) );
XOR2xp5_ASAP7_75t_L g1795 ( .A(n_87), .B(n_1796), .Y(n_1795) );
XNOR2xp5_ASAP7_75t_L g1320 ( .A(n_88), .B(n_1321), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1550 ( .A1(n_88), .A2(n_182), .B1(n_1534), .B2(n_1538), .Y(n_1550) );
INVx1_ASAP7_75t_L g1293 ( .A(n_89), .Y(n_1293) );
INVx1_ASAP7_75t_L g1826 ( .A(n_90), .Y(n_1826) );
OAI22xp33_ASAP7_75t_L g1391 ( .A1(n_91), .A2(n_122), .B1(n_454), .B2(n_462), .Y(n_1391) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_91), .A2(n_122), .B1(n_440), .B2(n_441), .Y(n_1397) );
XNOR2xp5_ASAP7_75t_L g1439 ( .A(n_92), .B(n_1440), .Y(n_1439) );
AOI22xp33_ASAP7_75t_L g1549 ( .A1(n_93), .A2(n_321), .B1(n_1526), .B2(n_1541), .Y(n_1549) );
OAI22xp33_ASAP7_75t_L g1317 ( .A1(n_94), .A2(n_198), .B1(n_580), .B2(n_921), .Y(n_1317) );
AOI22xp5_ASAP7_75t_L g1556 ( .A1(n_95), .A2(n_163), .B1(n_1534), .B2(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1428 ( .A(n_96), .Y(n_1428) );
OAI211xp5_ASAP7_75t_L g1433 ( .A1(n_96), .A2(n_642), .B(n_1434), .C(n_1436), .Y(n_1433) );
OAI22xp5_ASAP7_75t_L g1214 ( .A1(n_97), .A2(n_287), .B1(n_441), .B2(n_580), .Y(n_1214) );
OAI22xp5_ASAP7_75t_SL g1222 ( .A1(n_97), .A2(n_138), .B1(n_462), .B2(n_485), .Y(n_1222) );
INVx1_ASAP7_75t_L g1306 ( .A(n_98), .Y(n_1306) );
INVx1_ASAP7_75t_L g1507 ( .A(n_99), .Y(n_1507) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_100), .A2(n_365), .B1(n_512), .B2(n_525), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g1217 ( .A(n_101), .Y(n_1217) );
INVx1_ASAP7_75t_L g950 ( .A(n_102), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g1191 ( .A(n_103), .Y(n_1191) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_104), .Y(n_1151) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_105), .A2(n_639), .B(n_642), .C(n_643), .Y(n_638) );
INVx1_ASAP7_75t_L g656 ( .A(n_105), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g1350 ( .A1(n_106), .A2(n_263), .B1(n_1347), .B2(n_1351), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_106), .A2(n_174), .B1(n_549), .B2(n_1358), .Y(n_1357) );
XOR2xp5_ASAP7_75t_L g1146 ( .A(n_107), .B(n_1147), .Y(n_1146) );
XNOR2x2_ASAP7_75t_SL g632 ( .A(n_108), .B(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_108), .A2(n_350), .B1(n_1538), .B2(n_1541), .Y(n_1537) );
INVx1_ASAP7_75t_L g1099 ( .A(n_109), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_109), .A2(n_307), .B1(n_507), .B2(n_1127), .Y(n_1132) );
CKINVDCx5p33_ASAP7_75t_R g1453 ( .A(n_110), .Y(n_1453) );
CKINVDCx5p33_ASAP7_75t_R g1200 ( .A(n_111), .Y(n_1200) );
OAI22xp33_ASAP7_75t_L g1771 ( .A1(n_112), .A2(n_119), .B1(n_580), .B2(n_662), .Y(n_1771) );
OAI22xp33_ASAP7_75t_L g1778 ( .A1(n_112), .A2(n_119), .B1(n_1779), .B2(n_1780), .Y(n_1778) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_113), .A2(n_238), .B1(n_568), .B2(n_569), .Y(n_567) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_113), .Y(n_585) );
INVx1_ASAP7_75t_L g917 ( .A(n_114), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_115), .A2(n_304), .B1(n_512), .B2(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_115), .A2(n_278), .B1(n_619), .B2(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g810 ( .A(n_116), .Y(n_810) );
OAI211xp5_ASAP7_75t_L g1425 ( .A1(n_117), .A2(n_818), .B(n_914), .C(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1437 ( .A(n_117), .Y(n_1437) );
INVx1_ASAP7_75t_L g382 ( .A(n_118), .Y(n_382) );
INVx1_ASAP7_75t_L g1106 ( .A(n_120), .Y(n_1106) );
INVxp67_ASAP7_75t_SL g565 ( .A(n_121), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_121), .A2(n_238), .B1(n_587), .B2(n_590), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g1430 ( .A1(n_123), .A2(n_315), .B1(n_659), .B2(n_662), .Y(n_1430) );
OAI22xp33_ASAP7_75t_L g1438 ( .A1(n_123), .A2(n_168), .B1(n_454), .B2(n_462), .Y(n_1438) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_124), .Y(n_773) );
XOR2xp5_ASAP7_75t_L g1227 ( .A(n_125), .B(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1371 ( .A(n_126), .Y(n_1371) );
INVx1_ASAP7_75t_L g1368 ( .A(n_127), .Y(n_1368) );
INVx1_ASAP7_75t_L g1802 ( .A(n_128), .Y(n_1802) );
INVx1_ASAP7_75t_L g746 ( .A(n_129), .Y(n_746) );
INVx1_ASAP7_75t_L g791 ( .A(n_131), .Y(n_791) );
INVx1_ASAP7_75t_L g1095 ( .A(n_132), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1776 ( .A1(n_133), .A2(n_311), .B1(n_907), .B2(n_1120), .Y(n_1776) );
OAI22xp5_ASAP7_75t_L g1781 ( .A1(n_133), .A2(n_311), .B1(n_848), .B2(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1774 ( .A(n_134), .Y(n_1774) );
INVx1_ASAP7_75t_L g1818 ( .A(n_135), .Y(n_1818) );
AOI22xp33_ASAP7_75t_SL g1553 ( .A1(n_136), .A2(n_224), .B1(n_1526), .B2(n_1534), .Y(n_1553) );
INVx1_ASAP7_75t_L g1746 ( .A(n_136), .Y(n_1746) );
AOI22xp33_ASAP7_75t_L g1790 ( .A1(n_136), .A2(n_1791), .B1(n_1794), .B2(n_1832), .Y(n_1790) );
OAI22xp33_ASAP7_75t_SL g1219 ( .A1(n_137), .A2(n_138), .B1(n_440), .B2(n_921), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1225 ( .A1(n_137), .A2(n_142), .B1(n_1181), .B2(n_1182), .Y(n_1225) );
INVx1_ASAP7_75t_L g1511 ( .A(n_139), .Y(n_1511) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_140), .Y(n_1062) );
INVx1_ASAP7_75t_L g868 ( .A(n_141), .Y(n_868) );
INVx1_ASAP7_75t_L g1218 ( .A(n_142), .Y(n_1218) );
OAI22xp33_ASAP7_75t_L g647 ( .A1(n_143), .A2(n_359), .B1(n_485), .B2(n_648), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_143), .A2(n_359), .B1(n_580), .B2(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g694 ( .A(n_144), .Y(n_694) );
INVx1_ASAP7_75t_L g1324 ( .A(n_145), .Y(n_1324) );
INVx1_ASAP7_75t_L g1390 ( .A(n_146), .Y(n_1390) );
OAI211xp5_ASAP7_75t_L g1394 ( .A1(n_146), .A2(n_730), .B(n_914), .C(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g718 ( .A(n_147), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_148), .Y(n_1389) );
CKINVDCx5p33_ASAP7_75t_R g1066 ( .A(n_149), .Y(n_1066) );
CKINVDCx5p33_ASAP7_75t_R g1451 ( .A(n_150), .Y(n_1451) );
OAI22xp33_ASAP7_75t_L g1466 ( .A1(n_151), .A2(n_199), .B1(n_440), .B2(n_662), .Y(n_1466) );
OAI22xp33_ASAP7_75t_L g1472 ( .A1(n_151), .A2(n_190), .B1(n_454), .B2(n_462), .Y(n_1472) );
CKINVDCx5p33_ASAP7_75t_R g1195 ( .A(n_152), .Y(n_1195) );
CKINVDCx5p33_ASAP7_75t_R g1444 ( .A(n_153), .Y(n_1444) );
OAI211xp5_ASAP7_75t_L g1800 ( .A1(n_154), .A2(n_828), .B(n_1488), .C(n_1801), .Y(n_1800) );
INVx1_ASAP7_75t_L g1810 ( .A(n_154), .Y(n_1810) );
INVx1_ASAP7_75t_L g1803 ( .A(n_155), .Y(n_1803) );
OAI211xp5_ASAP7_75t_L g1807 ( .A1(n_155), .A2(n_642), .B(n_1808), .C(n_1809), .Y(n_1807) );
INVx1_ASAP7_75t_L g1502 ( .A(n_156), .Y(n_1502) );
INVx1_ASAP7_75t_L g689 ( .A(n_157), .Y(n_689) );
INVx1_ASAP7_75t_L g1482 ( .A(n_158), .Y(n_1482) );
INVx1_ASAP7_75t_L g1816 ( .A(n_159), .Y(n_1816) );
CKINVDCx5p33_ASAP7_75t_R g1154 ( .A(n_160), .Y(n_1154) );
INVx1_ASAP7_75t_L g1760 ( .A(n_161), .Y(n_1760) );
OAI211xp5_ASAP7_75t_L g827 ( .A1(n_162), .A2(n_704), .B(n_828), .C(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g845 ( .A(n_162), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_164), .A2(n_346), .B1(n_599), .B2(n_602), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g1352 ( .A1(n_165), .A2(n_219), .B1(n_735), .B2(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g830 ( .A(n_166), .Y(n_830) );
OAI211xp5_ASAP7_75t_L g1772 ( .A1(n_167), .A2(n_914), .B(n_1169), .C(n_1773), .Y(n_1772) );
INVx1_ASAP7_75t_L g1786 ( .A(n_167), .Y(n_1786) );
OAI22xp33_ASAP7_75t_L g1429 ( .A1(n_168), .A2(n_291), .B1(n_580), .B2(n_741), .Y(n_1429) );
INVx1_ASAP7_75t_L g1464 ( .A(n_169), .Y(n_1464) );
OAI211xp5_ASAP7_75t_L g1469 ( .A1(n_169), .A2(n_642), .B(n_1434), .C(n_1470), .Y(n_1469) );
CKINVDCx5p33_ASAP7_75t_R g1406 ( .A(n_170), .Y(n_1406) );
INVx1_ASAP7_75t_L g1290 ( .A(n_171), .Y(n_1290) );
INVx1_ASAP7_75t_L g1326 ( .A(n_172), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_173), .A2(n_303), .B1(n_833), .B2(n_834), .Y(n_832) );
OAI22xp33_ASAP7_75t_L g846 ( .A1(n_173), .A2(n_303), .B1(n_847), .B2(n_848), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g1343 ( .A1(n_174), .A2(n_281), .B1(n_1344), .B2(n_1345), .Y(n_1343) );
OAI211xp5_ASAP7_75t_L g1461 ( .A1(n_175), .A2(n_818), .B(n_914), .C(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1471 ( .A(n_175), .Y(n_1471) );
INVxp67_ASAP7_75t_SL g729 ( .A(n_176), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g767 ( .A1(n_176), .A2(n_284), .B1(n_768), .B2(n_769), .Y(n_767) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_177), .Y(n_731) );
CKINVDCx5p33_ASAP7_75t_R g1157 ( .A(n_180), .Y(n_1157) );
XNOR2xp5_ASAP7_75t_L g711 ( .A(n_181), .B(n_712), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g1330 ( .A(n_183), .Y(n_1330) );
INVx1_ASAP7_75t_L g1825 ( .A(n_185), .Y(n_1825) );
INVx1_ASAP7_75t_L g807 ( .A(n_186), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g1465 ( .A1(n_188), .A2(n_190), .B1(n_580), .B2(n_741), .Y(n_1465) );
OAI22xp33_ASAP7_75t_L g1468 ( .A1(n_188), .A2(n_199), .B1(n_485), .B2(n_1185), .Y(n_1468) );
INVx1_ASAP7_75t_L g1483 ( .A(n_189), .Y(n_1483) );
OAI211xp5_ASAP7_75t_L g1487 ( .A1(n_189), .A2(n_828), .B(n_1488), .C(n_1490), .Y(n_1487) );
OAI211xp5_ASAP7_75t_L g1387 ( .A1(n_191), .A2(n_642), .B(n_1105), .C(n_1388), .Y(n_1387) );
INVx1_ASAP7_75t_L g1396 ( .A(n_191), .Y(n_1396) );
OAI22xp33_ASAP7_75t_SL g1174 ( .A1(n_192), .A2(n_328), .B1(n_659), .B2(n_662), .Y(n_1174) );
INVx1_ASAP7_75t_L g1751 ( .A(n_193), .Y(n_1751) );
INVx1_ASAP7_75t_L g787 ( .A(n_194), .Y(n_787) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_196), .B(n_320), .Y(n_1528) );
INVx2_ASAP7_75t_L g1536 ( .A(n_196), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_196), .B(n_1540), .Y(n_1542) );
CKINVDCx5p33_ASAP7_75t_R g1448 ( .A(n_200), .Y(n_1448) );
INVx1_ASAP7_75t_L g748 ( .A(n_201), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g1198 ( .A(n_202), .Y(n_1198) );
INVx1_ASAP7_75t_L g1499 ( .A(n_203), .Y(n_1499) );
INVx1_ASAP7_75t_L g863 ( .A(n_204), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g1564 ( .A1(n_205), .A2(n_262), .B1(n_1534), .B2(n_1541), .Y(n_1564) );
INVx1_ASAP7_75t_L g411 ( .A(n_207), .Y(n_411) );
INVx1_ASAP7_75t_L g1247 ( .A(n_208), .Y(n_1247) );
XOR2xp5_ASAP7_75t_L g1279 ( .A(n_209), .B(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g1014 ( .A(n_210), .Y(n_1014) );
OAI22xp33_ASAP7_75t_L g1028 ( .A1(n_210), .A2(n_247), .B1(n_580), .B2(n_662), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_211), .A2(n_216), .B1(n_1538), .B2(n_1557), .Y(n_1565) );
INVx1_ASAP7_75t_L g1285 ( .A(n_212), .Y(n_1285) );
CKINVDCx5p33_ASAP7_75t_R g1412 ( .A(n_213), .Y(n_1412) );
INVx1_ASAP7_75t_L g916 ( .A(n_214), .Y(n_916) );
INVx1_ASAP7_75t_L g438 ( .A(n_215), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_217), .A2(n_278), .B1(n_602), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_217), .A2(n_304), .B1(n_549), .B2(n_619), .Y(n_618) );
XOR2x2_ASAP7_75t_L g909 ( .A(n_218), .B(n_910), .Y(n_909) );
AOI22xp33_ASAP7_75t_SL g1360 ( .A1(n_219), .A2(n_298), .B1(n_617), .B2(n_680), .Y(n_1360) );
INVx1_ASAP7_75t_L g860 ( .A(n_220), .Y(n_860) );
CKINVDCx5p33_ASAP7_75t_R g1037 ( .A(n_221), .Y(n_1037) );
OAI211xp5_ASAP7_75t_L g1230 ( .A1(n_222), .A2(n_899), .B(n_1231), .C(n_1239), .Y(n_1230) );
INVx1_ASAP7_75t_L g1265 ( .A(n_222), .Y(n_1265) );
INVx1_ASAP7_75t_L g794 ( .A(n_223), .Y(n_794) );
INVx1_ASAP7_75t_L g1288 ( .A(n_225), .Y(n_1288) );
OAI22xp33_ASAP7_75t_L g1799 ( .A1(n_226), .A2(n_306), .B1(n_391), .B2(n_662), .Y(n_1799) );
OAI22xp33_ASAP7_75t_L g1811 ( .A1(n_226), .A2(n_306), .B1(n_1049), .B2(n_1780), .Y(n_1811) );
INVx2_ASAP7_75t_L g495 ( .A(n_227), .Y(n_495) );
INVx1_ASAP7_75t_L g555 ( .A(n_227), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g1407 ( .A(n_228), .Y(n_1407) );
INVx1_ASAP7_75t_L g673 ( .A(n_229), .Y(n_673) );
XOR2xp5_ASAP7_75t_L g852 ( .A(n_230), .B(n_853), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g1558 ( .A1(n_230), .A2(n_360), .B1(n_1538), .B2(n_1541), .Y(n_1558) );
INVx1_ASAP7_75t_L g1764 ( .A(n_231), .Y(n_1764) );
INVx1_ASAP7_75t_L g989 ( .A(n_233), .Y(n_989) );
INVx1_ASAP7_75t_L g1375 ( .A(n_234), .Y(n_1375) );
INVx1_ASAP7_75t_L g1757 ( .A(n_235), .Y(n_1757) );
INVx1_ASAP7_75t_L g1238 ( .A(n_236), .Y(n_1238) );
OAI22xp5_ASAP7_75t_L g1263 ( .A1(n_236), .A2(n_268), .B1(n_454), .B2(n_462), .Y(n_1263) );
INVx1_ASAP7_75t_L g1232 ( .A(n_237), .Y(n_1232) );
BUFx3_ASAP7_75t_L g459 ( .A(n_239), .Y(n_459) );
INVx1_ASAP7_75t_L g1007 ( .A(n_240), .Y(n_1007) );
OA211x2_ASAP7_75t_L g1022 ( .A1(n_240), .A2(n_652), .B(n_1023), .C(n_1025), .Y(n_1022) );
INVx1_ASAP7_75t_L g1369 ( .A(n_241), .Y(n_1369) );
CKINVDCx5p33_ASAP7_75t_R g1416 ( .A(n_242), .Y(n_1416) );
CKINVDCx5p33_ASAP7_75t_R g1063 ( .A(n_243), .Y(n_1063) );
CKINVDCx5p33_ASAP7_75t_R g1454 ( .A(n_244), .Y(n_1454) );
OAI22xp5_ASAP7_75t_SL g971 ( .A1(n_245), .A2(n_972), .B1(n_1018), .B2(n_1031), .Y(n_971) );
NAND4xp25_ASAP7_75t_L g972 ( .A(n_245), .B(n_973), .C(n_991), .D(n_1001), .Y(n_972) );
XOR2xp5_ASAP7_75t_L g781 ( .A(n_246), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g1010 ( .A(n_247), .Y(n_1010) );
INVx1_ASAP7_75t_L g1101 ( .A(n_248), .Y(n_1101) );
INVx1_ASAP7_75t_L g1038 ( .A(n_249), .Y(n_1038) );
OAI211xp5_ASAP7_75t_L g1043 ( .A1(n_249), .A2(n_642), .B(n_1044), .C(n_1046), .Y(n_1043) );
INVx1_ASAP7_75t_L g1243 ( .A(n_251), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_251), .B(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g563 ( .A(n_253), .Y(n_563) );
INVx1_ASAP7_75t_L g788 ( .A(n_254), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g1447 ( .A(n_255), .Y(n_1447) );
INVx1_ASAP7_75t_L g982 ( .A(n_256), .Y(n_982) );
CKINVDCx5p33_ASAP7_75t_R g1409 ( .A(n_257), .Y(n_1409) );
INVx1_ASAP7_75t_L g867 ( .A(n_258), .Y(n_867) );
INVx1_ASAP7_75t_L g1819 ( .A(n_259), .Y(n_1819) );
INVx1_ASAP7_75t_L g432 ( .A(n_260), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_261), .Y(n_1060) );
AOI221xp5_ASAP7_75t_L g1361 ( .A1(n_263), .A2(n_281), .B1(n_549), .B2(n_619), .C(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1104 ( .A(n_264), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_264), .A2(n_322), .B1(n_1126), .B2(n_1127), .Y(n_1125) );
INVx1_ASAP7_75t_L g1374 ( .A(n_265), .Y(n_1374) );
INVx1_ASAP7_75t_L g942 ( .A(n_266), .Y(n_942) );
XOR2xp5_ASAP7_75t_L g1186 ( .A(n_267), .B(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1240 ( .A(n_268), .Y(n_1240) );
BUFx3_ASAP7_75t_L g399 ( .A(n_269), .Y(n_399) );
INVx1_ASAP7_75t_L g414 ( .A(n_269), .Y(n_414) );
XOR2x2_ASAP7_75t_L g1475 ( .A(n_270), .B(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1006 ( .A(n_272), .Y(n_1006) );
INVx1_ASAP7_75t_L g1284 ( .A(n_273), .Y(n_1284) );
INVx1_ASAP7_75t_L g990 ( .A(n_274), .Y(n_990) );
INVx1_ASAP7_75t_L g936 ( .A(n_275), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_276), .A2(n_318), .B1(n_531), .B2(n_535), .Y(n_530) );
INVx1_ASAP7_75t_L g644 ( .A(n_277), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_279), .A2(n_365), .B1(n_538), .B2(n_540), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_280), .A2(n_346), .B1(n_616), .B2(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g858 ( .A(n_283), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g1155 ( .A(n_285), .Y(n_1155) );
INVx1_ASAP7_75t_L g750 ( .A(n_286), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g1221 ( .A(n_287), .B(n_454), .Y(n_1221) );
INVx1_ASAP7_75t_L g669 ( .A(n_288), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g1202 ( .A(n_290), .Y(n_1202) );
OAI22xp33_ASAP7_75t_L g1432 ( .A1(n_291), .A2(n_315), .B1(n_485), .B2(n_1185), .Y(n_1432) );
CKINVDCx5p33_ASAP7_75t_R g1158 ( .A(n_292), .Y(n_1158) );
INVx1_ASAP7_75t_L g646 ( .A(n_293), .Y(n_646) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_293), .A2(n_651), .B(n_652), .C(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g562 ( .A(n_294), .Y(n_562) );
INVx1_ASAP7_75t_L g986 ( .A(n_295), .Y(n_986) );
CKINVDCx5p33_ASAP7_75t_R g1445 ( .A(n_296), .Y(n_1445) );
INVx1_ASAP7_75t_L g461 ( .A(n_299), .Y(n_461) );
INVx1_ASAP7_75t_L g465 ( .A(n_299), .Y(n_465) );
INVx1_ASAP7_75t_L g983 ( .A(n_300), .Y(n_983) );
INVx1_ASAP7_75t_L g682 ( .A(n_301), .Y(n_682) );
INVx1_ASAP7_75t_L g739 ( .A(n_302), .Y(n_739) );
OAI211xp5_ASAP7_75t_L g887 ( .A1(n_305), .A2(n_888), .B(n_889), .C(n_890), .Y(n_887) );
INVx1_ASAP7_75t_L g905 ( .A(n_305), .Y(n_905) );
INVx1_ASAP7_75t_L g1102 ( .A(n_307), .Y(n_1102) );
INVx1_ASAP7_75t_L g1171 ( .A(n_308), .Y(n_1171) );
OAI211xp5_ASAP7_75t_SL g1177 ( .A1(n_308), .A2(n_889), .B(n_1137), .C(n_1178), .Y(n_1177) );
OAI22xp33_ASAP7_75t_L g1040 ( .A1(n_310), .A2(n_312), .B1(n_391), .B2(n_662), .Y(n_1040) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_310), .A2(n_312), .B1(n_841), .B2(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1503 ( .A(n_313), .Y(n_1503) );
AOI22xp5_ASAP7_75t_SL g1561 ( .A1(n_314), .A2(n_367), .B1(n_1534), .B2(n_1557), .Y(n_1561) );
INVx1_ASAP7_75t_L g678 ( .A(n_316), .Y(n_678) );
INVx1_ASAP7_75t_L g1287 ( .A(n_317), .Y(n_1287) );
AOI22xp33_ASAP7_75t_SL g520 ( .A1(n_318), .A2(n_355), .B1(n_515), .B2(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g1333 ( .A(n_319), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1535 ( .A(n_320), .B(n_1536), .Y(n_1535) );
INVx1_ASAP7_75t_L g1540 ( .A(n_320), .Y(n_1540) );
INVx1_ASAP7_75t_L g1091 ( .A(n_322), .Y(n_1091) );
INVx1_ASAP7_75t_L g572 ( .A(n_323), .Y(n_572) );
INVx1_ASAP7_75t_L g1377 ( .A(n_325), .Y(n_1377) );
INVx1_ASAP7_75t_L g938 ( .A(n_326), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g1410 ( .A(n_327), .Y(n_1410) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_328), .A2(n_361), .B1(n_454), .B2(n_462), .Y(n_1176) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_329), .Y(n_1054) );
INVx1_ASAP7_75t_L g949 ( .A(n_330), .Y(n_949) );
INVx1_ASAP7_75t_L g1109 ( .A(n_331), .Y(n_1109) );
CKINVDCx5p33_ASAP7_75t_R g1463 ( .A(n_332), .Y(n_1463) );
CKINVDCx5p33_ASAP7_75t_R g1249 ( .A(n_333), .Y(n_1249) );
OAI211xp5_ASAP7_75t_SL g1215 ( .A1(n_334), .A2(n_914), .B(n_1169), .C(n_1216), .Y(n_1215) );
OAI211xp5_ASAP7_75t_SL g1223 ( .A1(n_334), .A2(n_756), .B(n_889), .C(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1372 ( .A(n_335), .Y(n_1372) );
INVx1_ASAP7_75t_L g1761 ( .A(n_336), .Y(n_1761) );
INVx1_ASAP7_75t_L g1305 ( .A(n_337), .Y(n_1305) );
OAI211xp5_ASAP7_75t_L g1035 ( .A1(n_339), .A2(n_652), .B(n_704), .C(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1047 ( .A(n_339), .Y(n_1047) );
INVx1_ASAP7_75t_L g742 ( .A(n_341), .Y(n_742) );
INVx1_ASAP7_75t_L g831 ( .A(n_342), .Y(n_831) );
OAI211xp5_ASAP7_75t_L g842 ( .A1(n_342), .A2(n_642), .B(n_843), .C(n_844), .Y(n_842) );
INVx1_ASAP7_75t_L g410 ( .A(n_343), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g1161 ( .A(n_344), .Y(n_1161) );
CKINVDCx5p33_ASAP7_75t_R g1056 ( .A(n_345), .Y(n_1056) );
INVx1_ASAP7_75t_L g976 ( .A(n_347), .Y(n_976) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_348), .Y(n_395) );
INVx1_ASAP7_75t_L g1822 ( .A(n_349), .Y(n_1822) );
INVx1_ASAP7_75t_L g802 ( .A(n_351), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_352), .Y(n_1059) );
OA22x2_ASAP7_75t_L g406 ( .A1(n_353), .A2(n_407), .B1(n_556), .B2(n_557), .Y(n_406) );
INVxp67_ASAP7_75t_SL g557 ( .A(n_353), .Y(n_557) );
INVx1_ASAP7_75t_L g865 ( .A(n_354), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g1427 ( .A(n_356), .Y(n_1427) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_357), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_358), .Y(n_1194) );
XOR2x2_ASAP7_75t_L g1032 ( .A(n_362), .B(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g450 ( .A(n_363), .Y(n_450) );
INVx2_ASAP7_75t_L g504 ( .A(n_363), .Y(n_504) );
INVx1_ASAP7_75t_L g626 ( .A(n_363), .Y(n_626) );
INVx1_ASAP7_75t_L g893 ( .A(n_364), .Y(n_893) );
INVx1_ASAP7_75t_L g1015 ( .A(n_366), .Y(n_1015) );
INVx1_ASAP7_75t_L g574 ( .A(n_368), .Y(n_574) );
INVx1_ASAP7_75t_L g1823 ( .A(n_369), .Y(n_1823) );
AOI21xp33_ASAP7_75t_L g1250 ( .A1(n_370), .A2(n_609), .B(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1268 ( .A(n_370), .Y(n_1268) );
INVx1_ASAP7_75t_L g1510 ( .A(n_371), .Y(n_1510) );
INVx1_ASAP7_75t_L g1008 ( .A(n_372), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g1417 ( .A(n_373), .Y(n_1417) );
CKINVDCx5p33_ASAP7_75t_R g1236 ( .A(n_374), .Y(n_1236) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_400), .B(n_1523), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_385), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g1789 ( .A(n_379), .B(n_388), .Y(n_1789) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1793 ( .A(n_381), .B(n_384), .Y(n_1793) );
INVx1_ASAP7_75t_L g1835 ( .A(n_381), .Y(n_1835) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g1837 ( .A(n_384), .B(n_1835), .Y(n_1837) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g446 ( .A(n_388), .B(n_447), .Y(n_446) );
AOI21xp5_ASAP7_75t_SL g1229 ( .A1(n_388), .A2(n_1230), .B(n_1241), .Y(n_1229) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g523 ( .A(n_389), .B(n_399), .Y(n_523) );
AND2x4_ASAP7_75t_L g1252 ( .A(n_389), .B(n_398), .Y(n_1252) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_390), .A2(n_410), .B1(n_411), .B2(n_412), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g749 ( .A1(n_390), .A2(n_412), .B1(n_750), .B2(n_751), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_390), .A2(n_412), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
AND2x4_ASAP7_75t_SL g1788 ( .A(n_390), .B(n_1789), .Y(n_1788) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
OR2x2_ASAP7_75t_L g440 ( .A(n_392), .B(n_413), .Y(n_440) );
OR2x6_ASAP7_75t_L g659 ( .A(n_392), .B(n_413), .Y(n_659) );
BUFx4f_ASAP7_75t_L g813 ( .A(n_392), .Y(n_813) );
INVx1_ASAP7_75t_L g963 ( .A(n_392), .Y(n_963) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g581 ( .A(n_393), .Y(n_581) );
BUFx4f_ASAP7_75t_L g825 ( .A(n_393), .Y(n_825) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g415 ( .A(n_395), .B(n_416), .Y(n_415) );
NAND2x1_ASAP7_75t_L g422 ( .A(n_395), .B(n_396), .Y(n_422) );
AND2x2_ASAP7_75t_L g428 ( .A(n_395), .B(n_396), .Y(n_428) );
INVx1_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
INVx2_ASAP7_75t_L g444 ( .A(n_395), .Y(n_444) );
INVx2_ASAP7_75t_L g510 ( .A(n_395), .Y(n_510) );
INVx2_ASAP7_75t_L g416 ( .A(n_396), .Y(n_416) );
BUFx2_ASAP7_75t_L g431 ( .A(n_396), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_396), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g511 ( .A(n_396), .Y(n_511) );
AND2x2_ASAP7_75t_L g513 ( .A(n_396), .B(n_444), .Y(n_513) );
OR2x2_ASAP7_75t_L g703 ( .A(n_396), .B(n_510), .Y(n_703) );
OR2x6_ASAP7_75t_L g580 ( .A(n_397), .B(n_581), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g1235 ( .A1(n_397), .A2(n_1236), .B1(n_1237), .B2(n_1238), .Y(n_1235) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g425 ( .A(n_398), .Y(n_425) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g435 ( .A(n_399), .B(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g589 ( .A(n_399), .Y(n_589) );
XNOR2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_966), .Y(n_400) );
XNOR2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_778), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_630), .B1(n_631), .B2(n_777), .Y(n_404) );
INVx1_ASAP7_75t_L g777 ( .A(n_405), .Y(n_777) );
XNOR2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_558), .Y(n_405) );
INVx1_ASAP7_75t_L g556 ( .A(n_407), .Y(n_556) );
NAND4xp75_ASAP7_75t_L g407 ( .A(n_408), .B(n_451), .C(n_499), .D(n_527), .Y(n_407) );
AO21x1_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_417), .B(n_445), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_410), .A2(n_411), .B1(n_484), .B2(n_486), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_412), .A2(n_562), .B1(n_563), .B2(n_579), .Y(n_578) );
CKINVDCx16_ASAP7_75t_R g662 ( .A(n_412), .Y(n_662) );
INVx3_ASAP7_75t_SL g899 ( .A(n_412), .Y(n_899) );
INVx4_ASAP7_75t_L g921 ( .A(n_412), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g1323 ( .A1(n_412), .A2(n_1324), .B1(n_1325), .B2(n_1326), .Y(n_1323) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_415), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_415), .Y(n_517) );
BUFx3_ASAP7_75t_L g601 ( .A(n_415), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_439), .Y(n_417) );
OAI22xp5_ASAP7_75t_SL g995 ( .A1(n_419), .A2(n_702), .B1(n_982), .B2(n_986), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_419), .A2(n_979), .B1(n_990), .B2(n_997), .Y(n_996) );
OAI221xp5_ASAP7_75t_L g1245 ( .A1(n_419), .A2(n_523), .B1(n_997), .B2(n_1246), .C(n_1247), .Y(n_1245) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g818 ( .A(n_420), .Y(n_818) );
INVx2_ASAP7_75t_L g958 ( .A(n_420), .Y(n_958) );
INVx2_ASAP7_75t_L g1211 ( .A(n_420), .Y(n_1211) );
INVx2_ASAP7_75t_L g1519 ( .A(n_420), .Y(n_1519) );
INVx4_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx4f_ASAP7_75t_L g651 ( .A(n_421), .Y(n_651) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_421), .Y(n_730) );
BUFx4f_ASAP7_75t_L g820 ( .A(n_421), .Y(n_820) );
BUFx4f_ASAP7_75t_L g903 ( .A(n_421), .Y(n_903) );
BUFx4f_ASAP7_75t_L g1169 ( .A(n_421), .Y(n_1169) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g705 ( .A(n_422), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g743 ( .A(n_423), .B(n_744), .C(n_747), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g1328 ( .A(n_423), .B(n_1329), .C(n_1332), .Y(n_1328) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI211xp5_ASAP7_75t_L g582 ( .A1(n_424), .A2(n_583), .B(n_585), .C(n_586), .Y(n_582) );
INVx2_ASAP7_75t_L g914 ( .A(n_424), .Y(n_914) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AND2x2_ASAP7_75t_L g430 ( .A(n_425), .B(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g441 ( .A(n_425), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g653 ( .A(n_425), .B(n_519), .Y(n_653) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g584 ( .A(n_427), .Y(n_584) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_428), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B1(n_433), .B2(n_438), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_430), .A2(n_433), .B1(n_745), .B2(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g1234 ( .A(n_430), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_430), .A2(n_435), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
AOI22xp5_ASAP7_75t_L g1426 ( .A1(n_430), .A2(n_433), .B1(n_1427), .B2(n_1428), .Y(n_1426) );
AOI22xp5_ASAP7_75t_L g1462 ( .A1(n_430), .A2(n_918), .B1(n_1463), .B2(n_1464), .Y(n_1462) );
AND2x4_ASAP7_75t_L g588 ( .A(n_431), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g655 ( .A(n_431), .B(n_589), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_432), .B(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_433), .A2(n_588), .B1(n_830), .B2(n_831), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g1170 ( .A1(n_433), .A2(n_655), .B1(n_1171), .B2(n_1172), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_433), .A2(n_655), .B1(n_1389), .B2(n_1396), .Y(n_1395) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g590 ( .A(n_435), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_435), .A2(n_588), .B1(n_893), .B2(n_905), .Y(n_904) );
BUFx3_ASAP7_75t_L g918 ( .A(n_435), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g1801 ( .A1(n_435), .A2(n_588), .B1(n_1802), .B2(n_1803), .Y(n_1801) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g1316 ( .A(n_441), .Y(n_1316) );
OR2x2_ASAP7_75t_L g594 ( .A(n_442), .B(n_589), .Y(n_594) );
BUFx2_ASAP7_75t_L g700 ( .A(n_442), .Y(n_700) );
INVx8_ASAP7_75t_L g709 ( .A(n_442), .Y(n_709) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI21xp33_ASAP7_75t_L g737 ( .A1(n_445), .A2(n_738), .B(n_749), .Y(n_737) );
AOI31xp33_ASAP7_75t_SL g1107 ( .A1(n_445), .A2(n_1108), .A3(n_1111), .B(n_1116), .Y(n_1107) );
AO21x1_ASAP7_75t_L g1322 ( .A1(n_445), .A2(n_1323), .B(n_1327), .Y(n_1322) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_SL g595 ( .A(n_446), .Y(n_595) );
BUFx3_ASAP7_75t_L g836 ( .A(n_446), .Y(n_836) );
BUFx2_ASAP7_75t_L g1030 ( .A(n_446), .Y(n_1030) );
OAI31xp33_ASAP7_75t_L g1213 ( .A1(n_446), .A2(n_1214), .A3(n_1215), .B(n_1219), .Y(n_1213) );
OAI21xp5_ASAP7_75t_L g1309 ( .A1(n_446), .A2(n_1310), .B(n_1317), .Y(n_1309) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g498 ( .A(n_449), .Y(n_498) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AO21x1_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_483), .B(n_491), .Y(n_451) );
NOR3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_466), .C(n_480), .Y(n_452) );
INVx2_ASAP7_75t_SL g573 ( .A(n_454), .Y(n_573) );
BUFx2_ASAP7_75t_L g761 ( .A(n_454), .Y(n_761) );
BUFx3_ASAP7_75t_L g847 ( .A(n_454), .Y(n_847) );
OR2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_458), .Y(n_454) );
AND2x4_ASAP7_75t_L g486 ( .A(n_455), .B(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_455), .B(n_487), .Y(n_1011) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x6_ASAP7_75t_L g462 ( .A(n_456), .B(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g480 ( .A(n_456), .B(n_481), .Y(n_480) );
OR2x4_ASAP7_75t_L g485 ( .A(n_456), .B(n_458), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_456), .B(n_555), .Y(n_554) );
NAND3x1_ASAP7_75t_L g624 ( .A(n_456), .B(n_555), .C(n_625), .Y(n_624) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g475 ( .A(n_457), .Y(n_475) );
NAND2xp33_ASAP7_75t_SL g667 ( .A(n_457), .B(n_495), .Y(n_667) );
INVx2_ASAP7_75t_L g672 ( .A(n_458), .Y(n_672) );
BUFx3_ASAP7_75t_L g859 ( .A(n_458), .Y(n_859) );
BUFx4f_ASAP7_75t_L g937 ( .A(n_458), .Y(n_937) );
BUFx3_ASAP7_75t_L g1072 ( .A(n_458), .Y(n_1072) );
OR2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_459), .B(n_465), .Y(n_464) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_459), .Y(n_471) );
AND2x4_ASAP7_75t_L g481 ( .A(n_459), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g490 ( .A(n_459), .Y(n_490) );
INVx1_ASAP7_75t_L g534 ( .A(n_460), .Y(n_534) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVxp67_ASAP7_75t_L g489 ( .A(n_461), .Y(n_489) );
INVx1_ASAP7_75t_L g575 ( .A(n_462), .Y(n_575) );
INVx1_ASAP7_75t_L g637 ( .A(n_462), .Y(n_637) );
INVx2_ASAP7_75t_L g762 ( .A(n_462), .Y(n_762) );
BUFx3_ASAP7_75t_L g765 ( .A(n_463), .Y(n_765) );
INVx1_ASAP7_75t_L g797 ( .A(n_463), .Y(n_797) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g685 ( .A(n_464), .Y(n_685) );
INVx1_ASAP7_75t_L g470 ( .A(n_465), .Y(n_470) );
INVx2_ASAP7_75t_L g482 ( .A(n_465), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_467), .A2(n_936), .B1(n_937), .B2(n_938), .Y(n_935) );
OAI22xp33_ASAP7_75t_L g988 ( .A1(n_467), .A2(n_859), .B1(n_989), .B2(n_990), .Y(n_988) );
INVx1_ASAP7_75t_L g1045 ( .A(n_467), .Y(n_1045) );
OAI22xp33_ASAP7_75t_L g1090 ( .A1(n_467), .A2(n_1091), .B1(n_1092), .B2(n_1095), .Y(n_1090) );
OAI22xp33_ASAP7_75t_L g1150 ( .A1(n_467), .A2(n_937), .B1(n_1151), .B2(n_1152), .Y(n_1150) );
OAI22xp33_ASAP7_75t_L g1292 ( .A1(n_467), .A2(n_937), .B1(n_1293), .B2(n_1294), .Y(n_1292) );
OAI22xp33_ASAP7_75t_L g1456 ( .A1(n_467), .A2(n_1094), .B1(n_1444), .B2(n_1450), .Y(n_1456) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx4_ASAP7_75t_L g809 ( .A(n_468), .Y(n_809) );
INVx3_ASAP7_75t_L g978 ( .A(n_468), .Y(n_978) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g641 ( .A(n_469), .Y(n_641) );
BUFx2_ASAP7_75t_L g676 ( .A(n_469), .Y(n_676) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
BUFx2_ASAP7_75t_L g476 ( .A(n_470), .Y(n_476) );
BUFx2_ASAP7_75t_L g479 ( .A(n_471), .Y(n_479) );
AND2x4_ASAP7_75t_L g542 ( .A(n_471), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g1182 ( .A(n_471), .Y(n_1182) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_473), .A2(n_644), .B1(n_645), .B2(n_646), .Y(n_643) );
AOI22xp33_ASAP7_75t_SL g844 ( .A1(n_473), .A2(n_645), .B1(n_830), .B2(n_845), .Y(n_844) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_473), .Y(n_894) );
AOI222xp33_ASAP7_75t_L g1005 ( .A1(n_473), .A2(n_478), .B1(n_551), .B2(n_1006), .C1(n_1007), .C2(n_1008), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_473), .A2(n_645), .B1(n_1037), .B2(n_1047), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g1785 ( .A1(n_473), .A2(n_645), .B1(n_1774), .B2(n_1786), .Y(n_1785) );
AOI22xp33_ASAP7_75t_L g1809 ( .A1(n_473), .A2(n_645), .B1(n_1802), .B2(n_1810), .Y(n_1809) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_476), .Y(n_473) );
AND2x4_ASAP7_75t_L g478 ( .A(n_474), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g570 ( .A(n_474), .B(n_476), .Y(n_570) );
AND2x4_ASAP7_75t_L g645 ( .A(n_474), .B(n_479), .Y(n_645) );
AND2x2_ASAP7_75t_L g892 ( .A(n_474), .B(n_479), .Y(n_892) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND3x4_ASAP7_75t_L g528 ( .A(n_475), .B(n_495), .C(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_475), .B(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g568 ( .A(n_478), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g1224 ( .A1(n_478), .A2(n_1179), .B1(n_1217), .B2(n_1225), .Y(n_1224) );
AOI222xp33_ASAP7_75t_L g1303 ( .A1(n_478), .A2(n_570), .B1(n_769), .B2(n_1304), .C1(n_1305), .C2(n_1306), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_478), .B(n_1330), .Y(n_1339) );
AOI22xp33_ASAP7_75t_SL g1388 ( .A1(n_478), .A2(n_570), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
AOI22xp33_ASAP7_75t_SL g1436 ( .A1(n_478), .A2(n_570), .B1(n_1427), .B2(n_1437), .Y(n_1436) );
AOI22xp33_ASAP7_75t_SL g1470 ( .A1(n_478), .A2(n_570), .B1(n_1463), .B2(n_1471), .Y(n_1470) );
AOI211xp5_ASAP7_75t_L g564 ( .A1(n_480), .A2(n_565), .B(n_566), .C(n_567), .Y(n_564) );
CKINVDCx8_ASAP7_75t_R g642 ( .A(n_480), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g753 ( .A1(n_480), .A2(n_746), .B(n_754), .C(n_755), .Y(n_753) );
CKINVDCx8_ASAP7_75t_R g889 ( .A(n_480), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g1003 ( .A(n_480), .B(n_1004), .Y(n_1003) );
AOI211xp5_ASAP7_75t_L g1134 ( .A1(n_480), .A2(n_619), .B(n_1135), .C(n_1136), .Y(n_1134) );
NOR3xp33_ASAP7_75t_L g1259 ( .A(n_480), .B(n_1260), .C(n_1263), .Y(n_1259) );
NOR3xp33_ASAP7_75t_L g1337 ( .A(n_480), .B(n_1338), .C(n_1340), .Y(n_1337) );
INVx2_ASAP7_75t_L g536 ( .A(n_481), .Y(n_536) );
BUFx2_ASAP7_75t_L g551 ( .A(n_481), .Y(n_551) );
BUFx2_ASAP7_75t_L g566 ( .A(n_481), .Y(n_566) );
BUFx3_ASAP7_75t_L g619 ( .A(n_481), .Y(n_619) );
BUFx2_ASAP7_75t_L g769 ( .A(n_481), .Y(n_769) );
BUFx2_ASAP7_75t_L g1272 ( .A(n_481), .Y(n_1272) );
INVx1_ASAP7_75t_L g543 ( .A(n_482), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_484), .A2(n_486), .B1(n_562), .B2(n_563), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_484), .A2(n_486), .B1(n_1109), .B2(n_1110), .Y(n_1138) );
AOI22xp5_ASAP7_75t_L g1336 ( .A1(n_484), .A2(n_1011), .B1(n_1324), .B2(n_1326), .Y(n_1336) );
INVx2_ASAP7_75t_SL g1779 ( .A(n_484), .Y(n_1779) );
INVx2_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g758 ( .A(n_485), .Y(n_758) );
INVx1_ASAP7_75t_L g840 ( .A(n_485), .Y(n_840) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_485), .Y(n_885) );
INVx1_ASAP7_75t_L g1050 ( .A(n_485), .Y(n_1050) );
INVx2_ASAP7_75t_L g648 ( .A(n_486), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_486), .A2(n_750), .B1(n_751), .B2(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g841 ( .A(n_486), .Y(n_841) );
INVx1_ASAP7_75t_L g886 ( .A(n_486), .Y(n_886) );
INVx1_ASAP7_75t_L g924 ( .A(n_486), .Y(n_924) );
INVx1_ASAP7_75t_L g1780 ( .A(n_486), .Y(n_1780) );
INVx2_ASAP7_75t_L g539 ( .A(n_487), .Y(n_539) );
INVx1_ASAP7_75t_L g546 ( .A(n_487), .Y(n_546) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_487), .Y(n_616) );
INVx2_ASAP7_75t_L g771 ( .A(n_487), .Y(n_771) );
BUFx6f_ASAP7_75t_L g1076 ( .A(n_487), .Y(n_1076) );
INVx2_ASAP7_75t_L g1078 ( .A(n_487), .Y(n_1078) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g681 ( .A(n_488), .Y(n_681) );
BUFx8_ASAP7_75t_L g688 ( .A(n_488), .Y(n_688) );
BUFx6f_ASAP7_75t_L g793 ( .A(n_488), .Y(n_793) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
AND2x4_ASAP7_75t_L g533 ( .A(n_490), .B(n_534), .Y(n_533) );
AOI31xp33_ASAP7_75t_L g752 ( .A1(n_491), .A2(n_753), .A3(n_757), .B(n_759), .Y(n_752) );
AO21x1_ASAP7_75t_L g1335 ( .A1(n_491), .A2(n_1336), .B(n_1337), .Y(n_1335) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI31xp33_ASAP7_75t_L g634 ( .A1(n_492), .A2(n_635), .A3(n_638), .B(n_647), .Y(n_634) );
OAI31xp33_ASAP7_75t_SL g1777 ( .A1(n_492), .A2(n_1778), .A3(n_1781), .B(n_1783), .Y(n_1777) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .Y(n_492) );
AND2x2_ASAP7_75t_SL g576 ( .A(n_493), .B(n_496), .Y(n_576) );
AND2x2_ASAP7_75t_L g849 ( .A(n_493), .B(n_496), .Y(n_849) );
AND2x2_ASAP7_75t_L g931 ( .A(n_493), .B(n_496), .Y(n_931) );
AND2x4_ASAP7_75t_L g1017 ( .A(n_493), .B(n_496), .Y(n_1017) );
INVx1_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_SL g522 ( .A(n_498), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g612 ( .A(n_498), .Y(n_612) );
OR2x2_ASAP7_75t_L g666 ( .A(n_498), .B(n_667), .Y(n_666) );
AOI33xp33_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_506), .A3(n_514), .B1(n_520), .B2(n_522), .B3(n_524), .Y(n_499) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_500), .Y(n_606) );
INVx1_ASAP7_75t_L g993 ( .A(n_500), .Y(n_993) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
OAI33xp33_ASAP7_75t_L g696 ( .A1(n_501), .A2(n_697), .A3(n_701), .B1(n_706), .B2(n_707), .B3(n_710), .Y(n_696) );
INVx2_ASAP7_75t_SL g1342 ( .A(n_501), .Y(n_1342) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g724 ( .A(n_502), .Y(n_724) );
INVx2_ASAP7_75t_L g955 ( .A(n_502), .Y(n_955) );
INVx1_ASAP7_75t_L g1057 ( .A(n_502), .Y(n_1057) );
INVx2_ASAP7_75t_L g1513 ( .A(n_502), .Y(n_1513) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
OR2x6_ASAP7_75t_L g553 ( .A(n_503), .B(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g951 ( .A(n_503), .B(n_554), .Y(n_951) );
INVx1_ASAP7_75t_L g1256 ( .A(n_503), .Y(n_1256) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g529 ( .A(n_504), .Y(n_529) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g526 ( .A(n_508), .Y(n_526) );
AND2x2_ASAP7_75t_L g592 ( .A(n_508), .B(n_589), .Y(n_592) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx3_ASAP7_75t_L g605 ( .A(n_509), .Y(n_605) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g722 ( .A(n_513), .Y(n_722) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_513), .Y(n_735) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_517), .Y(n_609) );
INVx2_ASAP7_75t_L g1348 ( .A(n_517), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_518), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g1113 ( .A(n_518), .Y(n_1113) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx3_ASAP7_75t_L g521 ( .A(n_519), .Y(n_521) );
BUFx3_ASAP7_75t_L g602 ( .A(n_519), .Y(n_602) );
O2A1O1Ixp33_ASAP7_75t_L g1231 ( .A1(n_521), .A2(n_589), .B(n_1232), .C(n_1233), .Y(n_1231) );
AOI222xp33_ASAP7_75t_L g1311 ( .A1(n_521), .A2(n_655), .B1(n_918), .B2(n_1305), .C1(n_1306), .C2(n_1312), .Y(n_1311) );
INVx2_ASAP7_75t_L g710 ( .A(n_522), .Y(n_710) );
INVx2_ASAP7_75t_L g960 ( .A(n_522), .Y(n_960) );
AOI33xp33_ASAP7_75t_L g1341 ( .A1(n_522), .A2(n_1342), .A3(n_1343), .B1(n_1346), .B2(n_1350), .B3(n_1352), .Y(n_1341) );
AND2x4_ASAP7_75t_L g610 ( .A(n_523), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_523), .B(n_611), .Y(n_736) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
AOI33xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_530), .A3(n_537), .B1(n_544), .B2(n_548), .B3(n_552), .Y(n_527) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_528), .B(n_615), .C(n_618), .Y(n_614) );
INVx1_ASAP7_75t_L g1362 ( .A(n_528), .Y(n_1362) );
BUFx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g629 ( .A(n_532), .Y(n_629) );
BUFx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx8_ASAP7_75t_L g550 ( .A(n_533), .Y(n_550) );
BUFx3_ASAP7_75t_L g1271 ( .A(n_533), .Y(n_1271) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g754 ( .A(n_536), .Y(n_754) );
INVx2_ASAP7_75t_L g1358 ( .A(n_536), .Y(n_1358) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_539), .A2(n_717), .B1(n_765), .B2(n_766), .C(n_767), .Y(n_764) );
INVx2_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g547 ( .A(n_541), .Y(n_547) );
INVx5_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx12f_ASAP7_75t_L g617 ( .A(n_542), .Y(n_617) );
BUFx2_ASAP7_75t_L g1274 ( .A(n_542), .Y(n_1274) );
INVx1_ASAP7_75t_L g1180 ( .A(n_543), .Y(n_1180) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_546), .A2(n_803), .B1(n_867), .B2(n_868), .Y(n_866) );
INVx8_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g768 ( .A(n_550), .Y(n_768) );
INVx2_ASAP7_75t_L g1278 ( .A(n_550), .Y(n_1278) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI33xp33_ASAP7_75t_L g664 ( .A1(n_553), .A2(n_665), .A3(n_668), .B1(n_677), .B2(n_686), .B3(n_693), .Y(n_664) );
OAI33xp33_ASAP7_75t_L g974 ( .A1(n_553), .A2(n_665), .A3(n_975), .B1(n_980), .B2(n_984), .B3(n_988), .Y(n_974) );
OAI33xp33_ASAP7_75t_L g1282 ( .A1(n_553), .A2(n_665), .A3(n_1283), .B1(n_1286), .B2(n_1289), .B3(n_1292), .Y(n_1282) );
INVx1_ASAP7_75t_L g1359 ( .A(n_553), .Y(n_1359) );
OAI33xp33_ASAP7_75t_L g1749 ( .A1(n_553), .A2(n_665), .A3(n_1750), .B1(n_1755), .B2(n_1759), .B3(n_1762), .Y(n_1749) );
AOI221xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_576), .B1(n_577), .B2(n_595), .C(n_596), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .C(n_571), .Y(n_560) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVxp67_ASAP7_75t_L g756 ( .A(n_570), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_570), .A2(n_645), .B1(n_916), .B2(n_927), .Y(n_926) );
AOI32xp33_ASAP7_75t_L g1178 ( .A1(n_570), .A2(n_1172), .A3(n_1179), .B1(n_1181), .B2(n_1183), .Y(n_1178) );
INVxp67_ASAP7_75t_L g1262 ( .A(n_570), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_574), .B2(n_575), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_572), .A2(n_574), .B1(n_592), .B2(n_593), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g1013 ( .A1(n_573), .A2(n_840), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_573), .A2(n_762), .B1(n_1117), .B2(n_1118), .Y(n_1139) );
INVx1_ASAP7_75t_L g1782 ( .A(n_573), .Y(n_1782) );
INVx1_ASAP7_75t_L g848 ( .A(n_575), .Y(n_848) );
AOI21xp5_ASAP7_75t_L g1257 ( .A1(n_576), .A2(n_1258), .B(n_1266), .Y(n_1257) );
BUFx2_ASAP7_75t_L g1485 ( .A(n_576), .Y(n_1485) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_582), .C(n_591), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g1325 ( .A(n_580), .Y(n_1325) );
INVx2_ASAP7_75t_SL g699 ( .A(n_581), .Y(n_699) );
BUFx3_ASAP7_75t_L g881 ( .A(n_581), .Y(n_881) );
BUFx3_ASAP7_75t_L g1206 ( .A(n_581), .Y(n_1206) );
BUFx6f_ASAP7_75t_L g1300 ( .A(n_581), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_583), .B(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g1349 ( .A(n_584), .Y(n_1349) );
INVx1_ASAP7_75t_L g1351 ( .A(n_584), .Y(n_1351) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g915 ( .A1(n_588), .A2(n_916), .B1(n_917), .B2(n_918), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_588), .A2(n_1006), .B1(n_1008), .B2(n_1026), .Y(n_1025) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_588), .A2(n_918), .B1(n_1217), .B2(n_1218), .Y(n_1216) );
INVx1_ASAP7_75t_L g1237 ( .A(n_589), .Y(n_1237) );
INVx2_ASAP7_75t_L g657 ( .A(n_590), .Y(n_657) );
INVx2_ASAP7_75t_L g1026 ( .A(n_590), .Y(n_1026) );
AOI221xp5_ASAP7_75t_L g738 ( .A1(n_592), .A2(n_739), .B1(n_740), .B2(n_742), .C(n_743), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_592), .A2(n_1117), .B1(n_1118), .B2(n_1119), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_592), .A2(n_1314), .B1(n_1315), .B2(n_1316), .Y(n_1313) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_593), .Y(n_660) );
INVx1_ASAP7_75t_L g834 ( .A(n_593), .Y(n_834) );
INVx2_ASAP7_75t_L g1021 ( .A(n_593), .Y(n_1021) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g741 ( .A(n_594), .Y(n_741) );
INVx1_ASAP7_75t_L g1121 ( .A(n_594), .Y(n_1121) );
OAI31xp33_ASAP7_75t_L g649 ( .A1(n_595), .A2(n_650), .A3(n_658), .B(n_661), .Y(n_649) );
OAI31xp33_ASAP7_75t_L g897 ( .A1(n_595), .A2(n_898), .A3(n_900), .B(n_906), .Y(n_897) );
OAI31xp33_ASAP7_75t_SL g911 ( .A1(n_595), .A2(n_912), .A3(n_919), .B(n_920), .Y(n_911) );
OAI31xp33_ASAP7_75t_L g1034 ( .A1(n_595), .A2(n_1035), .A3(n_1039), .B(n_1040), .Y(n_1034) );
OAI31xp33_ASAP7_75t_L g1798 ( .A1(n_595), .A2(n_1799), .A3(n_1800), .B(n_1804), .Y(n_1798) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_597), .B(n_607), .C(n_614), .D(n_620), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_603), .C(n_606), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g720 ( .A(n_605), .Y(n_720) );
INVx2_ASAP7_75t_L g1126 ( .A(n_605), .Y(n_1126) );
INVx2_ASAP7_75t_L g1254 ( .A(n_605), .Y(n_1254) );
INVx2_ASAP7_75t_SL g1344 ( .A(n_605), .Y(n_1344) );
INVx1_ASAP7_75t_L g1353 ( .A(n_605), .Y(n_1353) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .C(n_613), .Y(n_607) );
INVx2_ASAP7_75t_L g821 ( .A(n_610), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g1064 ( .A(n_610), .Y(n_1064) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_SL g1269 ( .A(n_616), .Y(n_1269) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_619), .Y(n_929) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .C(n_627), .Y(n_620) );
INVx1_ASAP7_75t_L g805 ( .A(n_622), .Y(n_805) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx2_ASAP7_75t_L g776 ( .A(n_623), .Y(n_776) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g870 ( .A(n_624), .Y(n_870) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_711), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_649), .C(n_663), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_637), .A2(n_1010), .B1(n_1011), .B2(n_1012), .Y(n_1009) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g1784 ( .A(n_640), .Y(n_1784) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_641), .A2(n_671), .B1(n_694), .B2(n_695), .Y(n_693) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_641), .Y(n_861) );
OAI22xp33_ASAP7_75t_L g948 ( .A1(n_641), .A2(n_937), .B1(n_949), .B2(n_950), .Y(n_948) );
BUFx6f_ASAP7_75t_L g1105 ( .A(n_641), .Y(n_1105) );
OAI22xp33_ASAP7_75t_L g1159 ( .A1(n_641), .A2(n_937), .B1(n_1160), .B2(n_1161), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1201 ( .A1(n_641), .A2(n_937), .B1(n_1202), .B2(n_1203), .Y(n_1201) );
OAI22xp33_ASAP7_75t_L g1373 ( .A1(n_641), .A2(n_937), .B1(n_1374), .B2(n_1375), .Y(n_1373) );
OAI22xp33_ASAP7_75t_L g1415 ( .A1(n_641), .A2(n_1094), .B1(n_1416), .B2(n_1417), .Y(n_1415) );
OAI22xp33_ASAP7_75t_L g1459 ( .A1(n_641), .A2(n_1094), .B1(n_1445), .B2(n_1451), .Y(n_1459) );
NAND3xp33_ASAP7_75t_L g925 ( .A(n_642), .B(n_926), .C(n_928), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_644), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g1137 ( .A(n_645), .Y(n_1137) );
OAI221xp5_ASAP7_75t_L g714 ( .A1(n_651), .A2(n_715), .B1(n_717), .B2(n_718), .C(n_719), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g878 ( .A1(n_651), .A2(n_817), .B1(n_863), .B2(n_867), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g1209 ( .A1(n_651), .A2(n_957), .B1(n_1194), .B2(n_1198), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1382 ( .A1(n_651), .A2(n_702), .B1(n_1368), .B2(n_1377), .Y(n_1382) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g828 ( .A(n_653), .Y(n_828) );
AOI211xp5_ASAP7_75t_L g1111 ( .A1(n_653), .A2(n_1112), .B(n_1114), .C(n_1115), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_655), .A2(n_657), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1490 ( .A1(n_655), .A2(n_1026), .B1(n_1482), .B2(n_1491), .Y(n_1490) );
AOI22xp33_ASAP7_75t_L g1773 ( .A1(n_655), .A2(n_657), .B1(n_1774), .B2(n_1775), .Y(n_1773) );
BUFx2_ASAP7_75t_L g833 ( .A(n_659), .Y(n_833) );
BUFx6f_ASAP7_75t_L g907 ( .A(n_659), .Y(n_907) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_696), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g763 ( .A1(n_665), .A2(n_764), .B1(n_770), .B2(n_775), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g1266 ( .A1(n_665), .A2(n_869), .B1(n_1267), .B2(n_1275), .Y(n_1266) );
OAI33xp33_ASAP7_75t_L g1496 ( .A1(n_665), .A2(n_869), .A3(n_1497), .B1(n_1501), .B2(n_1504), .B3(n_1509), .Y(n_1496) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx4f_ASAP7_75t_L g785 ( .A(n_666), .Y(n_785) );
BUFx8_ASAP7_75t_L g856 ( .A(n_666), .Y(n_856) );
BUFx4f_ASAP7_75t_L g934 ( .A(n_666), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_673), .B2(n_674), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_669), .A2(n_694), .B1(n_698), .B2(n_700), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g786 ( .A1(n_670), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g806 ( .A1(n_670), .A2(n_807), .B1(n_808), .B2(n_810), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g1750 ( .A1(n_670), .A2(n_1751), .B1(n_1752), .B2(n_1753), .Y(n_1750) );
OAI22xp33_ASAP7_75t_L g1828 ( .A1(n_670), .A2(n_1434), .B1(n_1815), .B2(n_1822), .Y(n_1828) );
OAI22xp33_ASAP7_75t_L g1831 ( .A1(n_670), .A2(n_843), .B1(n_1816), .B2(n_1823), .Y(n_1831) );
BUFx4f_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_671), .A2(n_976), .B1(n_977), .B2(n_979), .Y(n_975) );
INVx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_SL g1094 ( .A(n_672), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_673), .A2(n_695), .B1(n_702), .B2(n_704), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g1762 ( .A1(n_674), .A2(n_859), .B1(n_1763), .B2(n_1764), .Y(n_1762) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_675), .Y(n_789) );
INVx1_ASAP7_75t_L g888 ( .A(n_675), .Y(n_888) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g1435 ( .A(n_676), .Y(n_1435) );
INVx1_ASAP7_75t_L g1754 ( .A(n_676), .Y(n_1754) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_682), .B2(n_683), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_678), .A2(n_689), .B1(n_702), .B2(n_704), .Y(n_701) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g1413 ( .A(n_680), .Y(n_1413) );
INVx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx2_ASAP7_75t_L g981 ( .A(n_681), .Y(n_981) );
BUFx2_ASAP7_75t_L g1276 ( .A(n_681), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_682), .A2(n_692), .B1(n_698), .B2(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_683), .A2(n_1097), .B1(n_1098), .B2(n_1099), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1289 ( .A1(n_683), .A2(n_941), .B1(n_1290), .B2(n_1291), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_683), .A2(n_1199), .B1(n_1448), .B2(n_1454), .Y(n_1458) );
INVx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g772 ( .A(n_684), .Y(n_772) );
CKINVDCx8_ASAP7_75t_R g803 ( .A(n_684), .Y(n_803) );
INVx3_ASAP7_75t_L g1196 ( .A(n_684), .Y(n_1196) );
INVx1_ASAP7_75t_L g1758 ( .A(n_684), .Y(n_1758) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g691 ( .A(n_685), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_687), .A2(n_690), .B1(n_1101), .B2(n_1102), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g1759 ( .A1(n_687), .A2(n_772), .B1(n_1760), .B2(n_1761), .Y(n_1759) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx3_ASAP7_75t_L g941 ( .A(n_688), .Y(n_941) );
INVx2_ASAP7_75t_SL g945 ( .A(n_688), .Y(n_945) );
INVx3_ASAP7_75t_L g985 ( .A(n_688), .Y(n_985) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_690), .A2(n_945), .B1(n_946), .B2(n_947), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_690), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_690), .A2(n_985), .B1(n_986), .B2(n_987), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_690), .A2(n_792), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
OAI22xp5_ASAP7_75t_L g1286 ( .A1(n_690), .A2(n_1276), .B1(n_1287), .B2(n_1288), .Y(n_1286) );
BUFx3_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g994 ( .A1(n_700), .A2(n_813), .B1(n_976), .B2(n_989), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1768 ( .A1(n_700), .A2(n_813), .B1(n_1757), .B2(n_1761), .Y(n_1768) );
OAI22xp5_ASAP7_75t_L g1422 ( .A1(n_702), .A2(n_705), .B1(n_1407), .B2(n_1417), .Y(n_1422) );
OAI22xp5_ASAP7_75t_L g1766 ( .A1(n_702), .A2(n_903), .B1(n_1756), .B2(n_1760), .Y(n_1766) );
BUFx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g716 ( .A(n_703), .Y(n_716) );
BUFx2_ASAP7_75t_L g728 ( .A(n_703), .Y(n_728) );
INVx2_ASAP7_75t_L g999 ( .A(n_703), .Y(n_999) );
BUFx3_ASAP7_75t_L g1131 ( .A(n_703), .Y(n_1131) );
OAI221xp5_ASAP7_75t_L g1123 ( .A1(n_704), .A2(n_1097), .B1(n_1101), .B2(n_1124), .C(n_1125), .Y(n_1123) );
OAI221xp5_ASAP7_75t_L g1128 ( .A1(n_704), .A2(n_1095), .B1(n_1106), .B2(n_1129), .C(n_1132), .Y(n_1128) );
INVx1_ASAP7_75t_L g1489 ( .A(n_704), .Y(n_1489) );
BUFx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_705), .A2(n_726), .B1(n_860), .B2(n_874), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_705), .A2(n_938), .B1(n_950), .B2(n_957), .Y(n_959) );
INVx2_ASAP7_75t_SL g1024 ( .A(n_705), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g1446 ( .A1(n_705), .A2(n_1421), .B1(n_1447), .B2(n_1448), .Y(n_1446) );
OAI22xp5_ASAP7_75t_L g1000 ( .A1(n_708), .A2(n_813), .B1(n_983), .B2(n_987), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1443 ( .A1(n_708), .A2(n_954), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
INVx2_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_709), .Y(n_815) );
INVx1_ASAP7_75t_L g877 ( .A(n_709), .Y(n_877) );
INVx4_ASAP7_75t_L g964 ( .A(n_709), .Y(n_964) );
INVx2_ASAP7_75t_L g1208 ( .A(n_709), .Y(n_1208) );
INVx1_ASAP7_75t_L g1381 ( .A(n_709), .Y(n_1381) );
OAI33xp33_ASAP7_75t_L g992 ( .A1(n_710), .A2(n_993), .A3(n_994), .B1(n_995), .B2(n_996), .B3(n_1000), .Y(n_992) );
OAI33xp33_ASAP7_75t_L g1418 ( .A1(n_710), .A2(n_955), .A3(n_1419), .B1(n_1420), .B2(n_1422), .B3(n_1423), .Y(n_1418) );
OAI33xp33_ASAP7_75t_L g1442 ( .A1(n_710), .A2(n_724), .A3(n_1443), .B1(n_1446), .B2(n_1449), .B3(n_1452), .Y(n_1442) );
OAI33xp33_ASAP7_75t_L g1765 ( .A1(n_710), .A2(n_955), .A3(n_1766), .B1(n_1767), .B2(n_1768), .B3(n_1769), .Y(n_1765) );
NOR4xp25_ASAP7_75t_L g712 ( .A(n_713), .B(n_737), .C(n_752), .D(n_763), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_723), .B1(n_725), .B2(n_736), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_715), .A2(n_818), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_715), .A2(n_903), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1298 ( .A1(n_715), .A2(n_730), .B1(n_1285), .B2(n_1294), .Y(n_1298) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g957 ( .A(n_716), .Y(n_957) );
OAI221xp5_ASAP7_75t_L g770 ( .A1(n_718), .A2(n_771), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_770) );
INVx3_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g1345 ( .A(n_722), .Y(n_1345) );
OAI33xp33_ASAP7_75t_L g811 ( .A1(n_723), .A2(n_812), .A3(n_816), .B1(n_819), .B2(n_821), .B3(n_822), .Y(n_811) );
OAI33xp33_ASAP7_75t_L g875 ( .A1(n_723), .A2(n_821), .A3(n_876), .B1(n_878), .B2(n_879), .B3(n_880), .Y(n_875) );
OAI33xp33_ASAP7_75t_L g1813 ( .A1(n_723), .A2(n_1064), .A3(n_1814), .B1(n_1817), .B2(n_1820), .B3(n_1824), .Y(n_1813) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI33xp33_ASAP7_75t_L g1204 ( .A1(n_724), .A2(n_960), .A3(n_1205), .B1(n_1209), .B2(n_1210), .B3(n_1212), .Y(n_1204) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_729), .B1(n_730), .B2(n_731), .C(n_732), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx4_ASAP7_75t_L g817 ( .A(n_727), .Y(n_817) );
INVx4_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_730), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g1449 ( .A1(n_730), .A2(n_1421), .B1(n_1450), .B2(n_1451), .Y(n_1449) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx2_ASAP7_75t_L g1127 ( .A(n_735), .Y(n_1127) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_739), .A2(n_742), .B1(n_760), .B2(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g1493 ( .A(n_740), .Y(n_1493) );
INVx2_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g1479 ( .A(n_758), .Y(n_1479) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g1308 ( .A(n_762), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1504 ( .A1(n_765), .A2(n_1505), .B1(n_1507), .B2(n_1508), .Y(n_1504) );
OAI22xp5_ASAP7_75t_L g1193 ( .A1(n_771), .A2(n_1194), .B1(n_1195), .B2(n_1196), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_771), .A2(n_1196), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
OAI22xp5_ASAP7_75t_L g1457 ( .A1(n_771), .A2(n_1196), .B1(n_1447), .B2(n_1453), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1197 ( .A1(n_772), .A2(n_1198), .B1(n_1199), .B2(n_1200), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1367 ( .A1(n_772), .A2(n_792), .B1(n_1368), .B2(n_1369), .Y(n_1367) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
XNOR2xp5_ASAP7_75t_L g778 ( .A(n_779), .B(n_850), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NAND3xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_826), .C(n_837), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_811), .Y(n_783) );
OAI33xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_786), .A3(n_790), .B1(n_798), .B2(n_805), .B3(n_806), .Y(n_784) );
OAI33xp33_ASAP7_75t_L g1827 ( .A1(n_785), .A2(n_869), .A3(n_1828), .B1(n_1829), .B2(n_1830), .B3(n_1831), .Y(n_1827) );
OAI22xp33_ASAP7_75t_L g812 ( .A1(n_787), .A2(n_807), .B1(n_813), .B2(n_814), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_788), .A2(n_810), .B1(n_817), .B2(n_820), .Y(n_819) );
OAI22xp33_ASAP7_75t_SL g790 ( .A1(n_791), .A2(n_792), .B1(n_794), .B2(n_795), .Y(n_790) );
OAI22xp33_ASAP7_75t_L g816 ( .A1(n_791), .A2(n_802), .B1(n_817), .B2(n_818), .Y(n_816) );
INVx2_ASAP7_75t_L g1506 ( .A(n_792), .Y(n_1506) );
INVx3_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx5_ASAP7_75t_L g801 ( .A(n_793), .Y(n_801) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_793), .Y(n_1098) );
INVx2_ASAP7_75t_SL g1199 ( .A(n_793), .Y(n_1199) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_794), .A2(n_804), .B1(n_814), .B2(n_823), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_795), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_795), .A2(n_1059), .B1(n_1066), .B2(n_1075), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_795), .A2(n_1060), .B1(n_1067), .B2(n_1078), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g1829 ( .A1(n_795), .A2(n_1199), .B1(n_1818), .B2(n_1825), .Y(n_1829) );
INVx3_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
BUFx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g943 ( .A(n_797), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_802), .B1(n_803), .B2(n_804), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx8_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx3_ASAP7_75t_L g864 ( .A(n_801), .Y(n_864) );
OAI22xp5_ASAP7_75t_L g1830 ( .A1(n_801), .A2(n_803), .B1(n_1819), .B2(n_1826), .Y(n_1830) );
OAI221xp5_ASAP7_75t_L g1275 ( .A1(n_803), .A2(n_1244), .B1(n_1249), .B2(n_1276), .C(n_1277), .Y(n_1275) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_803), .A2(n_864), .B1(n_1502), .B2(n_1503), .Y(n_1501) );
OAI33xp33_ASAP7_75t_L g1088 ( .A1(n_805), .A2(n_1089), .A3(n_1090), .B1(n_1096), .B2(n_1100), .B3(n_1103), .Y(n_1088) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_808), .A2(n_1056), .B1(n_1063), .B2(n_1081), .Y(n_1080) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g843 ( .A(n_809), .Y(n_843) );
INVx1_ASAP7_75t_L g873 ( .A(n_809), .Y(n_873) );
INVx2_ASAP7_75t_L g1261 ( .A(n_809), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g1242 ( .A1(n_813), .A2(n_814), .B1(n_1243), .B2(n_1244), .Y(n_1242) );
OAI22xp33_ASAP7_75t_L g1814 ( .A1(n_813), .A2(n_814), .B1(n_1815), .B2(n_1816), .Y(n_1814) );
OAI22xp5_ASAP7_75t_L g1824 ( .A1(n_814), .A2(n_823), .B1(n_1825), .B2(n_1826), .Y(n_1824) );
INVx5_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx6_ASAP7_75t_L g882 ( .A(n_815), .Y(n_882) );
OAI22xp5_ASAP7_75t_L g1769 ( .A1(n_817), .A2(n_1211), .B1(n_1752), .B2(n_1764), .Y(n_1769) );
OAI22xp5_ASAP7_75t_L g1817 ( .A1(n_817), .A2(n_1023), .B1(n_1818), .B2(n_1819), .Y(n_1817) );
OAI22xp5_ASAP7_75t_L g1520 ( .A1(n_818), .A2(n_997), .B1(n_1499), .B2(n_1511), .Y(n_1520) );
OAI211xp5_ASAP7_75t_SL g1248 ( .A1(n_820), .A2(n_1249), .B(n_1250), .C(n_1253), .Y(n_1248) );
OAI22xp33_ASAP7_75t_L g1820 ( .A1(n_820), .A2(n_1821), .B1(n_1822), .B2(n_1823), .Y(n_1820) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_823), .A2(n_858), .B1(n_872), .B2(n_877), .Y(n_876) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx3_ASAP7_75t_L g1055 ( .A(n_824), .Y(n_1055) );
BUFx6f_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx4_ASAP7_75t_L g954 ( .A(n_825), .Y(n_954) );
INVx3_ASAP7_75t_L g1517 ( .A(n_825), .Y(n_1517) );
OAI31xp33_ASAP7_75t_SL g826 ( .A1(n_827), .A2(n_832), .A3(n_835), .B(n_836), .Y(n_826) );
OAI31xp33_ASAP7_75t_L g1486 ( .A1(n_836), .A2(n_1487), .A3(n_1492), .B(n_1494), .Y(n_1486) );
OAI31xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_842), .A3(n_846), .B(n_849), .Y(n_837) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
HB1xp67_ASAP7_75t_L g1808 ( .A(n_843), .Y(n_1808) );
OAI31xp33_ASAP7_75t_L g883 ( .A1(n_849), .A2(n_884), .A3(n_887), .B(n_896), .Y(n_883) );
OAI31xp33_ASAP7_75t_L g1041 ( .A1(n_849), .A2(n_1042), .A3(n_1043), .B(n_1048), .Y(n_1041) );
OAI31xp33_ASAP7_75t_L g1805 ( .A1(n_849), .A2(n_1806), .A3(n_1807), .B(n_1811), .Y(n_1805) );
OAI22xp5_ASAP7_75t_L g850 ( .A1(n_851), .A2(n_908), .B1(n_909), .B2(n_965), .Y(n_850) );
INVx1_ASAP7_75t_L g965 ( .A(n_851), .Y(n_965) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND3xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_883), .C(n_897), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_875), .Y(n_854) );
OAI33xp33_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .A3(n_862), .B1(n_866), .B2(n_869), .B3(n_871), .Y(n_855) );
OAI33xp33_ASAP7_75t_L g1068 ( .A1(n_856), .A2(n_1069), .A3(n_1074), .B1(n_1077), .B2(n_1079), .B3(n_1080), .Y(n_1068) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_859), .B1(n_860), .B2(n_861), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_859), .A2(n_872), .B1(n_873), .B2(n_874), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g1497 ( .A1(n_859), .A2(n_1498), .B1(n_1499), .B2(n_1500), .Y(n_1497) );
OAI22xp33_ASAP7_75t_L g1509 ( .A1(n_859), .A2(n_1434), .B1(n_1510), .B2(n_1511), .Y(n_1509) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_865), .A2(n_868), .B1(n_881), .B2(n_882), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g1079 ( .A(n_870), .Y(n_1079) );
OAI22xp33_ASAP7_75t_L g953 ( .A1(n_877), .A2(n_936), .B1(n_949), .B2(n_954), .Y(n_953) );
OAI22xp33_ASAP7_75t_L g1053 ( .A1(n_882), .A2(n_1054), .B1(n_1055), .B2(n_1056), .Y(n_1053) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_882), .A2(n_1055), .B1(n_1066), .B2(n_1067), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1514 ( .A1(n_882), .A2(n_1498), .B1(n_1510), .B2(n_1515), .Y(n_1514) );
OAI22xp5_ASAP7_75t_L g1521 ( .A1(n_882), .A2(n_1503), .B1(n_1508), .B2(n_1515), .Y(n_1521) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_893), .B1(n_894), .B2(n_895), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g1481 ( .A1(n_891), .A2(n_894), .B1(n_1482), .B2(n_1483), .Y(n_1481) );
BUFx3_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g910 ( .A(n_911), .B(n_922), .C(n_932), .Y(n_910) );
NAND3xp33_ASAP7_75t_SL g1310 ( .A(n_914), .B(n_1311), .C(n_1313), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_917), .B(n_929), .Y(n_928) );
OAI31xp33_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_925), .A3(n_930), .B(n_931), .Y(n_922) );
OAI31xp33_ASAP7_75t_SL g1175 ( .A1(n_931), .A2(n_1176), .A3(n_1177), .B(n_1184), .Y(n_1175) );
OAI31xp33_ASAP7_75t_SL g1220 ( .A1(n_931), .A2(n_1221), .A3(n_1222), .B(n_1223), .Y(n_1220) );
OAI21xp5_ASAP7_75t_L g1301 ( .A1(n_931), .A2(n_1302), .B(n_1307), .Y(n_1301) );
OAI31xp33_ASAP7_75t_L g1385 ( .A1(n_931), .A2(n_1386), .A3(n_1387), .B(n_1391), .Y(n_1385) );
OAI31xp33_ASAP7_75t_SL g1431 ( .A1(n_931), .A2(n_1432), .A3(n_1433), .B(n_1438), .Y(n_1431) );
OAI31xp33_ASAP7_75t_SL g1467 ( .A1(n_931), .A2(n_1468), .A3(n_1469), .B(n_1472), .Y(n_1467) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_952), .Y(n_932) );
OAI33xp33_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_935), .A3(n_939), .B1(n_944), .B2(n_948), .B3(n_951), .Y(n_933) );
BUFx3_ASAP7_75t_L g1089 ( .A(n_934), .Y(n_1089) );
OAI33xp33_ASAP7_75t_L g1149 ( .A1(n_934), .A2(n_951), .A3(n_1150), .B1(n_1153), .B2(n_1156), .B3(n_1159), .Y(n_1149) );
OAI33xp33_ASAP7_75t_L g1189 ( .A1(n_934), .A2(n_951), .A3(n_1190), .B1(n_1193), .B2(n_1197), .B3(n_1201), .Y(n_1189) );
OAI33xp33_ASAP7_75t_L g1366 ( .A1(n_934), .A2(n_951), .A3(n_1367), .B1(n_1370), .B2(n_1373), .B3(n_1376), .Y(n_1366) );
OAI33xp33_ASAP7_75t_L g1404 ( .A1(n_934), .A2(n_951), .A3(n_1405), .B1(n_1408), .B2(n_1411), .B3(n_1415), .Y(n_1404) );
OAI33xp33_ASAP7_75t_L g1455 ( .A1(n_934), .A2(n_951), .A3(n_1456), .B1(n_1457), .B2(n_1458), .B3(n_1459), .Y(n_1455) );
OAI22xp5_ASAP7_75t_L g1190 ( .A1(n_937), .A2(n_977), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
OAI22xp33_ASAP7_75t_L g1283 ( .A1(n_937), .A2(n_1261), .B1(n_1284), .B2(n_1285), .Y(n_1283) );
OAI22xp5_ASAP7_75t_SL g1370 ( .A1(n_937), .A2(n_977), .B1(n_1371), .B2(n_1372), .Y(n_1370) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_937), .A2(n_977), .B1(n_1406), .B2(n_1407), .Y(n_1405) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_941), .B1(n_942), .B2(n_943), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_940), .A2(n_946), .B1(n_957), .B2(n_958), .Y(n_956) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_942), .A2(n_947), .B1(n_962), .B2(n_964), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_943), .A2(n_945), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
OAI22xp5_ASAP7_75t_L g1376 ( .A1(n_943), .A2(n_1199), .B1(n_1377), .B2(n_1378), .Y(n_1376) );
OAI22xp5_ASAP7_75t_L g1411 ( .A1(n_943), .A2(n_1412), .B1(n_1413), .B2(n_1414), .Y(n_1411) );
OAI33xp33_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_955), .A3(n_956), .B1(n_959), .B2(n_960), .B3(n_961), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_954), .A2(n_964), .B1(n_1151), .B2(n_1160), .Y(n_1163) );
OAI22xp33_ASAP7_75t_L g1380 ( .A1(n_954), .A2(n_1371), .B1(n_1374), .B2(n_1381), .Y(n_1380) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_954), .A2(n_964), .B1(n_1369), .B2(n_1378), .Y(n_1384) );
OAI22xp5_ASAP7_75t_L g1419 ( .A1(n_954), .A2(n_1207), .B1(n_1406), .B2(n_1416), .Y(n_1419) );
OAI22xp5_ASAP7_75t_L g1423 ( .A1(n_954), .A2(n_964), .B1(n_1410), .B2(n_1414), .Y(n_1423) );
OAI22xp5_ASAP7_75t_L g1452 ( .A1(n_954), .A2(n_1207), .B1(n_1453), .B2(n_1454), .Y(n_1452) );
OAI22xp5_ASAP7_75t_SL g1122 ( .A1(n_955), .A2(n_1064), .B1(n_1123), .B2(n_1128), .Y(n_1122) );
OAI33xp33_ASAP7_75t_L g1162 ( .A1(n_955), .A2(n_960), .A3(n_1163), .B1(n_1164), .B2(n_1165), .B3(n_1166), .Y(n_1162) );
OAI33xp33_ASAP7_75t_L g1295 ( .A1(n_955), .A2(n_960), .A3(n_1296), .B1(n_1297), .B2(n_1298), .B3(n_1299), .Y(n_1295) );
OAI33xp33_ASAP7_75t_L g1379 ( .A1(n_955), .A2(n_960), .A3(n_1380), .B1(n_1382), .B2(n_1383), .B3(n_1384), .Y(n_1379) );
OAI22xp5_ASAP7_75t_L g1164 ( .A1(n_957), .A2(n_958), .B1(n_1154), .B2(n_1157), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_957), .A2(n_958), .B1(n_1152), .B2(n_1161), .Y(n_1165) );
OAI22xp5_ASAP7_75t_L g1383 ( .A1(n_957), .A2(n_958), .B1(n_1372), .B2(n_1375), .Y(n_1383) );
OAI22xp5_ASAP7_75t_L g1420 ( .A1(n_958), .A2(n_1409), .B1(n_1412), .B2(n_1421), .Y(n_1420) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_962), .A2(n_964), .B1(n_1155), .B2(n_1158), .Y(n_1166) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_964), .A2(n_1195), .B1(n_1200), .B2(n_1206), .Y(n_1212) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_964), .A2(n_1206), .B1(n_1284), .B2(n_1293), .Y(n_1296) );
OAI22xp33_ASAP7_75t_L g1767 ( .A1(n_964), .A2(n_1300), .B1(n_1751), .B2(n_1763), .Y(n_1767) );
XNOR2xp5_ASAP7_75t_L g966 ( .A(n_967), .B(n_1141), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_969), .B1(n_1085), .B2(n_1140), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
AOI22xp5_ASAP7_75t_L g969 ( .A1(n_970), .A2(n_1032), .B1(n_1083), .B2(n_1084), .Y(n_969) );
INVx1_ASAP7_75t_L g1083 ( .A(n_970), .Y(n_1083) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVxp67_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
NOR4xp25_ASAP7_75t_L g1031 ( .A(n_974), .B(n_992), .C(n_1002), .D(n_1018), .Y(n_1031) );
INVx3_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
INVx2_ASAP7_75t_L g1073 ( .A(n_978), .Y(n_1073) );
INVx2_ASAP7_75t_L g1500 ( .A(n_978), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g1755 ( .A1(n_981), .A2(n_1756), .B1(n_1757), .B2(n_1758), .Y(n_1755) );
INVxp67_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g1518 ( .A1(n_997), .A2(n_1502), .B1(n_1507), .B2(n_1519), .Y(n_1518) );
INVx4_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
BUFx2_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_L g1124 ( .A(n_999), .Y(n_1124) );
INVx2_ASAP7_75t_L g1421 ( .A(n_999), .Y(n_1421) );
INVxp67_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
AOI31xp33_ASAP7_75t_L g1002 ( .A1(n_1003), .A2(n_1009), .A3(n_1013), .B(n_1016), .Y(n_1002) );
INVxp67_ASAP7_75t_SL g1004 ( .A(n_1005), .Y(n_1004) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1011), .Y(n_1185) );
AOI22xp33_ASAP7_75t_SL g1264 ( .A1(n_1011), .A2(n_1050), .B1(n_1236), .B2(n_1265), .Y(n_1264) );
AOI31xp33_ASAP7_75t_L g1133 ( .A1(n_1016), .A2(n_1134), .A3(n_1138), .B(n_1139), .Y(n_1133) );
CKINVDCx14_ASAP7_75t_R g1016 ( .A(n_1017), .Y(n_1016) );
AOI31xp67_ASAP7_75t_SL g1018 ( .A1(n_1019), .A2(n_1022), .A3(n_1027), .B(n_1029), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx5_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVxp67_ASAP7_75t_SL g1027 ( .A(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
OAI31xp33_ASAP7_75t_L g1167 ( .A1(n_1030), .A2(n_1168), .A3(n_1173), .B(n_1174), .Y(n_1167) );
OAI31xp33_ASAP7_75t_SL g1392 ( .A1(n_1030), .A2(n_1393), .A3(n_1394), .B(n_1397), .Y(n_1392) );
OAI31xp33_ASAP7_75t_L g1424 ( .A1(n_1030), .A2(n_1425), .A3(n_1429), .B(n_1430), .Y(n_1424) );
OAI31xp33_ASAP7_75t_L g1460 ( .A1(n_1030), .A2(n_1461), .A3(n_1465), .B(n_1466), .Y(n_1460) );
OAI31xp33_ASAP7_75t_L g1770 ( .A1(n_1030), .A2(n_1771), .A3(n_1772), .B(n_1776), .Y(n_1770) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1032), .Y(n_1084) );
NAND3xp33_ASAP7_75t_SL g1033 ( .A(n_1034), .B(n_1041), .C(n_1051), .Y(n_1033) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
NOR2xp33_ASAP7_75t_SL g1051 ( .A(n_1052), .B(n_1068), .Y(n_1051) );
OAI33xp33_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1057), .A3(n_1058), .B1(n_1061), .B2(n_1064), .B3(n_1065), .Y(n_1052) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_1054), .A2(n_1062), .B1(n_1070), .B2(n_1073), .Y(n_1069) );
OAI33xp33_ASAP7_75t_L g1512 ( .A1(n_1064), .A2(n_1513), .A3(n_1514), .B1(n_1518), .B2(n_1520), .B3(n_1521), .Y(n_1512) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1072), .Y(n_1082) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1085), .Y(n_1140) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
NOR4xp25_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1107), .C(n_1122), .D(n_1133), .Y(n_1087) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_1094), .Y(n_1093) );
OAI22xp33_ASAP7_75t_L g1103 ( .A1(n_1094), .A2(n_1104), .B1(n_1105), .B2(n_1106), .Y(n_1103) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1098), .Y(n_1356) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
NAND2xp5_ASAP7_75t_SL g1239 ( .A(n_1121), .B(n_1240), .Y(n_1239) );
INVx3_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_1131), .A2(n_1192), .B1(n_1203), .B2(n_1211), .Y(n_1210) );
OAI22xp5_ASAP7_75t_L g1297 ( .A1(n_1131), .A2(n_1169), .B1(n_1287), .B2(n_1290), .Y(n_1297) );
HB1xp67_ASAP7_75t_L g1821 ( .A(n_1131), .Y(n_1821) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1143), .B1(n_1474), .B2(n_1522), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
XOR2x2_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1318), .Y(n_1143) );
XNOR2xp5_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1226), .Y(n_1144) );
XNOR2xp5_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1186), .Y(n_1145) );
NAND3xp33_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1167), .C(n_1175), .Y(n_1147) );
NOR2xp33_ASAP7_75t_SL g1148 ( .A(n_1149), .B(n_1162), .Y(n_1148) );
INVx3_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
NAND3xp33_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1213), .C(n_1220), .Y(n_1187) );
NOR2xp33_ASAP7_75t_SL g1188 ( .A(n_1189), .B(n_1204), .Y(n_1188) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_1191), .A2(n_1202), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_1207), .A2(n_1288), .B1(n_1291), .B2(n_1300), .Y(n_1299) );
BUFx6f_ASAP7_75t_L g1207 ( .A(n_1208), .Y(n_1207) );
XOR2xp5_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1279), .Y(n_1226) );
OAI21xp5_ASAP7_75t_L g1228 ( .A1(n_1229), .A2(n_1255), .B(n_1257), .Y(n_1228) );
OAI21xp5_ASAP7_75t_L g1241 ( .A1(n_1242), .A2(n_1245), .B(n_1248), .Y(n_1241) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
BUFx2_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
NAND2xp5_ASAP7_75t_SL g1258 ( .A(n_1259), .B(n_1264), .Y(n_1258) );
OAI211xp5_ASAP7_75t_L g1267 ( .A1(n_1268), .A2(n_1269), .B(n_1270), .C(n_1273), .Y(n_1267) );
NAND3xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1301), .C(n_1309), .Y(n_1280) );
NOR2xp33_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1295), .Y(n_1281) );
AOI22xp5_ASAP7_75t_L g1318 ( .A1(n_1319), .A2(n_1398), .B1(n_1399), .B2(n_1473), .Y(n_1318) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1319), .Y(n_1473) );
XNOR2x1_ASAP7_75t_SL g1319 ( .A(n_1320), .B(n_1363), .Y(n_1319) );
NAND4xp75_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1335), .C(n_1341), .D(n_1354), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1334), .Y(n_1327) );
INVx2_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
AOI32xp33_ASAP7_75t_L g1354 ( .A1(n_1355), .A2(n_1357), .A3(n_1359), .B1(n_1360), .B2(n_1361), .Y(n_1354) );
AND3x1_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1385), .C(n_1392), .Y(n_1364) );
NOR2xp33_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1379), .Y(n_1365) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
XNOR2x1_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1439), .Y(n_1399) );
XNOR2xp5_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1402), .Y(n_1400) );
AND3x1_ASAP7_75t_L g1402 ( .A(n_1403), .B(n_1424), .C(n_1431), .Y(n_1402) );
NOR2xp33_ASAP7_75t_SL g1403 ( .A(n_1404), .B(n_1418), .Y(n_1403) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
AND3x1_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1460), .C(n_1467), .Y(n_1440) );
NOR2xp33_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1455), .Y(n_1441) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
HB1xp67_ASAP7_75t_L g1522 ( .A(n_1475), .Y(n_1522) );
NAND3xp33_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1486), .C(n_1495), .Y(n_1476) );
OAI31xp33_ASAP7_75t_L g1477 ( .A1(n_1478), .A2(n_1480), .A3(n_1484), .B(n_1485), .Y(n_1477) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1489), .Y(n_1488) );
NOR2xp33_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1512), .Y(n_1495) );
INVx2_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
INVx2_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVx2_ASAP7_75t_SL g1516 ( .A(n_1517), .Y(n_1516) );
OAI221xp5_ASAP7_75t_SL g1523 ( .A1(n_1524), .A2(n_1529), .B1(n_1743), .B2(n_1787), .C(n_1790), .Y(n_1523) );
INVx4_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
HB1xp67_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1528), .Y(n_1526) );
AND2x6_ASAP7_75t_L g1534 ( .A(n_1527), .B(n_1535), .Y(n_1534) );
AND2x4_ASAP7_75t_L g1538 ( .A(n_1527), .B(n_1539), .Y(n_1538) );
AND2x6_ASAP7_75t_L g1541 ( .A(n_1527), .B(n_1542), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1557 ( .A(n_1527), .B(n_1528), .Y(n_1557) );
AND2x2_ASAP7_75t_L g1571 ( .A(n_1527), .B(n_1528), .Y(n_1571) );
OAI21xp5_ASAP7_75t_L g1834 ( .A1(n_1528), .A2(n_1835), .B(n_1836), .Y(n_1834) );
AOI211xp5_ASAP7_75t_L g1529 ( .A1(n_1530), .A2(n_1543), .B(n_1625), .C(n_1737), .Y(n_1529) );
NAND2xp5_ASAP7_75t_L g1677 ( .A(n_1530), .B(n_1678), .Y(n_1677) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1530), .Y(n_1728) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
NAND3xp33_ASAP7_75t_L g1719 ( .A(n_1531), .B(n_1581), .C(n_1663), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1736 ( .A(n_1531), .B(n_1679), .Y(n_1736) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
AOI32xp33_ASAP7_75t_L g1645 ( .A1(n_1532), .A2(n_1573), .A3(n_1615), .B1(n_1646), .B2(n_1648), .Y(n_1645) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1532), .Y(n_1649) );
NOR2xp33_ASAP7_75t_L g1660 ( .A(n_1532), .B(n_1555), .Y(n_1660) );
AOI211xp5_ASAP7_75t_L g1661 ( .A1(n_1532), .A2(n_1662), .B(n_1663), .C(n_1667), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1533), .B(n_1537), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1536), .B(n_1540), .Y(n_1539) );
NAND5xp2_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1603), .C(n_1613), .D(n_1618), .E(n_1621), .Y(n_1543) );
AOI221xp5_ASAP7_75t_SL g1544 ( .A1(n_1545), .A2(n_1559), .B1(n_1566), .B2(n_1581), .C(n_1583), .Y(n_1544) );
O2A1O1Ixp33_ASAP7_75t_L g1704 ( .A1(n_1545), .A2(n_1647), .B(n_1705), .C(n_1707), .Y(n_1704) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
OR2x2_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1551), .Y(n_1546) );
NOR3xp33_ASAP7_75t_L g1688 ( .A(n_1547), .B(n_1655), .C(n_1689), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1547), .B(n_1555), .Y(n_1692) );
OAI31xp33_ASAP7_75t_L g1723 ( .A1(n_1547), .A2(n_1602), .A3(n_1724), .B(n_1726), .Y(n_1723) );
INVx3_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1582 ( .A(n_1548), .B(n_1555), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_1548), .B(n_1586), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1592 ( .A(n_1548), .B(n_1593), .Y(n_1592) );
AND2x2_ASAP7_75t_L g1604 ( .A(n_1548), .B(n_1605), .Y(n_1604) );
INVx3_ASAP7_75t_L g1679 ( .A(n_1548), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1548), .B(n_1667), .Y(n_1685) );
OR2x2_ASAP7_75t_L g1697 ( .A(n_1548), .B(n_1555), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1548), .B(n_1649), .Y(n_1700) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1548), .B(n_1710), .Y(n_1722) );
AND2x4_ASAP7_75t_SL g1548 ( .A(n_1549), .B(n_1550), .Y(n_1548) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1551), .Y(n_1637) );
OR2x2_ASAP7_75t_L g1551 ( .A(n_1552), .B(n_1555), .Y(n_1551) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1552), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1552), .B(n_1555), .Y(n_1593) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1552), .Y(n_1607) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1552), .Y(n_1662) );
NAND2xp5_ASAP7_75t_L g1552 ( .A(n_1553), .B(n_1554), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1606 ( .A(n_1555), .B(n_1607), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1556), .B(n_1558), .Y(n_1555) );
AND2x4_ASAP7_75t_L g1615 ( .A(n_1556), .B(n_1558), .Y(n_1615) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1559), .B(n_1569), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_1559), .B(n_1620), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1633 ( .A(n_1559), .B(n_1568), .Y(n_1633) );
INVx1_ASAP7_75t_L g1725 ( .A(n_1559), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1563), .Y(n_1559) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1560), .Y(n_1576) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1560), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1562), .Y(n_1560) );
OR2x2_ASAP7_75t_L g1575 ( .A(n_1563), .B(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1563), .Y(n_1590) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1563), .Y(n_1599) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1563), .B(n_1576), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1565), .Y(n_1563) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
AOI221xp5_ASAP7_75t_SL g1737 ( .A1(n_1567), .A2(n_1614), .B1(n_1637), .B2(n_1738), .C(n_1742), .Y(n_1737) );
OR2x2_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1573), .Y(n_1567) );
AND2x2_ASAP7_75t_L g1647 ( .A(n_1568), .B(n_1574), .Y(n_1647) );
AND2x2_ASAP7_75t_L g1652 ( .A(n_1568), .B(n_1608), .Y(n_1652) );
AND2x2_ASAP7_75t_L g1665 ( .A(n_1568), .B(n_1666), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1671 ( .A(n_1568), .B(n_1598), .Y(n_1671) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1568), .B(n_1716), .Y(n_1732) );
CKINVDCx5p33_ASAP7_75t_R g1568 ( .A(n_1569), .Y(n_1568) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1569), .B(n_1589), .Y(n_1588) );
NOR2xp33_ASAP7_75t_L g1617 ( .A(n_1569), .B(n_1578), .Y(n_1617) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1569), .B(n_1578), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1569), .B(n_1599), .Y(n_1622) );
OR2x2_ASAP7_75t_L g1706 ( .A(n_1569), .B(n_1590), .Y(n_1706) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1569), .B(n_1716), .Y(n_1715) );
AND2x2_ASAP7_75t_L g1569 ( .A(n_1570), .B(n_1572), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1636 ( .A(n_1570), .B(n_1572), .Y(n_1636) );
NAND2xp5_ASAP7_75t_SL g1573 ( .A(n_1574), .B(n_1577), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1574), .B(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
NOR2xp33_ASAP7_75t_L g1608 ( .A(n_1575), .B(n_1597), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1576), .B(n_1599), .Y(n_1598) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1576), .Y(n_1666) );
OAI322xp33_ASAP7_75t_L g1583 ( .A1(n_1577), .A2(n_1584), .A3(n_1587), .B1(n_1591), .B2(n_1594), .C1(n_1600), .C2(n_1602), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1577), .B(n_1601), .Y(n_1600) );
OR2x2_ASAP7_75t_L g1631 ( .A(n_1577), .B(n_1632), .Y(n_1631) );
INVx2_ASAP7_75t_L g1676 ( .A(n_1577), .Y(n_1676) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1577), .B(n_1622), .Y(n_1687) );
INVx2_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx3_ASAP7_75t_L g1597 ( .A(n_1578), .Y(n_1597) );
OR2x2_ASAP7_75t_L g1655 ( .A(n_1578), .B(n_1607), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1578 ( .A(n_1579), .B(n_1580), .Y(n_1578) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
NOR2xp33_ASAP7_75t_L g1707 ( .A(n_1582), .B(n_1708), .Y(n_1707) );
A2O1A1Ixp33_ASAP7_75t_SL g1680 ( .A1(n_1584), .A2(n_1681), .B(n_1682), .C(n_1684), .Y(n_1680) );
OAI221xp5_ASAP7_75t_L g1720 ( .A1(n_1584), .A2(n_1616), .B1(n_1702), .B2(n_1721), .C(n_1723), .Y(n_1720) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1586), .Y(n_1629) );
NAND2xp5_ASAP7_75t_L g1639 ( .A(n_1586), .B(n_1616), .Y(n_1639) );
NAND2xp5_ASAP7_75t_L g1651 ( .A(n_1586), .B(n_1652), .Y(n_1651) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1586), .Y(n_1674) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
OAI22xp5_ASAP7_75t_SL g1698 ( .A1(n_1589), .A2(n_1699), .B1(n_1701), .B2(n_1703), .Y(n_1698) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1592), .Y(n_1591) );
CKINVDCx14_ASAP7_75t_R g1602 ( .A(n_1593), .Y(n_1602) );
AOI22xp5_ASAP7_75t_L g1668 ( .A1(n_1593), .A2(n_1669), .B1(n_1674), .B2(n_1675), .Y(n_1668) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
AOI321xp33_ASAP7_75t_L g1727 ( .A1(n_1595), .A2(n_1601), .A3(n_1696), .B1(n_1728), .B2(n_1729), .C(n_1730), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1596), .B(n_1598), .Y(n_1595) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1596), .B(n_1611), .Y(n_1658) );
AOI21xp33_ASAP7_75t_L g1729 ( .A1(n_1596), .A2(n_1606), .B(n_1678), .Y(n_1729) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1596), .B(n_1629), .Y(n_1734) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1612 ( .A(n_1597), .B(n_1605), .Y(n_1612) );
NAND2xp5_ASAP7_75t_L g1624 ( .A(n_1597), .B(n_1607), .Y(n_1624) );
NAND2xp5_ASAP7_75t_L g1664 ( .A(n_1597), .B(n_1665), .Y(n_1664) );
AND2x2_ASAP7_75t_L g1673 ( .A(n_1597), .B(n_1611), .Y(n_1673) );
NOR2xp33_ASAP7_75t_L g1705 ( .A(n_1597), .B(n_1706), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1598), .B(n_1636), .Y(n_1644) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1598), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1598), .B(n_1617), .Y(n_1702) );
AOI211xp5_ASAP7_75t_L g1653 ( .A1(n_1601), .A2(n_1654), .B(n_1656), .C(n_1659), .Y(n_1653) );
NAND2xp5_ASAP7_75t_L g1742 ( .A(n_1601), .B(n_1736), .Y(n_1742) );
AOI21xp5_ASAP7_75t_L g1603 ( .A1(n_1604), .A2(n_1608), .B(n_1609), .Y(n_1603) );
INVx2_ASAP7_75t_SL g1605 ( .A(n_1606), .Y(n_1605) );
OAI22xp5_ASAP7_75t_L g1738 ( .A1(n_1606), .A2(n_1667), .B1(n_1739), .B2(n_1741), .Y(n_1738) );
AND2x2_ASAP7_75t_L g1614 ( .A(n_1607), .B(n_1615), .Y(n_1614) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1608), .Y(n_1681) );
NOR2xp33_ASAP7_75t_L g1609 ( .A(n_1610), .B(n_1612), .Y(n_1609) );
OR2x2_ASAP7_75t_L g1642 ( .A(n_1610), .B(n_1636), .Y(n_1642) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
AND2x2_ASAP7_75t_L g1616 ( .A(n_1611), .B(n_1617), .Y(n_1616) );
AND2x2_ASAP7_75t_L g1695 ( .A(n_1611), .B(n_1620), .Y(n_1695) );
AOI211xp5_ASAP7_75t_L g1714 ( .A1(n_1612), .A2(n_1678), .B(n_1715), .C(n_1717), .Y(n_1714) );
NAND2xp5_ASAP7_75t_L g1613 ( .A(n_1614), .B(n_1616), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1618 ( .A(n_1614), .B(n_1619), .Y(n_1618) );
AOI21xp5_ASAP7_75t_L g1640 ( .A1(n_1614), .A2(n_1641), .B(n_1645), .Y(n_1640) );
NAND3xp33_ASAP7_75t_L g1699 ( .A(n_1614), .B(n_1676), .C(n_1700), .Y(n_1699) );
NOR2xp33_ASAP7_75t_L g1648 ( .A(n_1615), .B(n_1649), .Y(n_1648) );
INVx2_ASAP7_75t_L g1667 ( .A(n_1615), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1708 ( .A(n_1619), .B(n_1709), .Y(n_1708) );
CKINVDCx14_ASAP7_75t_R g1726 ( .A(n_1620), .Y(n_1726) );
NAND2xp5_ASAP7_75t_L g1621 ( .A(n_1622), .B(n_1623), .Y(n_1621) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
NAND5xp2_ASAP7_75t_L g1625 ( .A(n_1626), .B(n_1704), .C(n_1711), .D(n_1720), .E(n_1727), .Y(n_1625) );
AOI321xp33_ASAP7_75t_SL g1626 ( .A1(n_1627), .A2(n_1649), .A3(n_1650), .B1(n_1677), .B2(n_1680), .C(n_1690), .Y(n_1626) );
NAND3xp33_ASAP7_75t_SL g1627 ( .A(n_1628), .B(n_1634), .C(n_1640), .Y(n_1627) );
INVxp67_ASAP7_75t_L g1741 ( .A(n_1628), .Y(n_1741) );
NAND2xp5_ASAP7_75t_L g1628 ( .A(n_1629), .B(n_1630), .Y(n_1628) );
NAND2xp5_ASAP7_75t_L g1740 ( .A(n_1629), .B(n_1656), .Y(n_1740) );
INVx1_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
A2O1A1Ixp33_ASAP7_75t_L g1690 ( .A1(n_1631), .A2(n_1639), .B(n_1691), .C(n_1693), .Y(n_1690) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
AOI21xp5_ASAP7_75t_L g1634 ( .A1(n_1635), .A2(n_1637), .B(n_1638), .Y(n_1634) );
OR2x2_ASAP7_75t_L g1657 ( .A(n_1636), .B(n_1658), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_1636), .B(n_1673), .Y(n_1683) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
NAND2xp5_ASAP7_75t_L g1641 ( .A(n_1642), .B(n_1643), .Y(n_1641) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1642), .Y(n_1712) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
A2O1A1Ixp33_ASAP7_75t_L g1650 ( .A1(n_1651), .A2(n_1653), .B(n_1661), .C(n_1668), .Y(n_1650) );
CKINVDCx14_ASAP7_75t_R g1654 ( .A(n_1655), .Y(n_1654) );
INVx1_ASAP7_75t_L g1656 ( .A(n_1657), .Y(n_1656) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1662), .B(n_1695), .Y(n_1694) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1662), .Y(n_1710) );
INVx1_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1665), .Y(n_1717) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1670), .B(n_1672), .Y(n_1669) );
INVx1_ASAP7_75t_L g1670 ( .A(n_1671), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1671), .B(n_1676), .Y(n_1675) );
INVx1_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
AOI311xp33_ASAP7_75t_L g1711 ( .A1(n_1674), .A2(n_1712), .A3(n_1713), .B(n_1714), .C(n_1718), .Y(n_1711) );
INVxp67_ASAP7_75t_SL g1713 ( .A(n_1677), .Y(n_1713) );
INVx2_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
CKINVDCx14_ASAP7_75t_R g1682 ( .A(n_1683), .Y(n_1682) );
AOI21xp5_ASAP7_75t_L g1684 ( .A1(n_1685), .A2(n_1686), .B(n_1688), .Y(n_1684) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1685), .Y(n_1703) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
NAND2xp5_ASAP7_75t_L g1724 ( .A(n_1689), .B(n_1725), .Y(n_1724) );
AOI211xp5_ASAP7_75t_L g1730 ( .A1(n_1689), .A2(n_1731), .B(n_1733), .C(n_1735), .Y(n_1730) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
AOI21xp5_ASAP7_75t_L g1693 ( .A1(n_1694), .A2(n_1696), .B(n_1698), .Y(n_1693) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
INVxp67_ASAP7_75t_SL g1718 ( .A(n_1719), .Y(n_1718) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
INVx1_ASAP7_75t_L g1731 ( .A(n_1732), .Y(n_1731) );
INVxp67_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1736), .Y(n_1735) );
INVxp67_ASAP7_75t_L g1739 ( .A(n_1740), .Y(n_1739) );
INVx1_ASAP7_75t_L g1743 ( .A(n_1744), .Y(n_1743) );
HB1xp67_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
XNOR2xp5_ASAP7_75t_L g1745 ( .A(n_1746), .B(n_1747), .Y(n_1745) );
AND3x1_ASAP7_75t_L g1747 ( .A(n_1748), .B(n_1770), .C(n_1777), .Y(n_1747) );
NOR2xp33_ASAP7_75t_SL g1748 ( .A(n_1749), .B(n_1765), .Y(n_1748) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
CKINVDCx5p33_ASAP7_75t_R g1787 ( .A(n_1788), .Y(n_1787) );
HB1xp67_ASAP7_75t_SL g1791 ( .A(n_1792), .Y(n_1791) );
BUFx3_ASAP7_75t_L g1792 ( .A(n_1793), .Y(n_1792) );
INVxp33_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
HB1xp67_ASAP7_75t_L g1796 ( .A(n_1797), .Y(n_1796) );
NAND3xp33_ASAP7_75t_L g1797 ( .A(n_1798), .B(n_1805), .C(n_1812), .Y(n_1797) );
NOR2xp33_ASAP7_75t_L g1812 ( .A(n_1813), .B(n_1827), .Y(n_1812) );
INVx1_ASAP7_75t_L g1832 ( .A(n_1833), .Y(n_1832) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
endmodule