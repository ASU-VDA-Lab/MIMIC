module real_jpeg_21403_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_0),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_65),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_53),
.B1(n_55),
.B2(n_73),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_28),
.B1(n_30),
.B2(n_73),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_73),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_47),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_4),
.A2(n_65),
.B1(n_72),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_4),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_4),
.A2(n_53),
.B1(n_55),
.B2(n_97),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_97),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_97),
.Y(n_200)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_6),
.B(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_6),
.A2(n_211),
.B(n_235),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_7),
.A2(n_65),
.B1(n_72),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_7),
.A2(n_53),
.B1(n_55),
.B2(n_77),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_77),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_77),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_54),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_54),
.Y(n_168)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_10),
.A2(n_53),
.B(n_70),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_10),
.A2(n_65),
.B1(n_72),
.B2(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_10),
.B(n_75),
.Y(n_165)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_10),
.A2(n_36),
.B(n_41),
.C(n_178),
.D(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_10),
.B(n_36),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_10),
.B(n_59),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_10),
.A2(n_26),
.B(n_193),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_L g226 ( 
.A1(n_10),
.A2(n_55),
.B(n_56),
.C(n_127),
.D(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_10),
.B(n_55),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_39),
.B1(n_53),
.B2(n_55),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_39),
.Y(n_121)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_128),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_20),
.B(n_105),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_78),
.B2(n_79),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_49),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_25),
.B(n_34),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_26),
.A2(n_27),
.B(n_32),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_26),
.A2(n_29),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_26),
.A2(n_88),
.B1(n_91),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_26),
.A2(n_27),
.B1(n_121),
.B2(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_26),
.A2(n_192),
.B(n_193),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_26),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_26),
.B(n_195),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_27),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_27),
.A2(n_200),
.B(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_30),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_28),
.A2(n_43),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_30),
.B(n_42),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_30),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_35),
.A2(n_40),
.B1(n_48),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_37),
.B1(n_57),
.B2(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_36),
.A2(n_227),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_42),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_37),
.B(n_60),
.Y(n_232)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_40),
.A2(n_46),
.B1(n_48),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_40),
.A2(n_48),
.B1(n_190),
.B2(n_225),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_40),
.A2(n_225),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_41),
.B(n_142),
.Y(n_141)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_48),
.A2(n_93),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_48),
.B(n_143),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_48),
.A2(n_141),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_48),
.B(n_118),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B1(n_59),
.B2(n_61),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_53),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_57),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_55),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_58),
.Y(n_233)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_71),
.B(n_74),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_69),
.B1(n_71),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_67),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_67),
.B(n_118),
.C(n_119),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_96),
.B(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_74),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_94),
.C(n_98),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_92),
.Y(n_137)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_91),
.B(n_118),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_104),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_101),
.A2(n_124),
.B1(n_125),
.B2(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_101),
.A2(n_102),
.B(n_149),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_109),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_106),
.B(n_108),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_110),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_122),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_112),
.B1(n_122),
.B2(n_123),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_145),
.B(n_146),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

AOI22x1_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B(n_126),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_170),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_153),
.B(n_169),
.Y(n_132)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_133),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_150),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_150),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.C(n_138),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_138),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_144),
.C(n_147),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_140),
.B1(n_147),
.B2(n_148),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_154),
.B(n_156),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_157),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_159),
.A2(n_161),
.B1(n_162),
.B2(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_159),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_163),
.A2(n_164),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_165),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_168),
.Y(n_235)
);

NOR3xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_256),
.C(n_257),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_250),
.B(n_255),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_238),
.B(n_249),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_219),
.B(n_237),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_196),
.B(n_218),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_184),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_176),
.B(n_184),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_177),
.A2(n_180),
.B1(n_181),
.B2(n_205),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_179),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_189),
.C(n_191),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_206),
.B(n_217),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_204),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_198),
.B(n_204),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_212),
.B(n_216),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_209),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_220),
.B(n_221),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_230),
.B2(n_236),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_224),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_226),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_229),
.C(n_236),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_230),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_234),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_239),
.B(n_240),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_246),
.C(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);


endmodule