module fake_jpeg_4906_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_8),
.Y(n_37)
);

OAI21xp33_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_24),
.B(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_26),
.B1(n_36),
.B2(n_39),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_47),
.B1(n_18),
.B2(n_19),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_17),
.B1(n_32),
.B2(n_25),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_51),
.B1(n_25),
.B2(n_31),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_48),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_26),
.B1(n_19),
.B2(n_31),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_16),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_26),
.B1(n_32),
.B2(n_17),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_61),
.B1(n_18),
.B2(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_64),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_56),
.Y(n_93)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_72),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_23),
.B1(n_31),
.B2(n_19),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_78),
.B1(n_84),
.B2(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_22),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_79),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_23),
.B1(n_20),
.B2(n_2),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_83),
.B1(n_21),
.B2(n_9),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_33),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_81),
.B(n_33),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_0),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_59),
.A2(n_56),
.B1(n_50),
.B2(n_58),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_20),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_52),
.Y(n_98)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_58),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_96),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_110),
.B1(n_81),
.B2(n_77),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_105),
.B1(n_67),
.B2(n_60),
.Y(n_130)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_95),
.Y(n_131)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_80),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_108),
.B1(n_71),
.B2(n_77),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_57),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_66),
.Y(n_118)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_100),
.Y(n_125)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_101),
.Y(n_121)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_79),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_50),
.B1(n_20),
.B2(n_33),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_79),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_57),
.B1(n_60),
.B2(n_21),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_118),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_80),
.B1(n_73),
.B2(n_81),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_120),
.B1(n_124),
.B2(n_132),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_73),
.B(n_66),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_115),
.A2(n_135),
.B(n_6),
.Y(n_161)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_122),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_78),
.C(n_66),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_114),
.C(n_129),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_72),
.B1(n_68),
.B2(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_74),
.B1(n_69),
.B2(n_60),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_134),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_91),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_89),
.B(n_101),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_67),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_97),
.C(n_88),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_133),
.B1(n_106),
.B2(n_103),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_88),
.B1(n_90),
.B2(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_0),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_154),
.C(n_116),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_155),
.B(n_6),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_101),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_100),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_150),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_120),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_102),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_1),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_161),
.B(n_158),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_1),
.B(n_4),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_160),
.B1(n_134),
.B2(n_112),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_5),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_112),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_5),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_161),
.A2(n_152),
.B(n_147),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_168),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_135),
.B1(n_115),
.B2(n_118),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_166),
.A2(n_169),
.B1(n_177),
.B2(n_181),
.Y(n_190)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_154),
.C(n_138),
.Y(n_187)
);

NOR2xp67_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_125),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_171),
.B(n_7),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_159),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_155),
.B1(n_146),
.B2(n_149),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_121),
.B1(n_106),
.B2(n_103),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_148),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_187),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_154),
.C(n_160),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_191),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_139),
.C(n_151),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_192),
.B(n_193),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_166),
.B(n_149),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_144),
.B1(n_137),
.B2(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_140),
.C(n_136),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_196),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_136),
.C(n_153),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_197),
.A2(n_201),
.B(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_6),
.Y(n_199)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_165),
.C(n_182),
.Y(n_201)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_207),
.B(n_215),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_172),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_213),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_186),
.C(n_191),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_198),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_216),
.A2(n_200),
.B1(n_168),
.B2(n_162),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_189),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_220),
.C(n_222),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_223),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_193),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_224),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_184),
.C(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_225),
.B(n_226),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_179),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_176),
.B1(n_181),
.B2(n_162),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_203),
.B1(n_176),
.B2(n_210),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_236),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_217),
.A2(n_210),
.B1(n_213),
.B2(n_167),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_222),
.C(n_225),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_180),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_165),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_103),
.Y(n_242)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_173),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_242),
.C(n_228),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_239),
.B(n_241),
.Y(n_247)
);

NAND2x1p5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_229),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_173),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_231),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_178),
.B(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_214),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_246),
.Y(n_251)
);

AOI322xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_248),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_14),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_7),
.Y(n_248)
);

AO21x1_ASAP7_75t_SL g249 ( 
.A1(n_247),
.A2(n_238),
.B(n_10),
.Y(n_249)
);

OAI221xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_250),
.B1(n_10),
.B2(n_11),
.C(n_14),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_252),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_251),
.A2(n_11),
.B(n_15),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_253),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g256 ( 
.A(n_255),
.Y(n_256)
);


endmodule