module fake_ibex_1991_n_1242 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_250, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1242);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_250;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1242;

wire n_1084;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_875;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_662;
wire n_979;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_257;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_795;
wire n_592;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_499;
wire n_702;
wire n_971;
wire n_451;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1190;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_695;
wire n_639;
wire n_482;
wire n_282;
wire n_870;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_749;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1129;
wire n_449;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_291;
wire n_318;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_266;
wire n_485;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1048;
wire n_774;
wire n_588;
wire n_528;
wire n_260;
wire n_836;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_996;
wire n_915;
wire n_1174;
wire n_542;
wire n_900;
wire n_377;
wire n_647;
wire n_317;
wire n_326;
wire n_270;
wire n_259;
wire n_339;
wire n_276;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_838;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_768;
wire n_839;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_277;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_782;
wire n_616;
wire n_833;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_575;
wire n_313;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_302;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_587;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_478;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_632;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_333;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_987;
wire n_750;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_581;
wire n_416;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_405;
wire n_612;
wire n_955;
wire n_440;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1016;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_493;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_565;
wire n_1123;
wire n_271;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_117),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_33),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_176),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_21),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_138),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_175),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_214),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_110),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_185),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_53),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_61),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_56),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_188),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_177),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_34),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_124),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_181),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_96),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_200),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_121),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_150),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_230),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_146),
.Y(n_281)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_91),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_126),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_198),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_228),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_61),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_144),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_192),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_233),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_209),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_196),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_17),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_9),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_247),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_94),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_158),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_203),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_191),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_56),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_123),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_139),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_72),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_119),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_132),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_187),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_50),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_104),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_141),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_64),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_183),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_109),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_226),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_211),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_99),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_105),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_134),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_222),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_178),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_128),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_253),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_224),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_57),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_234),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_37),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_204),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_207),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_206),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_202),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_133),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_223),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_145),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_120),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_113),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_142),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_210),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_122),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_225),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_221),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_11),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_199),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_216),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_251),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_25),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_245),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_149),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_152),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_160),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_190),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_88),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_205),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_115),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_112),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_217),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_240),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_157),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_55),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_66),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_213),
.Y(n_360)
);

BUFx8_ASAP7_75t_SL g361 ( 
.A(n_246),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_92),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_32),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_237),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_35),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_249),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_82),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_23),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_90),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_159),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_65),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_241),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_153),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_154),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_88),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_252),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_118),
.Y(n_377)
);

BUFx10_ASAP7_75t_L g378 ( 
.A(n_129),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_184),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_94),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_20),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_201),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_7),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_195),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_64),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_111),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_73),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_197),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_179),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_193),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_189),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_22),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_26),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_140),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_243),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_250),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_244),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_125),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_89),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_74),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_232),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_86),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_2),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_114),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_43),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_231),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_208),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_93),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_172),
.Y(n_409)
);

BUFx10_ASAP7_75t_L g410 ( 
.A(n_220),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_107),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_84),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_182),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_43),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_86),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_227),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_12),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_93),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_218),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_34),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_40),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_5),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_83),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_90),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_194),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_76),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_151),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_212),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_215),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_116),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_60),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_3),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_58),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_162),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_8),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_229),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_53),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_31),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_219),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_103),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_186),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_235),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_127),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_239),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_48),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_46),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_137),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_161),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_76),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_147),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_25),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_131),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_143),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_238),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_180),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_171),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_33),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_65),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_248),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_17),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_165),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_36),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_270),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_337),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_361),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_449),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_344),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_386),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_404),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_360),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_361),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_264),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_267),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_362),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_362),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_412),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_412),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_435),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_458),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_266),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_428),
.B(n_0),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_435),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_363),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_280),
.B(n_1),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_408),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_282),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_417),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_278),
.B(n_1),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_313),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_333),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_349),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_364),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_282),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_267),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_398),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_282),
.Y(n_497)
);

BUFx10_ASAP7_75t_L g498 ( 
.A(n_256),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_441),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_444),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_282),
.B(n_2),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_455),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_314),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_282),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_257),
.B(n_260),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_304),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_394),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_281),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_326),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_267),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_268),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_281),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_345),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_272),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_367),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_278),
.B(n_3),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_275),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_383),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_393),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_286),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_293),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_273),
.B(n_4),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_297),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_301),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_308),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_298),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_341),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_402),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_415),
.Y(n_529)
);

INVxp33_ASAP7_75t_SL g530 ( 
.A(n_351),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_298),
.B(n_4),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_525),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_514),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_483),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_477),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_465),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_471),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_478),
.Y(n_540)
);

AND2x6_ASAP7_75t_L g541 ( 
.A(n_522),
.B(n_407),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_495),
.B(n_418),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_482),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_494),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_507),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_463),
.B(n_423),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_497),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_472),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_517),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_504),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_490),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_470),
.Y(n_552)
);

OA21x2_ASAP7_75t_L g553 ( 
.A1(n_501),
.A2(n_317),
.B(n_299),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_476),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_511),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_526),
.Y(n_556)
);

NOR2x1_ASAP7_75t_L g557 ( 
.A(n_464),
.B(n_269),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_474),
.B(n_299),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_491),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_467),
.B(n_426),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_468),
.B(n_431),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_484),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_506),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_492),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_509),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_513),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_486),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_515),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_483),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_518),
.B(n_317),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_493),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_519),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_496),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_505),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_469),
.B(n_445),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_473),
.B(n_528),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_530),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_480),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_529),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_470),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_498),
.B(n_311),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_498),
.B(n_311),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_488),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_470),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_498),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_481),
.B(n_462),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_489),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_520),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_524),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_500),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_485),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_489),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_516),
.B(n_531),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_502),
.Y(n_594)
);

NAND2x1_ASAP7_75t_L g595 ( 
.A(n_516),
.B(n_277),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_508),
.B(n_273),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_531),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_499),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_512),
.B(n_283),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_521),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_510),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_523),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_527),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_503),
.B(n_285),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_466),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_479),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_R g607 ( 
.A(n_465),
.B(n_358),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_465),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_R g609 ( 
.A(n_465),
.B(n_258),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_475),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_475),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_470),
.B(n_294),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_475),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_483),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_487),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_475),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_483),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_495),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_475),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_465),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_487),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_525),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_474),
.B(n_322),
.Y(n_623)
);

BUFx8_ASAP7_75t_L g624 ( 
.A(n_525),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_474),
.B(n_322),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_498),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_475),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_463),
.A2(n_368),
.B1(n_371),
.B2(n_359),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_465),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_474),
.B(n_339),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_487),
.Y(n_631)
);

AND2x6_ASAP7_75t_L g632 ( 
.A(n_522),
.B(n_407),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_465),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_508),
.B(n_384),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_475),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_475),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_475),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_495),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_475),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_465),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_495),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_526),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_525),
.B(n_384),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_487),
.A2(n_382),
.B(n_339),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_495),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_495),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_475),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_495),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_526),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_475),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_487),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_475),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_495),
.Y(n_653)
);

BUFx10_ASAP7_75t_L g654 ( 
.A(n_555),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_SL g655 ( 
.A(n_577),
.B(n_375),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_542),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_552),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_580),
.B(n_306),
.Y(n_658)
);

INVxp67_ASAP7_75t_SL g659 ( 
.A(n_622),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_532),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_535),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_622),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_642),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_574),
.A2(n_381),
.B1(n_385),
.B2(n_380),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_591),
.B(n_259),
.Y(n_665)
);

CKINVDCx11_ASAP7_75t_R g666 ( 
.A(n_578),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_549),
.B(n_387),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_585),
.B(n_450),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_552),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_580),
.B(n_591),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_540),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_533),
.B(n_306),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_543),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_533),
.B(n_378),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_642),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_SL g677 ( 
.A1(n_536),
.A2(n_399),
.B1(n_400),
.B2(n_392),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_642),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_610),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_611),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_613),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_626),
.B(n_450),
.Y(n_682)
);

INVx4_ASAP7_75t_SL g683 ( 
.A(n_541),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_638),
.B(n_261),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_624),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_616),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_587),
.B(n_296),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_584),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_576),
.B(n_403),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_584),
.B(n_410),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_646),
.B(n_262),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_584),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_588),
.B(n_405),
.Y(n_693)
);

XNOR2xp5_ASAP7_75t_L g694 ( 
.A(n_569),
.B(n_414),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_649),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_581),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_582),
.B(n_534),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_546),
.B(n_560),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_619),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_627),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_562),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_563),
.B(n_263),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_635),
.Y(n_703)
);

INVx6_ASAP7_75t_L g704 ( 
.A(n_562),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_636),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_637),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_562),
.Y(n_707)
);

INVx8_ASAP7_75t_L g708 ( 
.A(n_541),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_618),
.B(n_378),
.Y(n_709)
);

NAND2xp33_ASAP7_75t_L g710 ( 
.A(n_541),
.B(n_265),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_567),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_641),
.B(n_448),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_565),
.B(n_271),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_538),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_567),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_639),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_554),
.B(n_324),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_558),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_643),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_603),
.B(n_292),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_566),
.B(n_274),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_567),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_641),
.B(n_410),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_644),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_645),
.B(n_289),
.Y(n_725)
);

NOR3xp33_ASAP7_75t_L g726 ( 
.A(n_545),
.B(n_420),
.C(n_365),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_568),
.B(n_276),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_628),
.B(n_421),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_546),
.B(n_422),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_586),
.B(n_279),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_572),
.B(n_284),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_589),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_632),
.B(n_287),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_647),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_650),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_645),
.B(n_295),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_648),
.B(n_395),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_579),
.B(n_288),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_556),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_553),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_632),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_539),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_628),
.B(n_424),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_608),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_553),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_586),
.B(n_290),
.Y(n_746)
);

AND3x2_ASAP7_75t_L g747 ( 
.A(n_601),
.B(n_453),
.C(n_307),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_648),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_652),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_561),
.B(n_575),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_592),
.B(n_291),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_653),
.Y(n_752)
);

AND2x2_ASAP7_75t_SL g753 ( 
.A(n_603),
.B(n_369),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_599),
.B(n_397),
.Y(n_754)
);

AND2x6_ASAP7_75t_L g755 ( 
.A(n_597),
.B(n_557),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_595),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_570),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_605),
.B(n_602),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_570),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_548),
.B(n_432),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_547),
.Y(n_761)
);

XOR2x2_ASAP7_75t_SL g762 ( 
.A(n_614),
.B(n_433),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_632),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_558),
.B(n_300),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_593),
.A2(n_369),
.B1(n_303),
.B2(n_320),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_623),
.B(n_625),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_623),
.Y(n_767)
);

BUFx10_ASAP7_75t_L g768 ( 
.A(n_620),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_615),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_621),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_631),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_651),
.Y(n_772)
);

AND2x6_ASAP7_75t_L g773 ( 
.A(n_593),
.B(n_309),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_604),
.B(n_438),
.C(n_437),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_625),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_630),
.B(n_321),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_612),
.B(n_302),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_630),
.B(n_596),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_544),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_609),
.B(n_446),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_634),
.B(n_305),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_550),
.B(n_310),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_629),
.B(n_312),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_551),
.A2(n_564),
.B1(n_571),
.B2(n_559),
.Y(n_784)
);

INVx5_ASAP7_75t_L g785 ( 
.A(n_607),
.Y(n_785)
);

INVx6_ASAP7_75t_L g786 ( 
.A(n_633),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_640),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_573),
.Y(n_788)
);

AND3x2_ASAP7_75t_L g789 ( 
.A(n_583),
.B(n_325),
.C(n_323),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_590),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_594),
.B(n_315),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_606),
.B(n_451),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_598),
.B(n_316),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_617),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_600),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_542),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_580),
.B(n_318),
.Y(n_797)
);

NOR2x1_ASAP7_75t_L g798 ( 
.A(n_585),
.B(n_332),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_585),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_638),
.Y(n_800)
);

INVx4_ASAP7_75t_SL g801 ( 
.A(n_541),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_642),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_642),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_555),
.B(n_457),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_580),
.B(n_460),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_603),
.B(n_334),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_642),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_542),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_580),
.B(n_319),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_638),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_555),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_638),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_555),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_555),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_580),
.B(n_335),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_555),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_642),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_591),
.B(n_327),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_603),
.B(n_336),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_542),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_580),
.B(n_338),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_642),
.Y(n_822)
);

INVxp67_ASAP7_75t_SL g823 ( 
.A(n_811),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_718),
.A2(n_348),
.B1(n_350),
.B2(n_346),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_757),
.B(n_328),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_759),
.B(n_329),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_773),
.A2(n_776),
.B1(n_775),
.B2(n_767),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_766),
.B(n_330),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_701),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_773),
.A2(n_370),
.B1(n_372),
.B2(n_355),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_813),
.B(n_331),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_776),
.B(n_340),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_654),
.B(n_343),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_776),
.B(n_347),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_814),
.B(n_5),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_659),
.B(n_352),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_662),
.B(n_353),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_719),
.B(n_354),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_776),
.B(n_356),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_701),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_773),
.A2(n_379),
.B1(n_389),
.B2(n_373),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_656),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_763),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_749),
.A2(n_409),
.B(n_413),
.C(n_401),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_698),
.B(n_357),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_L g846 ( 
.A(n_774),
.B(n_425),
.C(n_416),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_755),
.B(n_671),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_654),
.Y(n_848)
);

AND2x6_ASAP7_75t_SL g849 ( 
.A(n_666),
.B(n_427),
.Y(n_849)
);

NOR2x1p5_ASAP7_75t_L g850 ( 
.A(n_685),
.B(n_366),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_701),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_796),
.Y(n_852)
);

OR2x6_ASAP7_75t_L g853 ( 
.A(n_708),
.B(n_439),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_698),
.B(n_374),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_660),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_773),
.B(n_376),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_696),
.B(n_377),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_655),
.B(n_388),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_808),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_816),
.B(n_6),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_687),
.A2(n_452),
.B1(n_456),
.B2(n_442),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_720),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_657),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_657),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_687),
.A2(n_461),
.B1(n_459),
.B2(n_390),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_815),
.B(n_391),
.Y(n_866)
);

BUFx5_ASAP7_75t_L g867 ( 
.A(n_739),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_815),
.B(n_396),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_820),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_715),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_749),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_750),
.A2(n_717),
.B(n_664),
.C(n_728),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_715),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_720),
.Y(n_874)
);

AOI21x1_ASAP7_75t_L g875 ( 
.A1(n_724),
.A2(n_411),
.B(n_390),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_821),
.B(n_406),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_667),
.A2(n_689),
.B1(n_743),
.B2(n_804),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_687),
.B(n_419),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_670),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_661),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_732),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_800),
.B(n_810),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_668),
.B(n_429),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_672),
.B(n_430),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_674),
.B(n_434),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_679),
.B(n_436),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_680),
.B(n_440),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_693),
.B(n_8),
.Y(n_888)
);

BUFx8_ASAP7_75t_L g889 ( 
.A(n_790),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_681),
.B(n_443),
.Y(n_890)
);

AND2x6_ASAP7_75t_SL g891 ( 
.A(n_762),
.B(n_9),
.Y(n_891)
);

NOR2xp67_ASAP7_75t_L g892 ( 
.A(n_785),
.B(n_97),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_779),
.A2(n_753),
.B1(n_686),
.B2(n_699),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_810),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_700),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_703),
.B(n_447),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_806),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_705),
.B(n_10),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_729),
.B(n_11),
.Y(n_899)
);

NOR2xp67_ASAP7_75t_L g900 ( 
.A(n_785),
.B(n_98),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_806),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_683),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_805),
.B(n_12),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_754),
.A2(n_454),
.B1(n_342),
.B2(n_15),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_758),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_706),
.B(n_13),
.Y(n_906)
);

AND2x6_ASAP7_75t_L g907 ( 
.A(n_812),
.B(n_342),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_819),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_716),
.B(n_14),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_683),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_734),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_735),
.B(n_16),
.Y(n_912)
);

OAI221xp5_ASAP7_75t_L g913 ( 
.A1(n_726),
.A2(n_454),
.B1(n_342),
.B2(n_19),
.C(n_16),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_764),
.B(n_18),
.Y(n_914)
);

NOR2x1p5_ASAP7_75t_L g915 ( 
.A(n_742),
.B(n_18),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_740),
.A2(n_101),
.B(n_100),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_748),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_819),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_730),
.B(n_24),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_746),
.B(n_27),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_741),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_795),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_741),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_665),
.B(n_30),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_752),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_745),
.A2(n_106),
.B(n_102),
.Y(n_926)
);

AOI21xp33_ASAP7_75t_L g927 ( 
.A1(n_710),
.A2(n_31),
.B(n_35),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_697),
.B(n_36),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_739),
.Y(n_929)
);

NOR2x1p5_ASAP7_75t_L g930 ( 
.A(n_744),
.B(n_37),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_799),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_802),
.Y(n_932)
);

NAND2xp33_ASAP7_75t_L g933 ( 
.A(n_669),
.B(n_682),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_794),
.B(n_38),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_723),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_704),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_756),
.B(n_39),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_788),
.B(n_41),
.Y(n_938)
);

BUFx12f_ASAP7_75t_L g939 ( 
.A(n_714),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_761),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_769),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_770),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_780),
.B(n_42),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_771),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_787),
.B(n_44),
.Y(n_945)
);

AO22x1_ASAP7_75t_L g946 ( 
.A1(n_785),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_778),
.A2(n_51),
.B1(n_48),
.B2(n_49),
.Y(n_947)
);

BUFx4f_ASAP7_75t_SL g948 ( 
.A(n_939),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_848),
.B(n_786),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_880),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_877),
.B(n_792),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_895),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_855),
.Y(n_953)
);

CKINVDCx8_ASAP7_75t_R g954 ( 
.A(n_849),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_911),
.B(n_823),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_871),
.B(n_738),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_889),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_872),
.B(n_818),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_842),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_881),
.B(n_751),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_897),
.B(n_760),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_901),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_888),
.B(n_852),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_929),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_908),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_873),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_891),
.Y(n_967)
);

NAND2x1p5_ASAP7_75t_L g968 ( 
.A(n_862),
.B(n_688),
.Y(n_968)
);

INVx5_ASAP7_75t_L g969 ( 
.A(n_907),
.Y(n_969)
);

NOR3xp33_ASAP7_75t_SL g970 ( 
.A(n_833),
.B(n_784),
.C(n_677),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_873),
.Y(n_971)
);

BUFx8_ASAP7_75t_L g972 ( 
.A(n_945),
.Y(n_972)
);

AND2x6_ASAP7_75t_L g973 ( 
.A(n_843),
.B(n_923),
.Y(n_973)
);

BUFx4f_ASAP7_75t_L g974 ( 
.A(n_853),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_847),
.A2(n_733),
.B(n_713),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_931),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_874),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_859),
.B(n_765),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_874),
.Y(n_979)
);

NOR2xp67_ASAP7_75t_L g980 ( 
.A(n_922),
.B(n_793),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_869),
.B(n_725),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_853),
.B(n_801),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_899),
.B(n_736),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_867),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_898),
.Y(n_985)
);

AND2x4_ASAP7_75t_SL g986 ( 
.A(n_918),
.B(n_768),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_906),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_909),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_943),
.B(n_737),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_902),
.B(n_692),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_867),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_828),
.B(n_835),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_873),
.Y(n_993)
);

OR2x6_ASAP7_75t_L g994 ( 
.A(n_915),
.B(n_690),
.Y(n_994)
);

INVx3_ASAP7_75t_SL g995 ( 
.A(n_934),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_SL g996 ( 
.A1(n_928),
.A2(n_768),
.B1(n_669),
.B2(n_682),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_863),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_860),
.B(n_831),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_912),
.Y(n_999)
);

NOR3xp33_ASAP7_75t_SL g1000 ( 
.A(n_846),
.B(n_694),
.C(n_783),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_940),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_941),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_930),
.B(n_791),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_942),
.Y(n_1004)
);

OR2x6_ASAP7_75t_L g1005 ( 
.A(n_850),
.B(n_798),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_905),
.A2(n_673),
.B(n_709),
.C(n_675),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_836),
.B(n_658),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_938),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_907),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_837),
.B(n_712),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_925),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_893),
.B(n_684),
.Y(n_1012)
);

BUFx8_ASAP7_75t_L g1013 ( 
.A(n_907),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_910),
.B(n_864),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_944),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_907),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_944),
.Y(n_1017)
);

BUFx10_ASAP7_75t_L g1018 ( 
.A(n_903),
.Y(n_1018)
);

OAI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_865),
.A2(n_825),
.B1(n_826),
.B2(n_913),
.Y(n_1019)
);

AND2x6_ASAP7_75t_SL g1020 ( 
.A(n_919),
.B(n_789),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_SL g1021 ( 
.A(n_920),
.B(n_781),
.C(n_782),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_827),
.A2(n_682),
.B1(n_669),
.B2(n_772),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_865),
.B(n_691),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_845),
.B(n_747),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_879),
.B(n_777),
.Y(n_1025)
);

NOR2xp67_ASAP7_75t_L g1026 ( 
.A(n_904),
.B(n_49),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_838),
.B(n_797),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_917),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_824),
.B(n_809),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_879),
.B(n_682),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_857),
.A2(n_721),
.B1(n_727),
.B2(n_702),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_844),
.B(n_731),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_946),
.B(n_722),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_914),
.Y(n_1034)
);

OR2x6_ASAP7_75t_L g1035 ( 
.A(n_921),
.B(n_937),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_875),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_854),
.B(n_707),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_924),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_950),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_948),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_1036),
.A2(n_916),
.B(n_926),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_975),
.A2(n_840),
.B(n_829),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_951),
.A2(n_866),
.B1(n_876),
.B2(n_868),
.Y(n_1043)
);

INVx6_ASAP7_75t_L g1044 ( 
.A(n_957),
.Y(n_1044)
);

OAI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_983),
.A2(n_861),
.B(n_841),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1006),
.A2(n_830),
.B(n_883),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_958),
.A2(n_935),
.B(n_927),
.C(n_947),
.Y(n_1047)
);

AOI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_1019),
.A2(n_1007),
.B(n_1029),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_974),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_953),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_952),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1015),
.B(n_1017),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_955),
.B(n_884),
.Y(n_1053)
);

AOI211x1_ASAP7_75t_L g1054 ( 
.A1(n_992),
.A2(n_858),
.B(n_886),
.C(n_885),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_964),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_984),
.A2(n_870),
.B(n_851),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_998),
.B(n_959),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1023),
.A2(n_890),
.B(n_887),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_973),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_981),
.A2(n_896),
.B(n_856),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_956),
.A2(n_989),
.B(n_1032),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_1012),
.A2(n_933),
.B(n_932),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_1026),
.A2(n_900),
.B(n_892),
.C(n_894),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_986),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_966),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1001),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1010),
.A2(n_878),
.B(n_834),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_1034),
.A2(n_676),
.A3(n_678),
.B(n_663),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_976),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_996),
.A2(n_839),
.B1(n_832),
.B2(n_932),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_SL g1071 ( 
.A1(n_1022),
.A2(n_900),
.B(n_892),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_949),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_949),
.Y(n_1073)
);

AOI31xp67_ASAP7_75t_L g1074 ( 
.A1(n_1031),
.A2(n_803),
.A3(n_807),
.B(n_695),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1038),
.A2(n_932),
.B(n_882),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_1013),
.Y(n_1076)
);

NAND2x1_ASAP7_75t_L g1077 ( 
.A(n_973),
.B(n_936),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1002),
.Y(n_1078)
);

AO31x2_ASAP7_75t_L g1079 ( 
.A1(n_985),
.A2(n_822),
.A3(n_711),
.B(n_817),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1004),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_960),
.B(n_1011),
.Y(n_1081)
);

INVx3_ASAP7_75t_SL g1082 ( 
.A(n_967),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_977),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_987),
.A2(n_988),
.A3(n_999),
.B(n_991),
.Y(n_1084)
);

NAND2x1_ASAP7_75t_L g1085 ( 
.A(n_973),
.B(n_108),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_982),
.B(n_991),
.Y(n_1086)
);

OA22x2_ASAP7_75t_L g1087 ( 
.A1(n_994),
.A2(n_55),
.B1(n_52),
.B2(n_54),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_963),
.B(n_1003),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_966),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_962),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1033),
.A2(n_58),
.B1(n_54),
.B2(n_57),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1033),
.A2(n_62),
.B1(n_59),
.B2(n_60),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_SL g1093 ( 
.A1(n_1008),
.A2(n_63),
.B(n_66),
.Y(n_1093)
);

BUFx2_ASAP7_75t_SL g1094 ( 
.A(n_1040),
.Y(n_1094)
);

INVx6_ASAP7_75t_L g1095 ( 
.A(n_1059),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_1059),
.B(n_969),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1042),
.A2(n_1028),
.B(n_997),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1048),
.A2(n_1035),
.B(n_995),
.C(n_1027),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1052),
.A2(n_1035),
.B1(n_994),
.B2(n_1016),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1045),
.A2(n_972),
.B1(n_1018),
.B2(n_961),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1050),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_1083),
.Y(n_1102)
);

AO21x2_ASAP7_75t_L g1103 ( 
.A1(n_1041),
.A2(n_1071),
.B(n_1046),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1039),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1061),
.B(n_978),
.Y(n_1105)
);

AOI21xp33_ASAP7_75t_L g1106 ( 
.A1(n_1070),
.A2(n_1037),
.B(n_1016),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1043),
.A2(n_1058),
.B(n_1053),
.C(n_1060),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1055),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1051),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1084),
.B(n_1025),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_SL g1111 ( 
.A1(n_1087),
.A2(n_972),
.B1(n_979),
.B2(n_977),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1081),
.B(n_1088),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_1047),
.A2(n_1063),
.A3(n_1062),
.B(n_1074),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_1065),
.Y(n_1114)
);

AO31x2_ASAP7_75t_L g1115 ( 
.A1(n_1075),
.A2(n_1009),
.A3(n_979),
.B(n_1024),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_1049),
.B(n_1059),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1054),
.A2(n_1091),
.B1(n_1092),
.B2(n_1057),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_1076),
.B(n_1009),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1086),
.B(n_1014),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1049),
.B(n_1020),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1080),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1066),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1056),
.A2(n_990),
.B(n_968),
.Y(n_1123)
);

BUFx4f_ASAP7_75t_SL g1124 ( 
.A(n_1082),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1084),
.B(n_1021),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1086),
.B(n_1078),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1084),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1067),
.A2(n_1005),
.B1(n_965),
.B2(n_980),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1127),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1110),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1097),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1110),
.B(n_1079),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1119),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1112),
.B(n_1090),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1107),
.B(n_1069),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_SL g1136 ( 
.A(n_1111),
.B(n_954),
.C(n_1064),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_1115),
.B(n_1079),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1122),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1099),
.A2(n_1093),
.B1(n_1072),
.B2(n_1073),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1104),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1100),
.B(n_970),
.C(n_1000),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_1095),
.Y(n_1142)
);

CKINVDCx16_ASAP7_75t_R g1143 ( 
.A(n_1094),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_SL g1144 ( 
.A1(n_1117),
.A2(n_1044),
.B1(n_969),
.B2(n_1030),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1121),
.B(n_1068),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1109),
.B(n_1068),
.Y(n_1146)
);

BUFx12f_ASAP7_75t_L g1147 ( 
.A(n_1124),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1120),
.B(n_1126),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1108),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1135),
.A2(n_1106),
.B(n_1098),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1129),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1141),
.A2(n_1125),
.B1(n_1106),
.B2(n_1126),
.Y(n_1152)
);

CKINVDCx8_ASAP7_75t_R g1153 ( 
.A(n_1143),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1138),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_L g1155 ( 
.A(n_1144),
.B(n_1128),
.C(n_1125),
.Y(n_1155)
);

OAI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1143),
.A2(n_1118),
.B1(n_1102),
.B2(n_1116),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1146),
.B(n_1103),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1132),
.B(n_1115),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1136),
.A2(n_1101),
.B1(n_1105),
.B2(n_1102),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1140),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1130),
.B(n_1103),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_1147),
.Y(n_1162)
);

AOI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1139),
.A2(n_1077),
.B(n_1085),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1133),
.A2(n_1123),
.B1(n_1014),
.B2(n_1114),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1138),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1134),
.A2(n_1096),
.B1(n_1065),
.B2(n_1089),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1145),
.B(n_1115),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1154),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1151),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1167),
.B(n_1132),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1167),
.B(n_1132),
.Y(n_1171)
);

AO31x2_ASAP7_75t_L g1172 ( 
.A1(n_1150),
.A2(n_1165),
.A3(n_1160),
.B(n_1131),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1157),
.B(n_1137),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1153),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1161),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1161),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1162),
.B(n_1148),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1157),
.B(n_1137),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_1158),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1158),
.B(n_1137),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1158),
.Y(n_1181)
);

OA21x2_ASAP7_75t_L g1182 ( 
.A1(n_1181),
.A2(n_1152),
.B(n_1155),
.Y(n_1182)
);

AO21x2_ASAP7_75t_L g1183 ( 
.A1(n_1174),
.A2(n_1156),
.B(n_1163),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1173),
.B(n_1159),
.Y(n_1184)
);

AO21x2_ASAP7_75t_L g1185 ( 
.A1(n_1181),
.A2(n_1166),
.B(n_1131),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1168),
.B(n_1149),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1179),
.A2(n_1142),
.B1(n_1164),
.B2(n_1162),
.Y(n_1187)
);

BUFx5_ASAP7_75t_L g1188 ( 
.A(n_1169),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1184),
.B(n_1173),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1188),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1188),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1188),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1182),
.B(n_1178),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1185),
.B(n_1180),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1186),
.B(n_1170),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1188),
.B(n_1170),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1188),
.B(n_1171),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1183),
.B(n_1175),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1187),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1193),
.B(n_1175),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1193),
.B(n_1176),
.Y(n_1201)
);

INVxp67_ASAP7_75t_SL g1202 ( 
.A(n_1198),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1200),
.B(n_1199),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1201),
.B(n_1199),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1202),
.B(n_1194),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1205),
.Y(n_1206)
);

OAI32xp33_ASAP7_75t_L g1207 ( 
.A1(n_1206),
.A2(n_1198),
.A3(n_1204),
.B1(n_1203),
.B2(n_1177),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1206),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1207),
.Y(n_1209)
);

INVxp33_ASAP7_75t_L g1210 ( 
.A(n_1208),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1210),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1209),
.A2(n_1189),
.B1(n_1197),
.B2(n_1196),
.Y(n_1212)
);

AOI211xp5_ASAP7_75t_L g1213 ( 
.A1(n_1211),
.A2(n_1191),
.B(n_1192),
.C(n_1190),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1212),
.B(n_1195),
.Y(n_1214)
);

NAND5xp2_ASAP7_75t_L g1215 ( 
.A(n_1211),
.B(n_67),
.C(n_68),
.D(n_69),
.E(n_70),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1211),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1216)
);

AOI321xp33_ASAP7_75t_L g1217 ( 
.A1(n_1211),
.A2(n_75),
.A3(n_77),
.B1(n_78),
.B2(n_79),
.C(n_80),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1216),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1217),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1214),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1215),
.B(n_81),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1213),
.B(n_85),
.Y(n_1222)
);

AND3x4_ASAP7_75t_L g1223 ( 
.A(n_1213),
.B(n_85),
.C(n_87),
.Y(n_1223)
);

OAI22x1_ASAP7_75t_L g1224 ( 
.A1(n_1219),
.A2(n_1223),
.B1(n_1218),
.B2(n_1221),
.Y(n_1224)
);

NOR2x1_ASAP7_75t_L g1225 ( 
.A(n_1222),
.B(n_95),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1220),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1224),
.A2(n_993),
.B(n_971),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1226),
.B(n_1172),
.Y(n_1228)
);

AND4x1_ASAP7_75t_L g1229 ( 
.A(n_1225),
.B(n_130),
.C(n_135),
.D(n_136),
.Y(n_1229)
);

CKINVDCx12_ASAP7_75t_R g1230 ( 
.A(n_1229),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1227),
.B(n_148),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1228),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1230),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1232),
.B(n_1231),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1234),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1235),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1236),
.B(n_1233),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1237),
.Y(n_1238)
);

OAI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1238),
.A2(n_1113),
.B1(n_155),
.B2(n_156),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1238),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_1240)
);

AOI221xp5_ASAP7_75t_L g1241 ( 
.A1(n_1239),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.C(n_170),
.Y(n_1241)
);

AOI211xp5_ASAP7_75t_L g1242 ( 
.A1(n_1241),
.A2(n_1240),
.B(n_173),
.C(n_174),
.Y(n_1242)
);


endmodule