module fake_jpeg_9440_n_94 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_94);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_94;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_62;
wire n_43;
wire n_82;

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

CKINVDCx9p33_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_4),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_6),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_7),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_52),
.C(n_47),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_45),
.B1(n_57),
.B2(n_49),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_8),
.B1(n_14),
.B2(n_15),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_76),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_56),
.C(n_54),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_77),
.Y(n_81)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_73),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_79),
.A2(n_74),
.B(n_70),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g84 ( 
.A(n_82),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_81),
.B1(n_83),
.B2(n_80),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_87),
.A2(n_71),
.B1(n_20),
.B2(n_21),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_26),
.B(n_28),
.Y(n_90)
);

OAI321xp33_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_30),
.A3(n_31),
.B1(n_32),
.B2(n_34),
.C(n_35),
.Y(n_91)
);

OAI21x1_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_36),
.B(n_37),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_38),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_39),
.Y(n_94)
);


endmodule