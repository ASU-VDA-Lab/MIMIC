module real_jpeg_24762_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_0),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_0),
.B(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_0),
.B(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_2),
.B(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_2),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_2),
.B(n_114),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_2),
.B(n_74),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_2),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_2),
.B(n_30),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_2),
.B(n_25),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_3),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_3),
.B(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_3),
.B(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_3),
.B(n_56),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_3),
.B(n_34),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_3),
.B(n_30),
.Y(n_241)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_3),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_3),
.B(n_217),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_6),
.B(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_6),
.B(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_6),
.B(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_6),
.B(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_6),
.B(n_34),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_6),
.B(n_30),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_6),
.B(n_25),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_6),
.B(n_217),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_9),
.B(n_34),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_9),
.B(n_30),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_9),
.B(n_56),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_9),
.B(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_9),
.B(n_25),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_37),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_10),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_10),
.B(n_114),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_10),
.B(n_74),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_10),
.B(n_34),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_10),
.B(n_30),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_11),
.B(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_34),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_11),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_11),
.B(n_114),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_11),
.B(n_74),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_11),
.B(n_56),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_12),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_12),
.B(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_12),
.B(n_74),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_12),
.B(n_56),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_12),
.B(n_34),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_12),
.B(n_30),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_12),
.B(n_217),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_15),
.B(n_30),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_15),
.B(n_211),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_15),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_15),
.B(n_74),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_15),
.B(n_56),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_15),
.B(n_34),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_16),
.B(n_56),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_16),
.B(n_34),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_16),
.B(n_74),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_16),
.B(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_16),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_30),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_16),
.B(n_25),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_16),
.B(n_217),
.Y(n_257)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_17),
.Y(n_111)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_17),
.Y(n_159)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_17),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_82),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_58),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_45),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_35),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_28),
.C(n_33),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_23),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_26),
.B(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_26),
.B(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_29),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_29),
.B1(n_33),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_52),
.C(n_54),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_33),
.A2(n_49),
.B1(n_54),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_34),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_40),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_44),
.B(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_44),
.B(n_253),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.C(n_51),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_51),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_53),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_71),
.C(n_73),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_54),
.A2(n_73),
.B1(n_78),
.B2(n_332),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_55),
.B(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_55),
.B(n_72),
.Y(n_265)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.C(n_80),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_59),
.B(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_70),
.C(n_76),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_60),
.B(n_376),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_61),
.B(n_80),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_63),
.CI(n_64),
.CON(n_61),
.SN(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.C(n_68),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_65),
.B(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_70),
.B(n_76),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_71),
.B(n_357),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_73),
.A2(n_303),
.B1(n_304),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_73),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_SL g361 ( 
.A(n_73),
.B(n_303),
.C(n_330),
.Y(n_361)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_380),
.C(n_381),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_371),
.C(n_372),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_349),
.C(n_350),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_325),
.C(n_326),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_293),
.C(n_294),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_259),
.C(n_260),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_223),
.C(n_224),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_190),
.C(n_191),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_164),
.C(n_165),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_125),
.C(n_136),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_106),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_94),
.B(n_101),
.C(n_106),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_99),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_96),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_102),
.B(n_104),
.C(n_105),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_116),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_107),
.B(n_117),
.C(n_118),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_114),
.Y(n_253)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_120),
.B(n_124),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_135),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_130),
.B1(n_135),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_160),
.C(n_161),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.C(n_150),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_143),
.C(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.C(n_155),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_153),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_179),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_180),
.C(n_189),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_175),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.C(n_175),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_170),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_173),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g384 ( 
.A(n_175),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_177),
.CI(n_178),
.CON(n_175),
.SN(n_175)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_177),
.C(n_178),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_187),
.B2(n_188),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_183),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_206),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_195),
.C(n_206),
.Y(n_223)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_202),
.C(n_205),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_197),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.CI(n_200),
.CON(n_197),
.SN(n_197)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_199),
.C(n_200),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_214),
.C(n_221),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_214),
.B1(n_221),
.B2(n_222),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_212),
.B(n_213),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_212),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_248),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_213),
.B(n_248),
.C(n_249),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_219),
.C(n_220),
.Y(n_243)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_244),
.B2(n_258),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_245),
.C(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_229),
.C(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_237),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_233),
.C(n_236),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_235),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_244),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_250),
.B(n_289),
.C(n_290),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_254),
.CI(n_257),
.CON(n_250),
.SN(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_291),
.B2(n_292),
.Y(n_260)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_283),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_283),
.C(n_291),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_264),
.B(n_272),
.C(n_273),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_265),
.B(n_267),
.C(n_269),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_282),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_274),
.Y(n_282)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_277),
.A2(n_278),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_281),
.C(n_282),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_277),
.B(n_300),
.C(n_303),
.Y(n_347)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_286),
.C(n_287),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_297),
.C(n_324),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_311),
.B2(n_324),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_305),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_306),
.C(n_307),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_303),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g385 ( 
.A(n_307),
.Y(n_385)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_309),
.CI(n_310),
.CON(n_307),
.SN(n_307)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_309),
.C(n_310),
.Y(n_334)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_314),
.C(n_315),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_323),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_319),
.C(n_321),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_318),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_319),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_320),
.A2(n_321),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_346),
.C(n_347),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_348),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_339),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_339),
.C(n_348),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_334),
.C(n_335),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g386 ( 
.A(n_335),
.Y(n_386)
);

FAx1_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.CI(n_338),
.CON(n_335),
.SN(n_335)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_337),
.C(n_338),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_342),
.C(n_343),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_345),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_353),
.C(n_363),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_362),
.B2(n_363),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_358),
.B2(n_359),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_360),
.C(n_361),
.Y(n_374)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_366),
.C(n_369),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_368),
.B2(n_369),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_369),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_372)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_373),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_374),
.B(n_375),
.C(n_379),
.Y(n_380)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);


endmodule