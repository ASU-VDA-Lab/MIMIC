module fake_jpeg_15441_n_163 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_54),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_49),
.B1(n_65),
.B2(n_56),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_84),
.B1(n_89),
.B2(n_92),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_52),
.B1(n_60),
.B2(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_49),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_0),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_60),
.B1(n_52),
.B2(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_58),
.B1(n_62),
.B2(n_61),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_55),
.B1(n_51),
.B2(n_66),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_98),
.B1(n_100),
.B2(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_57),
.B1(n_21),
.B2(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_15),
.B1(n_46),
.B2(n_44),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_112),
.B(n_110),
.C(n_106),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_14),
.B1(n_42),
.B2(n_41),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_112),
.B1(n_113),
.B2(n_47),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_12),
.B1(n_38),
.B2(n_36),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_3),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_120),
.B(n_124),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_115),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_127),
.Y(n_132)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_129),
.Y(n_133)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_131),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_95),
.C(n_116),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_135),
.B1(n_132),
.B2(n_29),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_127),
.A2(n_98),
.B1(n_96),
.B2(n_94),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_115),
.B1(n_114),
.B2(n_107),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_117),
.B(n_101),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_140),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_142),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_16),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_144),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_137),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_146),
.B(n_141),
.CI(n_143),
.CON(n_150),
.SN(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_148),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_150),
.C(n_149),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_10),
.B(n_35),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_34),
.Y(n_154)
);

NAND4xp25_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_32),
.C(n_31),
.D(n_27),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_4),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_5),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_117),
.C(n_7),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_6),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_9),
.C(n_7),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_6),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_8),
.Y(n_163)
);


endmodule