module fake_netlist_1_9099_n_578 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_578);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_578;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g74 ( .A(n_43), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_7), .Y(n_75) );
INVxp67_ASAP7_75t_SL g76 ( .A(n_41), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_57), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_67), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_51), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_48), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_7), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_59), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_68), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_53), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_39), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_14), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_69), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_46), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_61), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_24), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_31), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_52), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_3), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_36), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_12), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_20), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_23), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_70), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_16), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_29), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_4), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_38), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_6), .Y(n_103) );
INVxp33_ASAP7_75t_SL g104 ( .A(n_60), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_22), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_44), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_13), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_10), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_72), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_49), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_50), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_56), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_5), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_63), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_27), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_0), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_28), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_45), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_99), .B(n_0), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_75), .B(n_1), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_118), .Y(n_123) );
NOR2xp33_ASAP7_75t_R g124 ( .A(n_79), .B(n_83), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_75), .B(n_1), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_79), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_91), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_74), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_93), .B(n_2), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_93), .B(n_3), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_81), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_83), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_87), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_74), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_95), .B(n_4), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_96), .B(n_5), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_87), .Y(n_138) );
NAND2xp33_ASAP7_75t_L g139 ( .A(n_98), .B(n_34), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_101), .B(n_107), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_113), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_120), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_113), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_84), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_84), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_77), .B(n_6), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_118), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_98), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_85), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_103), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_102), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_85), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_108), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_89), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_102), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_109), .B(n_8), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_129), .B(n_156), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_124), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
NAND2x1p5_ASAP7_75t_L g167 ( .A(n_129), .B(n_119), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_129), .B(n_116), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_128), .A2(n_152), .B(n_135), .C(n_140), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_126), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_156), .B(n_119), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_128), .B(n_92), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_123), .Y(n_177) );
AOI22x1_ASAP7_75t_L g178 ( .A1(n_157), .A2(n_159), .B1(n_144), .B2(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_123), .B(n_115), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g181 ( .A1(n_131), .A2(n_86), .B1(n_114), .B2(n_117), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_130), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_132), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_133), .B(n_104), .Y(n_185) );
INVx4_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_130), .Y(n_187) );
INVx4_ASAP7_75t_L g188 ( .A(n_144), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_138), .B(n_106), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_150), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_149), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_140), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_142), .B(n_115), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_150), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_127), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_136), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_142), .B(n_89), .Y(n_200) );
AND2x6_ASAP7_75t_L g201 ( .A(n_136), .B(n_92), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_147), .B(n_97), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
INVxp33_ASAP7_75t_L g204 ( .A(n_141), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_147), .B(n_100), .Y(n_205) );
OAI22xp33_ASAP7_75t_L g206 ( .A1(n_122), .A2(n_117), .B1(n_105), .B2(n_111), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_150), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_155), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_152), .A2(n_112), .B1(n_110), .B2(n_94), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_155), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_155), .Y(n_212) );
NAND2x1p5_ASAP7_75t_L g213 ( .A(n_157), .B(n_80), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_155), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_155), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_158), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_151), .A2(n_105), .B1(n_90), .B2(n_76), .Y(n_217) );
AND2x4_ASAP7_75t_L g218 ( .A(n_141), .B(n_78), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_158), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_127), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_158), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_198), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_204), .B(n_154), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_186), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_163), .B(n_121), .Y(n_225) );
NOR2x1_ASAP7_75t_L g226 ( .A(n_206), .B(n_161), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_186), .Y(n_227) );
BUFx2_ASAP7_75t_L g228 ( .A(n_183), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_163), .B(n_161), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_198), .Y(n_230) );
NOR2xp33_ASAP7_75t_R g231 ( .A(n_172), .B(n_160), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_167), .A2(n_122), .B1(n_125), .B2(n_137), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_188), .Y(n_233) );
BUFx4f_ASAP7_75t_L g234 ( .A(n_201), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_188), .Y(n_235) );
NOR2x1_ASAP7_75t_L g236 ( .A(n_180), .B(n_137), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_218), .B(n_148), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_188), .Y(n_238) );
NOR3xp33_ASAP7_75t_SL g239 ( .A(n_184), .B(n_125), .C(n_148), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_192), .B(n_127), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_183), .B(n_159), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_173), .B(n_159), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_190), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_190), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_201), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_163), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_218), .B(n_139), .Y(n_247) );
NAND2xp33_ASAP7_75t_SL g248 ( .A(n_165), .B(n_158), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_173), .B(n_145), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_167), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_218), .B(n_145), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_173), .B(n_143), .Y(n_252) );
NOR3xp33_ASAP7_75t_SL g253 ( .A(n_181), .B(n_153), .C(n_11), .Y(n_253) );
OR2x6_ASAP7_75t_L g254 ( .A(n_177), .B(n_143), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_195), .B(n_134), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_179), .B(n_182), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_202), .B(n_134), .Y(n_257) );
INVxp67_ASAP7_75t_SL g258 ( .A(n_167), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_177), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_175), .Y(n_260) );
INVx2_ASAP7_75t_SL g261 ( .A(n_201), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_202), .B(n_158), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_175), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_175), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_164), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_200), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_213), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_187), .B(n_158), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_196), .B(n_37), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_193), .B(n_35), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_202), .B(n_9), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_162), .Y(n_272) );
AND2x6_ASAP7_75t_SL g273 ( .A(n_185), .B(n_12), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_193), .B(n_47), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_199), .B(n_15), .Y(n_275) );
OR2x6_ASAP7_75t_L g276 ( .A(n_169), .B(n_16), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_201), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_200), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_213), .B(n_54), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_213), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_164), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_260), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_227), .Y(n_284) );
NAND2xp33_ASAP7_75t_L g285 ( .A(n_250), .B(n_178), .Y(n_285) );
BUFx5_ASAP7_75t_L g286 ( .A(n_281), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_228), .B(n_217), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_229), .B(n_205), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_229), .B(n_205), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_258), .A2(n_189), .B1(n_205), .B2(n_169), .Y(n_290) );
AOI21x1_ASAP7_75t_L g291 ( .A1(n_280), .A2(n_203), .B(n_169), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_229), .A2(n_210), .B1(n_220), .B2(n_170), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_263), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_227), .Y(n_294) );
AND2x6_ASAP7_75t_L g295 ( .A(n_245), .B(n_221), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_264), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_266), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_241), .B(n_178), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_278), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_259), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_242), .B(n_221), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_227), .B(n_221), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_227), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
BUFx12f_ASAP7_75t_L g306 ( .A(n_276), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_240), .B(n_171), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_256), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_232), .B(n_171), .Y(n_309) );
OAI22xp33_ASAP7_75t_L g310 ( .A1(n_276), .A2(n_174), .B1(n_216), .B2(n_176), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_223), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_267), .A2(n_176), .B1(n_216), .B2(n_174), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_267), .A2(n_214), .B1(n_166), .B2(n_211), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_233), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_281), .Y(n_316) );
INVx6_ASAP7_75t_L g317 ( .A(n_256), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_225), .B(n_17), .Y(n_318) );
INVx4_ASAP7_75t_L g319 ( .A(n_234), .Y(n_319) );
NOR2xp33_ASAP7_75t_SL g320 ( .A(n_234), .B(n_166), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_233), .Y(n_321) );
AND2x2_ASAP7_75t_SL g322 ( .A(n_271), .B(n_219), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_233), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_233), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_244), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_249), .A2(n_211), .B(n_214), .C(n_215), .Y(n_326) );
INVx2_ASAP7_75t_SL g327 ( .A(n_254), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_261), .B(n_171), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_245), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_244), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_237), .B(n_18), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_311), .B(n_254), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_291), .A2(n_280), .B(n_270), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_283), .Y(n_334) );
AOI21xp33_ASAP7_75t_L g335 ( .A1(n_310), .A2(n_269), .B(n_226), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_318), .A2(n_256), .B1(n_275), .B2(n_249), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_321), .Y(n_338) );
AOI22xp33_ASAP7_75t_SL g339 ( .A1(n_306), .A2(n_231), .B1(n_225), .B2(n_247), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_318), .A2(n_253), .B1(n_239), .B2(n_225), .C(n_251), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_294), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_287), .A2(n_252), .B1(n_268), .B2(n_255), .C(n_257), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_296), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_286), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_294), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_300), .B(n_236), .Y(n_346) );
AO21x2_ASAP7_75t_L g347 ( .A1(n_326), .A2(n_274), .B(n_270), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_304), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
NAND2xp33_ASAP7_75t_SL g350 ( .A(n_327), .B(n_277), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_299), .Y(n_351) );
AOI221x1_ASAP7_75t_L g352 ( .A1(n_326), .A2(n_268), .B1(n_248), .B2(n_219), .C(n_168), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_306), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_288), .B(n_238), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_308), .A2(n_262), .B1(n_248), .B2(n_230), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_301), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_317), .A2(n_235), .B1(n_224), .B2(n_243), .Y(n_357) );
AO21x1_ASAP7_75t_L g358 ( .A1(n_285), .A2(n_274), .B(n_212), .Y(n_358) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_290), .A2(n_222), .B1(n_230), .B2(n_273), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_304), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_344), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_334), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_359), .A2(n_282), .B1(n_305), .B2(n_289), .C(n_292), .Y(n_363) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_332), .A2(n_313), .B1(n_331), .B2(n_317), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_334), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_337), .A2(n_316), .B1(n_322), .B2(n_309), .Y(n_366) );
AOI21x1_ASAP7_75t_L g367 ( .A1(n_358), .A2(n_298), .B(n_303), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_337), .A2(n_316), .B1(n_322), .B2(n_329), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_342), .A2(n_321), .B1(n_315), .B2(n_324), .Y(n_369) );
INVx5_ASAP7_75t_SL g370 ( .A(n_344), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_336), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_333), .A2(n_312), .B(n_314), .Y(n_372) );
OAI22xp5_ASAP7_75t_SL g373 ( .A1(n_339), .A2(n_265), .B1(n_319), .B2(n_284), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_342), .A2(n_302), .B1(n_307), .B2(n_285), .C(n_325), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_354), .B(n_286), .Y(n_375) );
AOI22xp5_ASAP7_75t_SL g376 ( .A1(n_353), .A2(n_295), .B1(n_319), .B2(n_284), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g377 ( .A1(n_340), .A2(n_325), .B1(n_319), .B2(n_323), .C(n_284), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_344), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_339), .A2(n_286), .B1(n_330), .B2(n_323), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_335), .A2(n_323), .B1(n_330), .B2(n_324), .C(n_315), .Y(n_380) );
OR2x6_ASAP7_75t_L g381 ( .A(n_332), .B(n_286), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_338), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_333), .A2(n_303), .B(n_328), .Y(n_383) );
OA21x2_ASAP7_75t_L g384 ( .A1(n_352), .A2(n_208), .B(n_209), .Y(n_384) );
AOI22xp33_ASAP7_75t_SL g385 ( .A1(n_353), .A2(n_286), .B1(n_295), .B2(n_320), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_363), .A2(n_346), .B1(n_343), .B2(n_336), .C(n_351), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_364), .A2(n_349), .B1(n_351), .B2(n_343), .C(n_356), .Y(n_387) );
AO21x2_ASAP7_75t_L g388 ( .A1(n_367), .A2(n_358), .B(n_335), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_375), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_375), .B(n_362), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_373), .A2(n_354), .B1(n_356), .B2(n_349), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_365), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_381), .A2(n_338), .B1(n_357), .B2(n_350), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_371), .B(n_338), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_382), .B(n_360), .Y(n_395) );
INVx2_ASAP7_75t_SL g396 ( .A(n_378), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_381), .B(n_338), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_366), .A2(n_355), .B1(n_360), .B2(n_348), .C(n_345), .Y(n_398) );
OAI31xp33_ASAP7_75t_L g399 ( .A1(n_368), .A2(n_355), .A3(n_360), .B(n_348), .Y(n_399) );
OA21x2_ASAP7_75t_L g400 ( .A1(n_372), .A2(n_352), .B(n_333), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_382), .Y(n_401) );
AOI21x1_ASAP7_75t_L g402 ( .A1(n_367), .A2(n_384), .B(n_372), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_383), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_381), .B(n_348), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_379), .A2(n_345), .B1(n_341), .B2(n_328), .C(n_330), .Y(n_405) );
AND2x4_ASAP7_75t_L g406 ( .A(n_381), .B(n_345), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_383), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_361), .Y(n_408) );
OR2x6_ASAP7_75t_L g409 ( .A(n_378), .B(n_341), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_374), .B(n_162), .C(n_168), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_377), .B(n_330), .Y(n_411) );
AO21x2_ASAP7_75t_L g412 ( .A1(n_369), .A2(n_347), .B(n_207), .Y(n_412) );
INVx4_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_380), .A2(n_347), .B1(n_295), .B2(n_162), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_376), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_384), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_413), .B(n_378), .Y(n_417) );
AOI33xp33_ASAP7_75t_L g418 ( .A1(n_391), .A2(n_385), .A3(n_215), .B1(n_209), .B2(n_208), .B3(n_207), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_389), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_392), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_392), .B(n_361), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_413), .B(n_378), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_395), .B(n_370), .Y(n_423) );
INVx4_ASAP7_75t_L g424 ( .A(n_406), .Y(n_424) );
INVx5_ASAP7_75t_L g425 ( .A(n_409), .Y(n_425) );
AND2x4_ASAP7_75t_SL g426 ( .A(n_406), .B(n_370), .Y(n_426) );
INVx5_ASAP7_75t_L g427 ( .A(n_409), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_395), .B(n_390), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_416), .Y(n_429) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_406), .B(n_370), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_403), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_416), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_401), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_390), .B(n_370), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_407), .Y(n_435) );
CKINVDCx16_ASAP7_75t_R g436 ( .A(n_413), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_386), .A2(n_197), .B(n_194), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_407), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_394), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_408), .Y(n_442) );
INVx4_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_394), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_402), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_412), .B(n_404), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_412), .B(n_347), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_400), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_415), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_400), .Y(n_451) );
OAI31xp33_ASAP7_75t_L g452 ( .A1(n_410), .A2(n_19), .A3(n_20), .B(n_21), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_397), .B(n_19), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_396), .Y(n_454) );
BUFx5_ASAP7_75t_L g455 ( .A(n_399), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_396), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_412), .B(n_71), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_388), .B(n_25), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_387), .B(n_295), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_453), .B(n_411), .C(n_405), .Y(n_461) );
NOR3xp33_ASAP7_75t_SL g462 ( .A(n_453), .B(n_398), .C(n_393), .Y(n_462) );
INVx4_ASAP7_75t_L g463 ( .A(n_426), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_424), .B(n_388), .Y(n_464) );
OR2x6_ASAP7_75t_L g465 ( .A(n_443), .B(n_414), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_450), .B(n_26), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_450), .B(n_30), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_420), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_436), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_419), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_426), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_428), .B(n_32), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_444), .B(n_219), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_446), .B(n_33), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_444), .B(n_219), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_446), .B(n_40), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_424), .B(n_42), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_440), .B(n_55), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_439), .B(n_219), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_433), .B(n_168), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_429), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_442), .B(n_58), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_434), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_421), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_448), .B(n_62), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_448), .B(n_64), .Y(n_486) );
NOR2xp33_ASAP7_75t_R g487 ( .A(n_436), .B(n_65), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_421), .B(n_66), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_434), .B(n_168), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_454), .Y(n_490) );
NAND4xp25_ASAP7_75t_L g491 ( .A(n_452), .B(n_191), .C(n_272), .D(n_73), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_431), .Y(n_492) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_443), .B(n_162), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_435), .B(n_438), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_435), .B(n_438), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_432), .B(n_451), .Y(n_496) );
NAND2x1_ASAP7_75t_L g497 ( .A(n_443), .B(n_457), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_458), .B(n_451), .Y(n_498) );
NAND2xp33_ASAP7_75t_R g499 ( .A(n_417), .B(n_422), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_449), .B(n_458), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_496), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_469), .B(n_441), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_470), .B(n_455), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_468), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_490), .B(n_423), .Y(n_505) );
INVx2_ASAP7_75t_SL g506 ( .A(n_471), .Y(n_506) );
INVxp33_ASAP7_75t_L g507 ( .A(n_487), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_463), .A2(n_460), .B1(n_425), .B2(n_427), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g509 ( .A1(n_463), .A2(n_460), .B1(n_425), .B2(n_427), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_498), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_494), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_494), .Y(n_512) );
AOI21xp33_ASAP7_75t_L g513 ( .A1(n_466), .A2(n_459), .B(n_457), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_496), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g515 ( .A1(n_462), .A2(n_456), .B1(n_458), .B2(n_441), .C(n_449), .Y(n_515) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_467), .A2(n_457), .B(n_456), .Y(n_516) );
AOI322xp5_ASAP7_75t_L g517 ( .A1(n_472), .A2(n_430), .A3(n_449), .B1(n_458), .B2(n_447), .C1(n_445), .C2(n_425), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_483), .B(n_484), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_495), .Y(n_519) );
O2A1O1Ixp5_ASAP7_75t_L g520 ( .A1(n_463), .A2(n_417), .B(n_422), .C(n_447), .Y(n_520) );
AND2x2_ASAP7_75t_SL g521 ( .A(n_477), .B(n_430), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_492), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_474), .B(n_455), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_491), .B(n_418), .C(n_437), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_499), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_461), .A2(n_455), .B1(n_417), .B2(n_427), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_497), .A2(n_425), .B(n_427), .Y(n_527) );
OAI21xp33_ASAP7_75t_SL g528 ( .A1(n_493), .A2(n_425), .B(n_427), .Y(n_528) );
AOI221x1_ASAP7_75t_SL g529 ( .A1(n_464), .A2(n_455), .B1(n_477), .B2(n_473), .C(n_475), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_511), .B(n_476), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_512), .B(n_485), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_525), .B(n_465), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_519), .B(n_486), .Y(n_533) );
AND2x4_ASAP7_75t_SL g534 ( .A(n_502), .B(n_488), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_525), .B(n_465), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_507), .B(n_480), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_518), .B(n_500), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_506), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_510), .B(n_500), .Y(n_539) );
HAxp5_ASAP7_75t_SL g540 ( .A(n_526), .B(n_465), .CON(n_540), .SN(n_540) );
OAI211xp5_ASAP7_75t_L g541 ( .A1(n_528), .A2(n_488), .B(n_489), .C(n_479), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_520), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_521), .B(n_478), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_515), .B(n_505), .Y(n_544) );
NAND2xp33_ASAP7_75t_R g545 ( .A(n_527), .B(n_482), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_520), .B(n_481), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_501), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_514), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_503), .B(n_455), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_504), .B(n_455), .Y(n_550) );
INVxp67_ASAP7_75t_SL g551 ( .A(n_546), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_544), .B(n_522), .Y(n_552) );
XNOR2xp5_ASAP7_75t_L g553 ( .A(n_543), .B(n_529), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_541), .A2(n_524), .B(n_517), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_536), .A2(n_513), .B1(n_523), .B2(n_516), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_539), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_538), .B(n_509), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_548), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_542), .B(n_508), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_536), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_537), .Y(n_561) );
NOR2xp33_ASAP7_75t_R g562 ( .A(n_553), .B(n_545), .Y(n_562) );
AO22x2_ASAP7_75t_L g563 ( .A1(n_551), .A2(n_535), .B1(n_532), .B2(n_546), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_553), .A2(n_534), .B1(n_547), .B2(n_530), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_560), .Y(n_565) );
AOI321xp33_ASAP7_75t_L g566 ( .A1(n_559), .A2(n_540), .A3(n_549), .B1(n_533), .B2(n_531), .C(n_550), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_557), .B(n_534), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_552), .A2(n_561), .B1(n_555), .B2(n_556), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_558), .A2(n_554), .B(n_553), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_565), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_567), .B(n_563), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_563), .B(n_562), .Y(n_572) );
OAI22x1_ASAP7_75t_L g573 ( .A1(n_572), .A2(n_569), .B1(n_568), .B2(n_566), .Y(n_573) );
XNOR2xp5_ASAP7_75t_L g574 ( .A(n_570), .B(n_564), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_574), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_575), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_576), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_577), .A2(n_573), .B(n_571), .Y(n_578) );
endmodule