module fake_jpeg_12827_n_262 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_35),
.B1(n_28),
.B2(n_21),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_54),
.B1(n_64),
.B2(n_70),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_18),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_18),
.B1(n_22),
.B2(n_28),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_22),
.B1(n_32),
.B2(n_30),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_55),
.A2(n_65),
.B1(n_75),
.B2(n_26),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_22),
.B1(n_33),
.B2(n_29),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_19),
.B1(n_17),
.B2(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_22),
.B1(n_32),
.B2(n_30),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_26),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_33),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_73),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_34),
.B1(n_27),
.B2(n_20),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_37),
.A2(n_34),
.B1(n_20),
.B2(n_27),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_64),
.B1(n_54),
.B2(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_29),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_19),
.B1(n_17),
.B2(n_26),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_77),
.A2(n_81),
.B(n_91),
.Y(n_126)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_97),
.Y(n_117)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_14),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_13),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_44),
.B1(n_26),
.B2(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_100),
.B1(n_62),
.B2(n_51),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_14),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_12),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_63),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_96),
.Y(n_133)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_103),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_50),
.B(n_13),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_104),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_44),
.B1(n_38),
.B2(n_36),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_68),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_31),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_67),
.C(n_49),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_107),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_66),
.B(n_63),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_105),
.B(n_77),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_68),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_127),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_103),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_84),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_131),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_63),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_120),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_62),
.B1(n_24),
.B2(n_31),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_88),
.B(n_95),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_62),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_24),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_12),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_144),
.C(n_132),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_109),
.B(n_114),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_137),
.B(n_140),
.Y(n_182)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_86),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_113),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_147),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_105),
.C(n_90),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_153),
.B1(n_118),
.B2(n_116),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_96),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_154),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_80),
.B1(n_83),
.B2(n_82),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_132),
.B1(n_125),
.B2(n_112),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_120),
.B(n_78),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_100),
.B1(n_38),
.B2(n_24),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_158),
.B1(n_1),
.B2(n_3),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_108),
.B(n_0),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_170),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_184),
.B1(n_141),
.B2(n_158),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_167),
.C(n_173),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_127),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_171),
.A2(n_153),
.B(n_150),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_144),
.C(n_157),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_175),
.B(n_180),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_6),
.C(n_7),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_145),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_125),
.B1(n_119),
.B2(n_128),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_156),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_118),
.B(n_128),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_146),
.B(n_139),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_136),
.A2(n_112),
.B1(n_118),
.B2(n_38),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_185),
.A2(n_152),
.B1(n_141),
.B2(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_189),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_190),
.A2(n_161),
.B1(n_10),
.B2(n_11),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_194),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_199),
.B1(n_202),
.B2(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_135),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g198 ( 
.A1(n_169),
.A2(n_3),
.B(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_199)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_6),
.Y(n_201)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_179),
.C(n_167),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_178),
.B(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_7),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_205),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_187),
.B(n_173),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_193),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_194),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_202),
.A2(n_185),
.B1(n_171),
.B2(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_220),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_176),
.C(n_179),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_203),
.C(n_186),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_190),
.A2(n_177),
.B1(n_184),
.B2(n_183),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_228),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_211),
.B(n_191),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_211),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_192),
.C(n_197),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_212),
.C(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

AOI221xp5_ASAP7_75t_L g228 ( 
.A1(n_207),
.A2(n_195),
.B1(n_188),
.B2(n_201),
.C(n_200),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_232),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_235),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_222),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_219),
.C(n_215),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_237),
.C(n_225),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_208),
.B1(n_218),
.B2(n_209),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_241),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_246),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_224),
.B1(n_218),
.B2(n_217),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_244),
.A2(n_242),
.B1(n_199),
.B2(n_215),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_239),
.A2(n_231),
.B(n_226),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_240),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_249),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_248),
.A2(n_213),
.B1(n_238),
.B2(n_205),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_252),
.C(n_253),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_240),
.B1(n_198),
.B2(n_161),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_250),
.A2(n_245),
.B(n_246),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_243),
.B(n_250),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_257),
.A2(n_258),
.B(n_254),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_256),
.B(n_252),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_198),
.B(n_10),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_9),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_261),
.B(n_11),
.Y(n_262)
);


endmodule