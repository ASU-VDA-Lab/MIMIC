module fake_jpeg_13302_n_426 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_426);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_44),
.B(n_60),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_67),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_47),
.Y(n_132)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_20),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_53),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_16),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_62),
.B(n_81),
.Y(n_99)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_14),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_68),
.Y(n_111)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_77),
.B(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_22),
.B(n_14),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_39),
.B(n_13),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_83),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_22),
.B(n_13),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_9),
.Y(n_124)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_18),
.C(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_32),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_51),
.A2(n_26),
.B1(n_37),
.B2(n_36),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_93),
.A2(n_104),
.B1(n_107),
.B2(n_117),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_40),
.Y(n_96)
);

OR2x2_ASAP7_75t_SL g175 ( 
.A(n_96),
.B(n_31),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_37),
.B1(n_36),
.B2(n_43),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_100),
.A2(n_130),
.B1(n_24),
.B2(n_31),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_46),
.A2(n_43),
.B1(n_42),
.B2(n_28),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_47),
.A2(n_37),
.B1(n_27),
.B2(n_19),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_115),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_63),
.A2(n_37),
.B1(n_27),
.B2(n_19),
.Y(n_117)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_139),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_75),
.A2(n_19),
.B1(n_27),
.B2(n_38),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_141),
.B1(n_32),
.B2(n_70),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_42),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_1),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_54),
.A2(n_28),
.B1(n_34),
.B2(n_18),
.Y(n_130)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_55),
.Y(n_137)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_49),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_56),
.A2(n_40),
.B1(n_34),
.B2(n_16),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_48),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_143),
.B(n_145),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_87),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_146),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_115),
.A2(n_109),
.B(n_116),
.C(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_147),
.B(n_152),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_148),
.B(n_180),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_89),
.B(n_88),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_151),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_92),
.B(n_0),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_0),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_153),
.B(n_174),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_106),
.A2(n_85),
.B1(n_72),
.B2(n_76),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_154),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_108),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_155),
.B(n_170),
.Y(n_197)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_158),
.A2(n_163),
.B1(n_172),
.B2(n_192),
.Y(n_198)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_107),
.A2(n_79),
.B1(n_74),
.B2(n_73),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_93),
.A2(n_71),
.B1(n_64),
.B2(n_58),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_64),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_169),
.C(n_171),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVx4_ASAP7_75t_SL g202 ( 
.A(n_166),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_94),
.A2(n_31),
.B1(n_24),
.B2(n_49),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_167),
.A2(n_193),
.B1(n_157),
.B2(n_184),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_103),
.B(n_118),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_99),
.B(n_13),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_103),
.B(n_0),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_175),
.B(n_181),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_176),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_111),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_177),
.B(n_178),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_131),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_2),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_2),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_95),
.B(n_9),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_183),
.B(n_186),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_187),
.B1(n_123),
.B2(n_138),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_102),
.B(n_12),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_102),
.A2(n_31),
.B1(n_4),
.B2(n_5),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_94),
.B(n_10),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_188),
.B(n_166),
.Y(n_235)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_191),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_117),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_151),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_235),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_149),
.A2(n_97),
.B1(n_113),
.B2(n_120),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_201),
.A2(n_203),
.B1(n_208),
.B2(n_213),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_97),
.B1(n_113),
.B2(n_120),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_204),
.A2(n_230),
.B1(n_234),
.B2(n_231),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_143),
.B1(n_145),
.B2(n_162),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_205),
.A2(n_229),
.B1(n_234),
.B2(n_169),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_162),
.A2(n_132),
.B1(n_138),
.B2(n_135),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_162),
.A2(n_119),
.B1(n_6),
.B2(n_8),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_152),
.A2(n_3),
.B1(n_153),
.B2(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_214),
.A2(n_221),
.B1(n_225),
.B2(n_236),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_171),
.B1(n_181),
.B2(n_151),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_171),
.B1(n_181),
.B2(n_164),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_144),
.A2(n_150),
.B1(n_146),
.B2(n_160),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_159),
.A2(n_147),
.B1(n_193),
.B2(n_179),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_164),
.A2(n_169),
.B1(n_190),
.B2(n_168),
.Y(n_236)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_173),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_242),
.B(n_246),
.Y(n_293)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_245),
.A2(n_254),
.B1(n_257),
.B2(n_275),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_156),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_226),
.A2(n_189),
.B1(n_165),
.B2(n_161),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_247),
.A2(n_265),
.B1(n_244),
.B2(n_261),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_220),
.A2(n_166),
.B(n_215),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_249),
.A2(n_252),
.B(n_267),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_217),
.B(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_251),
.B(n_256),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_215),
.A2(n_231),
.B(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_205),
.A2(n_230),
.B1(n_215),
.B2(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_214),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_198),
.A2(n_201),
.B1(n_208),
.B2(n_203),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_258),
.A2(n_272),
.B1(n_248),
.B2(n_253),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_259),
.B(n_260),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_221),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_195),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_266),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_219),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_264),
.Y(n_297)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_211),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_219),
.C(n_204),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_267),
.C(n_263),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_232),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_269),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_200),
.B(n_232),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_273),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_200),
.B(n_233),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_271),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_198),
.A2(n_213),
.B1(n_226),
.B2(n_206),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_195),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_206),
.A2(n_216),
.B1(n_222),
.B2(n_223),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_254),
.B(n_223),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_292),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_202),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_290),
.C(n_292),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_243),
.A2(n_222),
.B(n_210),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_283),
.A2(n_294),
.B(n_300),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_255),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_249),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_243),
.A2(n_259),
.B(n_245),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_308),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_256),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_277),
.C(n_289),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_272),
.A2(n_238),
.B(n_260),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_241),
.A2(n_239),
.B(n_240),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_302),
.A2(n_300),
.B(n_304),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_262),
.A2(n_248),
.B(n_275),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_303),
.A2(n_294),
.B(n_283),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_250),
.B1(n_265),
.B2(n_303),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_250),
.B(n_273),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_310),
.A2(n_328),
.B(n_320),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_258),
.C(n_266),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_327),
.C(n_329),
.Y(n_341)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_317),
.A2(n_334),
.B1(n_315),
.B2(n_332),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_324),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_285),
.Y(n_319)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_276),
.Y(n_320)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_321),
.A2(n_299),
.B(n_309),
.Y(n_349)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

XOR2x2_ASAP7_75t_SL g324 ( 
.A(n_282),
.B(n_307),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_276),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_330),
.Y(n_356)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_289),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_297),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_301),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_331),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_280),
.B(n_286),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_333),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_306),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_287),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_288),
.A2(n_286),
.B1(n_287),
.B2(n_291),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_335),
.A2(n_299),
.B1(n_322),
.B2(n_323),
.Y(n_348)
);

XNOR2x1_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_313),
.Y(n_368)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_284),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_353),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_331),
.A2(n_284),
.B1(n_291),
.B2(n_288),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_346),
.A2(n_348),
.B1(n_350),
.B2(n_317),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_349),
.A2(n_355),
.B1(n_312),
.B2(n_329),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_321),
.A2(n_315),
.B1(n_309),
.B2(n_325),
.Y(n_350)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_326),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_356),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_313),
.B(n_327),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_347),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g359 ( 
.A1(n_355),
.A2(n_324),
.B(n_319),
.Y(n_359)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_359),
.Y(n_378)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_316),
.Y(n_361)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_361),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_362),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_347),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_368),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_367),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_350),
.A2(n_314),
.B1(n_312),
.B2(n_318),
.Y(n_365)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_336),
.A2(n_342),
.B1(n_345),
.B2(n_337),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_345),
.A2(n_335),
.B1(n_333),
.B2(n_311),
.Y(n_369)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_369),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_377),
.C(n_363),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_371),
.B(n_372),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_346),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_339),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_373),
.B(n_374),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_343),
.A2(n_349),
.B1(n_351),
.B2(n_354),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_341),
.A2(n_342),
.B1(n_350),
.B2(n_331),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_375),
.A2(n_376),
.B(n_365),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_357),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_358),
.C(n_313),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_375),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_377),
.B(n_370),
.C(n_368),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_385),
.Y(n_398)
);

FAx1_ASAP7_75t_SL g385 ( 
.A(n_359),
.B(n_373),
.CI(n_361),
.CON(n_385),
.SN(n_385)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_384),
.C(n_388),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_381),
.B(n_364),
.C(n_360),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_397),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_383),
.A2(n_366),
.B1(n_372),
.B2(n_371),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_395),
.A2(n_378),
.B1(n_390),
.B2(n_383),
.Y(n_409)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_379),
.Y(n_396)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_396),
.Y(n_402)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_391),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_385),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_399),
.B(n_400),
.Y(n_408)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_389),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_376),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_385),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_388),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_404),
.B(n_406),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_405),
.B(n_393),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_380),
.C(n_390),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_407),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_409),
.B(n_401),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_410),
.B(n_415),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_413),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_395),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_392),
.C(n_382),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_414),
.B(n_408),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_419),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_411),
.B(n_414),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_418),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_420),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_422),
.A2(n_421),
.B(n_416),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_419),
.C(n_408),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_402),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_392),
.Y(n_426)
);


endmodule