module real_jpeg_2559_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_3),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_3),
.B(n_24),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_3),
.A2(n_87),
.B(n_90),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_3),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_3),
.B(n_54),
.C(n_64),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_34),
.B1(n_36),
.B2(n_92),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_3),
.B(n_51),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_103),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_3),
.A2(n_24),
.B(n_76),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_4),
.A2(n_34),
.B1(n_36),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_72),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_5),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_6),
.A2(n_34),
.B1(n_36),
.B2(n_40),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_6),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_147)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_11),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_11),
.A2(n_34),
.B1(n_36),
.B2(n_59),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_13),
.A2(n_34),
.B1(n_36),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_69),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_14),
.A2(n_26),
.B1(n_87),
.B2(n_88),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_14),
.A2(n_26),
.B1(n_34),
.B2(n_36),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_14),
.A2(n_26),
.B1(n_53),
.B2(n_54),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_118),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_116),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_82),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_82),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_61),
.C(n_73),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_20),
.B(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_41),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_21),
.B(n_43),
.C(n_48),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_37),
.B2(n_38),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_23),
.A2(n_28),
.B1(n_33),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_24),
.A2(n_25),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g74 ( 
.A1(n_24),
.A2(n_30),
.A3(n_34),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_24),
.B(n_46),
.C(n_88),
.Y(n_115)
);

CKINVDCx6p67_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_25),
.A2(n_47),
.B(n_91),
.C(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_28),
.A2(n_33),
.B1(n_39),
.B2(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

OA22x2_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_33),
.B(n_92),
.Y(n_127)
);

CKINVDCx6p67_ASAP7_75t_R g36 ( 
.A(n_34),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_36),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_34),
.B(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_48),
.B2(n_49),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_86),
.B1(n_93),
.B2(n_95),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_94),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_46),
.A2(n_47),
.B1(n_87),
.B2(n_88),
.Y(n_94)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B(n_57),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_50),
.B(n_80),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_50),
.A2(n_79),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_58),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_51),
.A2(n_60),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_51),
.A2(n_60),
.B1(n_92),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_51),
.A2(n_60),
.B1(n_144),
.B2(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_54),
.B(n_142),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_60),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_61),
.B(n_73),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_67),
.B(n_70),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_62),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_62),
.A2(n_103),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_62),
.A2(n_103),
.B1(n_129),
.B2(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_66),
.A2(n_68),
.B1(n_100),
.B2(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_74),
.B(n_78),
.Y(n_161)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B(n_81),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_104),
.B2(n_105),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_96),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_114),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_168),
.B(n_172),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_157),
.B(n_167),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_138),
.B(n_156),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_131),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_131),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_128),
.C(n_159),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_150),
.B(n_155),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_145),
.B(n_149),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_148),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_154),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_160),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_163),
.C(n_165),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_171),
.Y(n_172)
);


endmodule