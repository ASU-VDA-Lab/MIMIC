module fake_jpeg_8718_n_285 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_285);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_218;
wire n_63;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_19),
.B(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_27),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx9p33_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_24),
.B1(n_14),
.B2(n_15),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_14),
.B1(n_23),
.B2(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_15),
.B1(n_14),
.B2(n_37),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_68),
.B(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_64),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_26),
.B1(n_27),
.B2(n_51),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_37),
.B1(n_17),
.B2(n_23),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_44),
.B(n_49),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_45),
.A2(n_37),
.B1(n_36),
.B2(n_24),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_39),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_52),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_83),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_99),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_87),
.Y(n_109)
);

AOI22x1_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_36),
.B1(n_52),
.B2(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_86),
.B(n_89),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_77),
.B1(n_26),
.B2(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_56),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_0),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_30),
.C(n_34),
.Y(n_112)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_97),
.Y(n_115)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_96),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_107),
.B1(n_119),
.B2(n_90),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_82),
.A2(n_75),
.B1(n_65),
.B2(n_47),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_97),
.B1(n_87),
.B2(n_95),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_108),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_55),
.B1(n_48),
.B2(n_30),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_106),
.A2(n_110),
.B1(n_117),
.B2(n_118),
.Y(n_137)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_80),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_48),
.B1(n_55),
.B2(n_36),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_90),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_88),
.CI(n_20),
.CON(n_138),
.SN(n_138)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_34),
.C(n_73),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_121),
.C(n_80),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_48),
.B1(n_55),
.B2(n_76),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_64),
.B1(n_59),
.B2(n_67),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_29),
.C(n_28),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_56),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_78),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_140),
.Y(n_153)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_81),
.B(n_86),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_127),
.A2(n_132),
.B(n_138),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx5_ASAP7_75t_SL g162 ( 
.A(n_129),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_85),
.B1(n_93),
.B2(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_133),
.B(n_120),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_99),
.C(n_98),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_112),
.C(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_22),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_67),
.A3(n_29),
.B1(n_38),
.B2(n_20),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_144),
.B(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_22),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_114),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_20),
.B(n_18),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_16),
.B(n_18),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_107),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_111),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_151),
.C(n_165),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_119),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_157),
.Y(n_184)
);

OAI22x1_ASAP7_75t_SL g156 ( 
.A1(n_137),
.A2(n_120),
.B1(n_102),
.B2(n_105),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_13),
.B(n_22),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_167),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_164),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_102),
.B1(n_114),
.B2(n_119),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_163),
.A2(n_74),
.B1(n_77),
.B2(n_53),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_13),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_129),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_129),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_146),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_70),
.B(n_96),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_170),
.A2(n_145),
.B(n_125),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_123),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_182),
.C(n_191),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_183),
.B(n_165),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_168),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_177),
.B(n_190),
.Y(n_198)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_136),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_132),
.Y(n_181)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_135),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_170),
.A2(n_142),
.B(n_138),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_29),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_193),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_152),
.B1(n_159),
.B2(n_169),
.Y(n_201)
);

INVxp33_ASAP7_75t_SL g189 ( 
.A(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_70),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_39),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_192),
.B(n_157),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_167),
.B1(n_162),
.B2(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_163),
.C(n_153),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_175),
.A2(n_152),
.B1(n_158),
.B2(n_171),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_13),
.Y(n_229)
);

NOR2xp67_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_171),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_173),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_153),
.B1(n_162),
.B2(n_166),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_184),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_205),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_218),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_174),
.C(n_193),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_221),
.C(n_224),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_16),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_187),
.C(n_182),
.Y(n_221)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_176),
.C(n_179),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_191),
.C(n_183),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_230),
.C(n_16),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_162),
.B(n_11),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_0),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_63),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_38),
.C(n_53),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_207),
.A3(n_209),
.B1(n_206),
.B2(n_198),
.C1(n_211),
.C2(n_195),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_7),
.Y(n_253)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_11),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_195),
.B1(n_196),
.B2(n_201),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_236),
.B1(n_223),
.B2(n_226),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_242),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_240),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_224),
.B(n_18),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_244),
.C(n_1),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_227),
.A2(n_63),
.B(n_9),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_63),
.C(n_22),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_219),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_251),
.C(n_240),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_225),
.B(n_230),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_237),
.B(n_236),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_250),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_13),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_11),
.B1(n_10),
.B2(n_7),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_252),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_253),
.B(n_254),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_7),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_2),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_1),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_258),
.Y(n_267)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_3),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_239),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_265),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_263),
.A2(n_247),
.B(n_249),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_270),
.B(n_4),
.Y(n_275)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_237),
.B(n_249),
.C(n_251),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_266),
.C(n_259),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_273),
.C(n_4),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_261),
.B(n_264),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_272),
.B(n_3),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_276),
.B(n_277),
.C(n_267),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_4),
.C(n_5),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_278),
.B(n_5),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

OAI221xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_5),
.B1(n_6),
.B2(n_71),
.C(n_279),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_71),
.Y(n_285)
);


endmodule