module fake_jpeg_25525_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_3),
.B(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_14),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_20),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_5),
.Y(n_21)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_5),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_11),
.B1(n_16),
.B2(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_10),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_17),
.A2(n_16),
.B1(n_15),
.B2(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_16),
.B1(n_19),
.B2(n_9),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_33),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_34),
.B(n_24),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_23),
.B1(n_24),
.B2(n_10),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_24),
.A2(n_12),
.B1(n_10),
.B2(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_21),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_26),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_23),
.C(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_33),
.B1(n_30),
.B2(n_28),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_38),
.B(n_42),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_36),
.B1(n_20),
.B2(n_6),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_40),
.B(n_39),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_47),
.B(n_49),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_20),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_34),
.B(n_24),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_42),
.B(n_41),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_52),
.B(n_51),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_36),
.B(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_53),
.B(n_7),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_61),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_4),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_20),
.C(n_4),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_7),
.C(n_8),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_65),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_7),
.B(n_8),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

OAI21x1_ASAP7_75t_SL g67 ( 
.A1(n_66),
.A2(n_57),
.B(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_8),
.Y(n_71)
);

OA21x2_ASAP7_75t_SL g70 ( 
.A1(n_68),
.A2(n_69),
.B(n_65),
.Y(n_70)
);

AOI311xp33_ASAP7_75t_SL g73 ( 
.A1(n_70),
.A2(n_71),
.A3(n_0),
.B(n_1),
.C(n_2),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

OAI21x1_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B(n_0),
.Y(n_74)
);

BUFx24_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);


endmodule