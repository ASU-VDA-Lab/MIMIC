module fake_jpeg_7975_n_23 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_3),
.Y(n_7)
);

INVx13_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

NAND2x1_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_6),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_4),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_20)
);

A2O1A1O1Ixp25_ASAP7_75t_L g16 ( 
.A1(n_10),
.A2(n_1),
.B(n_11),
.C(n_12),
.D(n_7),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_18),
.C(n_9),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_14),
.B1(n_9),
.B2(n_8),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_13),
.B(n_8),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_19),
.A2(n_20),
.B(n_18),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_13),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_16),
.C(n_13),
.Y(n_23)
);


endmodule