module fake_jpeg_15294_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_0),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_1),
.Y(n_73)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_38),
.C(n_40),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_1),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_74),
.B(n_70),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_51),
.B1(n_49),
.B2(n_53),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_67),
.B1(n_71),
.B2(n_75),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_51),
.B1(n_39),
.B2(n_52),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_58),
.B1(n_38),
.B2(n_41),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_2),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_50),
.B1(n_48),
.B2(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_87),
.B1(n_3),
.B2(n_5),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_88),
.Y(n_89)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

OAI22x1_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_44),
.B1(n_47),
.B2(n_4),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_92),
.B1(n_84),
.B2(n_7),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_97),
.B1(n_94),
.B2(n_11),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_6),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_102),
.A2(n_9),
.B(n_10),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_22),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_6),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_107),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_113),
.B(n_94),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_111),
.A2(n_103),
.B1(n_109),
.B2(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_110),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_116),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_113),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_115),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_118),
.C(n_14),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_13),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_17),
.B(n_18),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_20),
.C(n_21),
.Y(n_124)
);

AOI321xp33_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_25),
.A3(n_26),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_33),
.Y(n_126)
);


endmodule