module fake_jpeg_13469_n_575 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_575);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_575;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_3),
.B(n_17),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_56),
.B(n_70),
.Y(n_117)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_57),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_18),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_71),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_60),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_67),
.Y(n_170)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_68),
.Y(n_127)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_31),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_31),
.B(n_17),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_24),
.B1(n_21),
.B2(n_32),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_79),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_32),
.Y(n_146)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

BUFx24_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx2_ASAP7_75t_R g168 ( 
.A(n_105),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_112),
.A2(n_155),
.B1(n_27),
.B2(n_35),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_70),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_118),
.B(n_125),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_56),
.B(n_46),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_123),
.B(n_138),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_59),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_25),
.B1(n_45),
.B2(n_41),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_129),
.A2(n_150),
.B1(n_34),
.B2(n_35),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_85),
.B(n_24),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_105),
.A2(n_54),
.B(n_45),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_139),
.B(n_22),
.C(n_54),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_146),
.B(n_1),
.C(n_2),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_79),
.B(n_21),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_149),
.B(n_158),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_57),
.A2(n_35),
.B1(n_45),
.B2(n_34),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_100),
.B(n_46),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_152),
.B(n_172),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_55),
.A2(n_41),
.B1(n_38),
.B2(n_28),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_72),
.B(n_36),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_65),
.B(n_36),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_20),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_74),
.B(n_50),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_119),
.Y(n_175)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_131),
.B(n_23),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_176),
.A2(n_194),
.B(n_157),
.Y(n_251)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_168),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_178),
.B(n_212),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_179),
.A2(n_136),
.B1(n_4),
.B2(n_5),
.Y(n_280)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_180),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_150),
.B1(n_76),
.B2(n_104),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_181),
.A2(n_185),
.B1(n_190),
.B2(n_174),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_126),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_182),
.B(n_183),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_29),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_117),
.A2(n_41),
.B1(n_38),
.B2(n_99),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_108),
.B1(n_106),
.B2(n_97),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_187),
.A2(n_200),
.B1(n_220),
.B2(n_235),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_133),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_188),
.B(n_195),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_173),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_189),
.B(n_196),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_130),
.A2(n_84),
.B1(n_94),
.B2(n_92),
.Y(n_190)
);

INVx13_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_191),
.Y(n_254)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_135),
.A2(n_34),
.B1(n_28),
.B2(n_50),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_114),
.B(n_42),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_127),
.B(n_42),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_197),
.B(n_205),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_134),
.B(n_29),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_198),
.B(n_218),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_201),
.Y(n_272)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_202),
.Y(n_293)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_204),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_168),
.B(n_14),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_127),
.B(n_27),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_206),
.B(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_141),
.Y(n_211)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_211),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_22),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_213),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_236),
.Y(n_242)
);

CKINVDCx12_ASAP7_75t_R g215 ( 
.A(n_113),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_215),
.Y(n_285)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_116),
.Y(n_217)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_217),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_159),
.B(n_0),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_219),
.B(n_228),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_132),
.A2(n_77),
.B1(n_90),
.B2(n_82),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_124),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_222),
.B(n_225),
.Y(n_238)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_223),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_170),
.B(n_51),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_144),
.B(n_51),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_110),
.B(n_1),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_229),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_110),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_132),
.B(n_2),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_116),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_230),
.B(n_231),
.Y(n_289)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_120),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_137),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_232),
.B(n_234),
.Y(n_247)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_120),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_128),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_171),
.A2(n_51),
.B1(n_80),
.B2(n_22),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_51),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_200),
.A2(n_111),
.B1(n_154),
.B2(n_143),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_249),
.A2(n_262),
.B1(n_268),
.B2(n_270),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_196),
.B(n_141),
.C(n_135),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_250),
.B(n_9),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_251),
.B(n_213),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_253),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_258),
.A2(n_267),
.B1(n_273),
.B2(n_280),
.Y(n_297)
);

AOI32xp33_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_102),
.A3(n_137),
.B1(n_66),
.B2(n_161),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g333 ( 
.A1(n_259),
.A2(n_11),
.B(n_12),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_183),
.A2(n_111),
.B1(n_143),
.B2(n_154),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_181),
.A2(n_174),
.B1(n_160),
.B2(n_151),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_189),
.A2(n_160),
.B1(n_151),
.B2(n_121),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_198),
.A2(n_121),
.B1(n_156),
.B2(n_22),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_190),
.A2(n_156),
.B1(n_54),
.B2(n_22),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_218),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_279),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_229),
.B(n_2),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_194),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_282),
.A2(n_288),
.B1(n_239),
.B2(n_238),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_186),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_212),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_221),
.B1(n_216),
.B2(n_233),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_212),
.B(n_12),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_288),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_175),
.B(n_207),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_204),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_184),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_295),
.B(n_304),
.Y(n_349)
);

INVx6_ASAP7_75t_SL g296 ( 
.A(n_264),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_296),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_264),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_299),
.Y(n_363)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_241),
.Y(n_300)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_300),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_247),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_301),
.B(n_329),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_302),
.A2(n_308),
.B1(n_246),
.B2(n_284),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_240),
.B(n_226),
.Y(n_304)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_254),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_177),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_306),
.B(n_313),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_258),
.A2(n_223),
.B1(n_231),
.B2(n_176),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_251),
.A2(n_209),
.B(n_211),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g354 ( 
.A1(n_309),
.A2(n_328),
.B(n_334),
.C(n_250),
.Y(n_354)
);

INVx13_ASAP7_75t_L g310 ( 
.A(n_285),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_310),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_325),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_245),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_242),
.B(n_261),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_316),
.C(n_320),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_282),
.A2(n_180),
.B1(n_202),
.B2(n_199),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_315),
.A2(n_319),
.B1(n_323),
.B2(n_343),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_242),
.B(n_203),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_291),
.Y(n_318)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_242),
.B(n_192),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_321),
.A2(n_333),
.B(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_266),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_322),
.B(n_324),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_270),
.A2(n_217),
.B1(n_213),
.B2(n_230),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_248),
.B(n_201),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_327),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_261),
.B(n_9),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_239),
.A2(n_191),
.B(n_11),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_243),
.B(n_210),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_328),
.Y(n_347)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_252),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_331),
.B(n_332),
.Y(n_374)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_239),
.A2(n_253),
.B(n_280),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_335),
.A2(n_286),
.B1(n_256),
.B2(n_244),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_265),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_338),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_289),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_245),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_341),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_269),
.B(n_275),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_340),
.B(n_342),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_248),
.B(n_269),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_279),
.B(n_281),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_293),
.A2(n_277),
.B1(n_256),
.B2(n_276),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_347),
.B(n_350),
.C(n_345),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_377),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_320),
.C(n_316),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_354),
.A2(n_372),
.B(n_361),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_355),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_296),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_358),
.B(n_364),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_297),
.A2(n_253),
.B1(n_267),
.B2(n_288),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_361),
.A2(n_380),
.B1(n_383),
.B2(n_348),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_310),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_367),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_321),
.Y(n_364)
);

NOR2x1_ASAP7_75t_L g365 ( 
.A(n_321),
.B(n_312),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_365),
.B(n_330),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_366),
.A2(n_368),
.B1(n_375),
.B2(n_379),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_310),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_336),
.A2(n_271),
.B1(n_272),
.B2(n_284),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_305),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_369),
.B(n_386),
.Y(n_419)
);

OA21x2_ASAP7_75t_L g372 ( 
.A1(n_308),
.A2(n_287),
.B(n_274),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_336),
.A2(n_334),
.B1(n_340),
.B2(n_294),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_298),
.B(n_257),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_294),
.A2(n_271),
.B1(n_257),
.B2(n_277),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_297),
.A2(n_293),
.B1(n_287),
.B2(n_276),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_298),
.B(n_255),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_382),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_255),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_338),
.A2(n_302),
.B1(n_307),
.B2(n_311),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_305),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_307),
.A2(n_301),
.B1(n_311),
.B2(n_309),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_387),
.B(n_366),
.Y(n_418)
);

OAI32xp33_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_300),
.A3(n_322),
.B1(n_317),
.B2(n_332),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_390),
.B(n_404),
.Y(n_435)
);

INVx13_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_391),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_339),
.B(n_313),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_392),
.A2(n_398),
.B(n_409),
.Y(n_432)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_349),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_393),
.B(n_399),
.Y(n_429)
);

INVx6_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_394),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_357),
.Y(n_442)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_374),
.Y(n_396)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

INVx13_ASAP7_75t_L g397 ( 
.A(n_353),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_397),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_387),
.B(n_299),
.Y(n_398)
);

AOI32xp33_ASAP7_75t_L g399 ( 
.A1(n_354),
.A2(n_325),
.A3(n_326),
.B1(n_331),
.B2(n_318),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g401 ( 
.A(n_375),
.B(n_319),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_401),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_356),
.B(n_303),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_405),
.Y(n_436)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_374),
.Y(n_403)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_371),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_351),
.B(n_303),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_406),
.B(n_410),
.C(n_347),
.Y(n_427)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_344),
.Y(n_407)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_407),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_383),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_414),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_345),
.B(n_350),
.C(n_354),
.Y(n_410)
);

BUFx5_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_413),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_376),
.B(n_381),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_379),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_354),
.B(n_376),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_423),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_417),
.A2(n_368),
.B1(n_372),
.B2(n_380),
.Y(n_453)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_418),
.Y(n_443)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_420),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_352),
.Y(n_421)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_362),
.B(n_367),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_346),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_354),
.A2(n_372),
.B(n_384),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_427),
.B(n_444),
.C(n_445),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_352),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_442),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_388),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_390),
.Y(n_470)
);

HAxp5_ASAP7_75t_SL g441 ( 
.A(n_389),
.B(n_355),
.CON(n_441),
.SN(n_441)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_441),
.B(n_449),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_410),
.B(n_357),
.C(n_385),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_395),
.B(n_382),
.C(n_346),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_402),
.B(n_386),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_405),
.B(n_369),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_450),
.B(n_419),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_453),
.A2(n_425),
.B1(n_399),
.B2(n_400),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_384),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_454),
.B(n_458),
.C(n_424),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_400),
.A2(n_378),
.B1(n_360),
.B2(n_373),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_455),
.A2(n_417),
.B1(n_434),
.B2(n_401),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_363),
.Y(n_456)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_456),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_419),
.B(n_363),
.Y(n_457)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_457),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_396),
.B(n_360),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_459),
.A2(n_460),
.B1(n_469),
.B2(n_476),
.Y(n_491)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_465),
.Y(n_498)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_456),
.Y(n_466)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_466),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_429),
.A2(n_425),
.B1(n_413),
.B2(n_403),
.Y(n_467)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_467),
.Y(n_506)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_457),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_468),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_435),
.A2(n_394),
.B1(n_421),
.B2(n_416),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_470),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_436),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_472),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_436),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_435),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_473),
.B(n_484),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_447),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_474),
.A2(n_412),
.B(n_398),
.Y(n_504)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_433),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_401),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_443),
.A2(n_401),
.B1(n_409),
.B2(n_392),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_478),
.A2(n_480),
.B1(n_482),
.B2(n_483),
.Y(n_503)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_433),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_430),
.B(n_416),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_485),
.Y(n_496)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_446),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_446),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_430),
.B(n_394),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_448),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_439),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_463),
.B(n_427),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_488),
.B(n_507),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_431),
.C(n_444),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_490),
.B(n_492),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_461),
.B(n_445),
.C(n_458),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_463),
.B(n_454),
.C(n_438),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_494),
.B(n_500),
.Y(n_522)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_499),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_438),
.C(n_432),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_432),
.C(n_442),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_501),
.B(n_505),
.Y(n_512)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_504),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_464),
.B(n_426),
.C(n_428),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_478),
.B(n_415),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_437),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_437),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_481),
.Y(n_526)
);

OAI21xp33_ASAP7_75t_L g510 ( 
.A1(n_506),
.A2(n_468),
.B(n_466),
.Y(n_510)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_510),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_513),
.B(n_514),
.Y(n_536)
);

BUFx12_ASAP7_75t_L g514 ( 
.A(n_497),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_498),
.A2(n_472),
.B1(n_475),
.B2(n_455),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_515),
.A2(n_434),
.B1(n_489),
.B2(n_485),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_508),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_523),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_493),
.B(n_490),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_519),
.B(n_520),
.Y(n_531)
);

BUFx24_ASAP7_75t_SL g520 ( 
.A(n_487),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_451),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_505),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_524),
.A2(n_525),
.B1(n_527),
.B2(n_462),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_495),
.A2(n_459),
.B1(n_453),
.B2(n_502),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_526),
.B(n_503),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_491),
.Y(n_527)
);

OA21x2_ASAP7_75t_SL g528 ( 
.A1(n_488),
.A2(n_479),
.B(n_462),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_528),
.B(n_496),
.C(n_428),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_492),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_533),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_532),
.B(n_539),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_511),
.B(n_494),
.C(n_500),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_522),
.B(n_509),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_534),
.B(n_538),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_535),
.B(n_540),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_526),
.B(n_507),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_516),
.C(n_521),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_542),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_513),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_517),
.B(n_527),
.C(n_496),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_543),
.B(n_544),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_510),
.B(n_443),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_536),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_546),
.B(n_543),
.Y(n_556)
);

FAx1_ASAP7_75t_L g547 ( 
.A(n_544),
.B(n_514),
.CI(n_452),
.CON(n_547),
.SN(n_547)
);

AOI31xp67_ASAP7_75t_L g562 ( 
.A1(n_547),
.A2(n_514),
.A3(n_542),
.B(n_448),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_531),
.B(n_533),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_539),
.Y(n_559)
);

AO21x1_ASAP7_75t_L g552 ( 
.A1(n_529),
.A2(n_452),
.B(n_484),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_552),
.A2(n_483),
.B(n_482),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_537),
.B(n_451),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_555),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_558),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_554),
.B(n_532),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_559),
.B(n_560),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_545),
.B(n_553),
.Y(n_560)
);

AOI322xp5_ASAP7_75t_L g563 ( 
.A1(n_561),
.A2(n_562),
.A3(n_547),
.B1(n_486),
.B2(n_552),
.C1(n_397),
.C2(n_391),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_563),
.B(n_565),
.Y(n_567)
);

AOI322xp5_ASAP7_75t_L g565 ( 
.A1(n_557),
.A2(n_553),
.A3(n_559),
.B1(n_480),
.B2(n_476),
.C1(n_550),
.C2(n_397),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_564),
.B(n_549),
.C(n_551),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_566),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_569),
.A2(n_570),
.B(n_448),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_567),
.B(n_407),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_420),
.C(n_423),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_360),
.B(n_391),
.Y(n_573)
);

BUFx24_ASAP7_75t_SL g574 ( 
.A(n_573),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_411),
.Y(n_575)
);


endmodule