module fake_jpeg_4598_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_10),
.C(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_1),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_22),
.B1(n_12),
.B2(n_20),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_36),
.B1(n_19),
.B2(n_21),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_12),
.B1(n_20),
.B2(n_19),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_14),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_18),
.Y(n_52)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

AOI32xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_29),
.A3(n_27),
.B1(n_31),
.B2(n_14),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_40),
.C(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_14),
.Y(n_63)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_54),
.B(n_37),
.C(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_63),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_17),
.B(n_16),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_41),
.B1(n_11),
.B2(n_13),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_69),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_65),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_43),
.B1(n_67),
.B2(n_5),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_75),
.B1(n_76),
.B2(n_62),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_49),
.C(n_48),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_74),
.B(n_37),
.Y(n_82)
);

XNOR2x1_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_52),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_54),
.B1(n_53),
.B2(n_50),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_44),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_64),
.B(n_56),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_79),
.B1(n_75),
.B2(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_63),
.B1(n_64),
.B2(n_56),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_2),
.B(n_4),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_13),
.B(n_11),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_74),
.B(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_89),
.B(n_90),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_80),
.C(n_87),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_77),
.C(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_77),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_2),
.C(n_4),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_8),
.B(n_10),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_100),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_98),
.B(n_9),
.C(n_6),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_5),
.B(n_6),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_104),
.A2(n_102),
.B(n_5),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_67),
.Y(n_106)
);


endmodule