module real_jpeg_6361_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_2),
.A2(n_28),
.B1(n_46),
.B2(n_49),
.Y(n_45)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_2),
.A2(n_49),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_2),
.A2(n_49),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_2),
.A2(n_49),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_2),
.A2(n_262),
.B(n_265),
.C(n_268),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_2),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_2),
.B(n_54),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_2),
.B(n_304),
.C(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_2),
.B(n_112),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_2),
.B(n_77),
.C(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_2),
.B(n_30),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_3),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_3),
.A2(n_79),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_3),
.A2(n_79),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_3),
.A2(n_79),
.B1(n_173),
.B2(n_177),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_4),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_4),
.A2(n_27),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_4),
.A2(n_27),
.B1(n_74),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_4),
.A2(n_27),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_5),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_5),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_5),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_5),
.A2(n_124),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_5),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_5),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_7),
.Y(n_96)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_8),
.Y(n_170)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_8),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_8),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_8),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_9),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_9),
.Y(n_267)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_13),
.Y(n_304)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_418),
.B(n_420),
.Y(n_18)
);

AO21x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_133),
.B(n_417),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_127),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_21),
.B(n_127),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_118),
.C(n_125),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_22),
.B(n_414),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.C(n_81),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_23),
.A2(n_141),
.B1(n_142),
.B2(n_155),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_23),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_23),
.B(n_142),
.C(n_156),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_23),
.B(n_243),
.C(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_23),
.A2(n_155),
.B1(n_243),
.B2(n_342),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_23),
.A2(n_155),
.B1(n_389),
.B2(n_390),
.Y(n_388)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_45),
.B2(n_50),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_24),
.A2(n_29),
.B1(n_45),
.B2(n_50),
.Y(n_231)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_28),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_29),
.A2(n_45),
.B1(n_50),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_29),
.A2(n_50),
.B1(n_119),
.B2(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_29),
.A2(n_45),
.B(n_50),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g419 ( 
.A1(n_29),
.A2(n_50),
.B(n_128),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_38),
.Y(n_29)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_31),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_32),
.Y(n_148)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_33),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_33),
.Y(n_154)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_40),
.Y(n_132)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_49),
.A2(n_144),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_51),
.A2(n_81),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_51),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_51),
.B(n_231),
.C(n_394),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_51),
.A2(n_392),
.B1(n_394),
.B2(n_401),
.Y(n_400)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_76),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_52),
.B(n_191),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_64),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_53),
.A2(n_64),
.B1(n_185),
.B2(n_190),
.Y(n_184)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_54),
.A2(n_199),
.B(n_206),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_54),
.B(n_186),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_54),
.A2(n_65),
.B1(n_76),
.B2(n_199),
.Y(n_242)
);

AO22x1_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_67),
.B1(n_70),
.B2(n_73),
.Y(n_66)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_58),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_58),
.Y(n_228)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_58),
.Y(n_275)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_61),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_61),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_65),
.B(n_191),
.Y(n_207)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_69),
.Y(n_205)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_75),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_75),
.Y(n_195)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_78),
.Y(n_193)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_81),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_89),
.B1(n_112),
.B2(n_113),
.Y(n_81)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_82),
.Y(n_395)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_89),
.B(n_230),
.Y(n_396)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_104),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_90),
.A2(n_104),
.B1(n_143),
.B2(n_149),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_90),
.A2(n_104),
.B1(n_143),
.B2(n_149),
.Y(n_243)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_104),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_97),
.B1(n_99),
.B2(n_102),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_101),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_104),
.A2(n_395),
.B(n_396),
.Y(n_394)
);

AOI22x1_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_110),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_118),
.B(n_125),
.Y(n_414)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_126),
.B(n_230),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_127),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_127),
.B(n_419),
.Y(n_421)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_412),
.B(n_416),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_383),
.B(n_409),
.Y(n_134)
);

OAI211xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_279),
.B(n_377),
.C(n_382),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_248),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_137),
.A2(n_248),
.B(n_378),
.C(n_381),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_232),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_138),
.B(n_232),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_196),
.C(n_214),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_139),
.B(n_196),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_156),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_141),
.A2(n_142),
.B1(n_217),
.B2(n_298),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_141),
.B(n_298),
.C(n_319),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_141),
.A2(n_142),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_142),
.B(n_231),
.C(n_352),
.Y(n_369)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_154),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_183),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_157),
.A2(n_183),
.B1(n_184),
.B2(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_157),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_163),
.B1(n_171),
.B2(n_180),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_159),
.A2(n_220),
.B(n_223),
.Y(n_219)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_162),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_163),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_164),
.A2(n_225),
.B1(n_271),
.B2(n_276),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_164),
.A2(n_221),
.B1(n_225),
.B2(n_271),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_170),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_209),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_177),
.Y(n_305)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_179),
.Y(n_272)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_183),
.A2(n_184),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_183),
.A2(n_184),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_184),
.B(n_270),
.C(n_312),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_184),
.B(n_334),
.C(n_336),
.Y(n_347)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_208),
.B2(n_213),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_208),
.Y(n_239)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_205),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_208),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_213),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_208),
.A2(n_238),
.B(n_239),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_209),
.B(n_225),
.Y(n_327)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_229),
.C(n_231),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_254),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_217),
.A2(n_298),
.B1(n_299),
.B2(n_306),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_217),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_217),
.A2(n_219),
.B1(n_298),
.B2(n_368),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_219),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_231),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_231),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_231),
.A2(n_255),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_231),
.A2(n_255),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_231),
.A2(n_255),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_231),
.B(n_388),
.C(n_393),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_246),
.B2(n_247),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_240),
.B1(n_241),
.B2(n_245),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_240),
.B(n_245),
.C(n_247),
.Y(n_408)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_243),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_243),
.A2(n_338),
.B1(n_339),
.B2(n_342),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_243),
.Y(n_342)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_244),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_244),
.A2(n_398),
.B1(n_402),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_249),
.B(n_251),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.C(n_259),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_252),
.A2(n_253),
.B1(n_257),
.B2(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_257),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_259),
.B(n_375),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_260),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_269),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_261),
.A2(n_269),
.B1(n_270),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_261),
.Y(n_359)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_SL g266 ( 
.A(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_269),
.A2(n_270),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_361),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_346),
.B(n_360),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_331),
.B(n_345),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_316),
.B(n_330),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_308),
.B(n_315),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_295),
.B(n_307),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_292),
.B(n_294),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_291),
.A2(n_296),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_296),
.B(n_340),
.C(n_342),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_306),
.Y(n_314)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_314),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_314),
.Y(n_315)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_318),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_329),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_327),
.B2(n_328),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_328),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_344),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_344),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_336),
.B1(n_337),
.B2(n_343),
.Y(n_332)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_348),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_354),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_356),
.C(n_357),
.Y(n_370)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NOR2x1_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_371),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_370),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_370),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_369),
.C(n_373),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_371),
.A2(n_379),
.B(n_380),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_374),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_404),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_410),
.B(n_411),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_397),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_397),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_393),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_394),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_402),
.C(n_403),
.Y(n_397)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_398),
.Y(n_407)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_406),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_405),
.B(n_408),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_415),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_413),
.B(n_415),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_421),
.Y(n_420)
);


endmodule