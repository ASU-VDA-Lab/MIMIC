module real_jpeg_24475_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_210;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_1),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_1),
.B(n_75),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_1),
.B(n_31),
.C(n_49),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_1),
.B(n_121),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_1),
.A2(n_91),
.B1(n_92),
.B2(n_231),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_2),
.A2(n_45),
.B1(n_67),
.B2(n_68),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_45),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_3),
.A2(n_35),
.B1(n_67),
.B2(n_68),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_3),
.A2(n_35),
.B1(n_42),
.B2(n_43),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_3),
.A2(n_35),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_4),
.A2(n_32),
.B1(n_60),
.B2(n_71),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_4),
.A2(n_32),
.B1(n_67),
.B2(n_68),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_4),
.A2(n_32),
.B1(n_42),
.B2(n_43),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_7),
.A2(n_59),
.B1(n_67),
.B2(n_68),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_59),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_59),
.Y(n_254)
);

INVx8_ASAP7_75t_SL g66 ( 
.A(n_8),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_9),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_163),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_163),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_163),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_54),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_10),
.A2(n_54),
.B1(n_67),
.B2(n_68),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_115),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_14),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_115),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_115),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_115),
.Y(n_224)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_15),
.Y(n_92)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_146),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_144),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_116),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_19),
.B(n_116),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_88),
.C(n_99),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_20),
.A2(n_21),
.B1(n_88),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_22),
.B(n_76),
.C(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_25),
.A2(n_91),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_29),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_29),
.A2(n_91),
.B(n_104),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_37),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_31),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_30),
.B(n_236),
.Y(n_235)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_33),
.A2(n_177),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_34),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_36),
.A2(n_103),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_36),
.A2(n_191),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_37),
.Y(n_179)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_52),
.B2(n_53),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_41),
.A2(n_51),
.B(n_108),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_43),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_42),
.A2(n_80),
.B(n_245),
.C(n_247),
.Y(n_244)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_43),
.B(n_206),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_L g247 ( 
.A(n_43),
.B(n_67),
.C(n_79),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_46),
.B(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_46),
.A2(n_96),
.B(n_125),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_46),
.A2(n_52),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_46),
.A2(n_52),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_47),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_47),
.A2(n_51),
.B1(n_210),
.B2(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_47),
.A2(n_124),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_51),
.B(n_159),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_52),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_53),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_76),
.B1(n_77),
.B2(n_87),
.Y(n_55)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_62),
.B(n_73),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_58),
.A2(n_63),
.B1(n_75),
.B2(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_62),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_62),
.A2(n_64),
.B1(n_162),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_63),
.A2(n_75),
.B1(n_158),
.B2(n_161),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_66),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_65),
.A2(n_68),
.B(n_160),
.C(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_66),
.B(n_67),
.C(n_72),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_68),
.B1(n_79),
.B2(n_80),
.Y(n_84)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

HAxp5_ASAP7_75t_SL g246 ( 
.A(n_68),
.B(n_159),
.CON(n_246),
.SN(n_246)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_72),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_75),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_82),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_78),
.A2(n_171),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_83),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_83),
.A2(n_121),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_83),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_83),
.A2(n_121),
.B1(n_196),
.B2(n_246),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_88),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_98),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_90),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_93),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_91),
.A2(n_224),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_99),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_110),
.C(n_113),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_100),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_107),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_107),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_105),
.Y(n_232)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_106),
.B(n_159),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_110),
.B(n_113),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_111),
.B(n_121),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_114),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_127),
.B1(n_139),
.B2(n_140),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_123),
.B(n_126),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_119),
.B(n_123),
.Y(n_126)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_138),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_136),
.B(n_159),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_141),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_287),
.B(n_292),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_198),
.B(n_278),
.C(n_286),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_183),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_149),
.B(n_183),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_164),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_151),
.B(n_152),
.C(n_164),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.C(n_157),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_185),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_173),
.B2(n_182),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_167),
.B(n_169),
.C(n_182),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_180),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_175),
.B1(n_180),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_184),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_186),
.B(n_188),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_189),
.Y(n_263)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_194),
.B(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_277),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_272),
.B(n_276),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_257),
.B(n_271),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_240),
.B(n_256),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_220),
.B(n_239),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_211),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_211),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_207),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_215),
.C(n_218),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_227),
.B(n_238),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_226),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_237),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_255),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_255),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_250),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_251),
.C(n_252),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_249),
.Y(n_266)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_259),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_264),
.B2(n_265),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_267),
.C(n_269),
.Y(n_275)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_275),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_285),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_283),
.C(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);


endmodule