module fake_jpeg_7835_n_46 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_46);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_46;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_24),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_25),
.A2(n_28),
.B(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_11),
.C(n_17),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_6),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_4),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_19),
.B(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_36),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_27),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_37),
.B(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_8),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_10),
.B(n_12),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_32),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_35),
.B1(n_41),
.B2(n_40),
.Y(n_45)
);

AOI322xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_14),
.A3(n_16),
.B1(n_18),
.B2(n_39),
.C1(n_40),
.C2(n_42),
.Y(n_46)
);


endmodule