module real_jpeg_23665_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_286;
wire n_215;
wire n_288;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_293;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_216;
wire n_167;
wire n_213;
wire n_202;
wire n_133;
wire n_179;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

INVx3_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_1),
.A2(n_29),
.B1(n_43),
.B2(n_44),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_3),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_5),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_5),
.A2(n_66),
.B1(n_73),
.B2(n_81),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_66),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_66),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_7),
.A2(n_75),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_7),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_136),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_136),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_136),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_10),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_10),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_71),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_71),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_71),
.Y(n_243)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_12),
.A2(n_81),
.B1(n_87),
.B2(n_89),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_12),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_89),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_89),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_89),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_13),
.B(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_13),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_13),
.B(n_83),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_13),
.B(n_44),
.C(n_58),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_184),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_13),
.B(n_156),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_184),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_13),
.B(n_28),
.C(n_49),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_13),
.A2(n_30),
.B(n_244),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_15),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_99)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_16),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_16),
.B(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_16),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_138),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_117),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_20),
.B(n_117),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_90),
.B2(n_116),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.C(n_68),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_23),
.A2(n_24),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_25),
.A2(n_39),
.B1(n_40),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_25),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_26),
.A2(n_30),
.B1(n_36),
.B2(n_125),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_28),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_27),
.B(n_269),
.Y(n_268)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_30),
.A2(n_34),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_30),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_30),
.A2(n_165),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_30),
.B(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_30),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_31),
.Y(n_166)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_38),
.B(n_184),
.Y(n_269)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_42),
.A2(n_51),
.B1(n_96),
.B2(n_128),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_44),
.B(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_47),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_47),
.A2(n_54),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_51),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_51),
.A2(n_128),
.B(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_51),
.A2(n_180),
.B(n_217),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_51),
.B(n_184),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_54),
.B(n_181),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_55),
.B(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_65),
.B2(n_67),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_56),
.A2(n_57),
.B1(n_67),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_56),
.A2(n_153),
.B(n_155),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_56),
.A2(n_155),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_57),
.A2(n_65),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_57),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_57),
.A2(n_131),
.B(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_62),
.B1(n_79),
.B2(n_80),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g158 ( 
.A1(n_61),
.A2(n_72),
.A3(n_80),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_62),
.B(n_79),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_62),
.B(n_210),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_76),
.B(n_84),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_70),
.A2(n_77),
.B1(n_83),
.B2(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_72),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_78)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_77),
.A2(n_85),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_113),
.B(n_114),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_82),
.A2(n_114),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_101),
.B2(n_102),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B(n_100),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_95),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_96),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_96),
.A2(n_232),
.B(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.C(n_122),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_121),
.Y(n_168)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.C(n_134),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_124),
.B(n_127),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_154),
.B1(n_156),
.B2(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_135),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_169),
.B(n_293),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_167),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_142),
.B(n_167),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.C(n_149),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_147),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_149),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_157),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_152),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_162),
.Y(n_186)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_163),
.A2(n_255),
.B1(n_257),
.B2(n_259),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_166),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_202),
.B(n_287),
.C(n_292),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_196),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_196),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_186),
.C(n_187),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_172),
.A2(n_173),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_178),
.C(n_182),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_177),
.Y(n_189)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_186),
.B(n_187),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_192),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_197),
.B(n_200),
.C(n_201),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_281),
.B(n_286),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_233),
.B(n_280),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_222),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_207),
.B(n_222),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_215),
.C(n_219),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_208),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_211),
.Y(n_229)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_215),
.A2(n_219),
.B1(n_220),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_215),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_218),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_228),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_223),
.B(n_229),
.C(n_230),
.Y(n_285)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_274),
.B(n_279),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_252),
.B(n_273),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_246),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_246),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_278)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_243),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_248),
.B1(n_250),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_250),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_262),
.B(n_272),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_260),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_260),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_258),
.B(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_267),
.B(n_271),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_265),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_278),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);


endmodule