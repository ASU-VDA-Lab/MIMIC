module real_jpeg_24733_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_179;
wire n_244;
wire n_167;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_59),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_1),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_48),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_5),
.A2(n_48),
.B1(n_66),
.B2(n_67),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_5),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_6),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_6),
.A2(n_38),
.B1(n_66),
.B2(n_67),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_8),
.B(n_66),
.C(n_85),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_76),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_8),
.B(n_60),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_8),
.A2(n_68),
.B1(n_72),
.B2(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_8),
.B(n_99),
.Y(n_217)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_71),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_11),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_11),
.A2(n_66),
.B1(n_67),
.B2(n_93),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_93),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_13),
.A2(n_44),
.B1(n_53),
.B2(n_54),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_13),
.A2(n_44),
.B1(n_66),
.B2(n_67),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_65),
.Y(n_108)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_15),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_139),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_111),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_19),
.B(n_111),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_80),
.C(n_101),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_20),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_61),
.B2(n_79),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_45),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_23),
.B(n_45),
.C(n_79),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_26),
.B1(n_37),
.B2(n_42),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_25),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_25),
.A2(n_43),
.B1(n_99),
.B2(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_28),
.B1(n_33),
.B2(n_36),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_27),
.A2(n_30),
.B(n_75),
.C(n_78),
.Y(n_74)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_28),
.B(n_29),
.C(n_77),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_29),
.A2(n_30),
.B1(n_52),
.B2(n_55),
.Y(n_56)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g194 ( 
.A(n_30),
.B(n_76),
.CON(n_194),
.SN(n_194)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_30),
.B(n_53),
.C(n_55),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_39),
.A2(n_75),
.B(n_76),
.Y(n_98)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B(n_57),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_47),
.A2(n_50),
.B1(n_60),
.B2(n_96),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_49),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_49),
.A2(n_51),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_50),
.A2(n_60),
.B1(n_194),
.B2(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_52),
.A2(n_54),
.B(n_194),
.C(n_195),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_54),
.B1(n_85),
.B2(n_87),
.Y(n_84)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_54),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_58),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_60),
.B(n_123),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_74),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_62),
.B(n_74),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_68),
.B1(n_70),
.B2(n_72),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_64),
.A2(n_130),
.B(n_169),
.Y(n_218)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_69),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_67),
.B1(n_85),
.B2(n_87),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_67),
.B(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_70),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_68),
.B(n_106),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_68),
.A2(n_128),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_68),
.A2(n_168),
.B1(n_176),
.B2(n_185),
.Y(n_184)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_69),
.Y(n_169)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_69),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_76),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_76),
.B(n_88),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_80),
.A2(n_101),
.B1(n_102),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_80),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_95),
.C(n_97),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_81),
.A2(n_82),
.B1(n_95),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_89),
.B(n_91),
.Y(n_82)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_83),
.A2(n_88),
.B1(n_108),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_83),
.A2(n_88),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_83),
.A2(n_88),
.B1(n_153),
.B2(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_83),
.A2(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_88),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_90),
.B(n_94),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_94),
.A2(n_110),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_95),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_96),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_97),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_107),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_107),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_105),
.A2(n_129),
.B(n_166),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_136),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_124),
.B1(n_134),
.B2(n_135),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_131),
.B2(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_244),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_239),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_229),
.B(n_238),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_207),
.B(n_228),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_190),
.B(n_206),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_163),
.B(n_189),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_154),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_162),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_173),
.B(n_188),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_182),
.B(n_187),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_183),
.B(n_184),
.Y(n_187)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_205),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_205),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_199),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_200),
.C(n_203),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_193),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_220),
.B2(n_221),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_223),
.C(n_226),
.Y(n_237)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_216),
.C(n_219),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_218),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_237),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);


endmodule