module fake_netlist_1_4280_n_708 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_708);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_708;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_6), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_82), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_63), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_44), .Y(n_90) );
INVx3_ASAP7_75t_L g91 ( .A(n_28), .Y(n_91) );
NOR2xp67_ASAP7_75t_L g92 ( .A(n_3), .B(n_37), .Y(n_92) );
XNOR2x1_ASAP7_75t_L g93 ( .A(n_13), .B(n_3), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_17), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_13), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_76), .Y(n_96) );
INVx1_ASAP7_75t_SL g97 ( .A(n_14), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_22), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_85), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_58), .Y(n_100) );
CKINVDCx14_ASAP7_75t_R g101 ( .A(n_36), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_16), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_64), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_57), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_55), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_32), .Y(n_106) );
INVx3_ASAP7_75t_L g107 ( .A(n_39), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_15), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_19), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_53), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_59), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_72), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_62), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_7), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_1), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_79), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_83), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_2), .Y(n_119) );
XOR2xp5_ASAP7_75t_L g120 ( .A(n_75), .B(n_27), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_41), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_23), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_26), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_121), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_88), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_121), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_121), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_121), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_91), .B(n_0), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_116), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_120), .A2(n_102), .B1(n_109), .B2(n_119), .Y(n_132) );
INVx4_ASAP7_75t_L g133 ( .A(n_91), .Y(n_133) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_91), .A2(n_46), .B(n_84), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_91), .B(n_0), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_107), .B(n_1), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_107), .B(n_47), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_110), .B(n_2), .Y(n_139) );
BUFx8_ASAP7_75t_L g140 ( .A(n_121), .Y(n_140) );
AO22x1_ASAP7_75t_L g141 ( .A1(n_102), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_107), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_121), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_133), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_133), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_135), .B(n_110), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_135), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_133), .B(n_101), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_133), .B(n_87), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_135), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_136), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_136), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_125), .B(n_99), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_125), .B(n_104), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_142), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_135), .B(n_131), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_142), .Y(n_160) );
OR2x2_ASAP7_75t_L g161 ( .A(n_139), .B(n_93), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_130), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_124), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_124), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_138), .A2(n_145), .B1(n_131), .B2(n_143), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_124), .Y(n_167) );
AND2x6_ASAP7_75t_L g168 ( .A(n_139), .B(n_90), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_143), .B(n_116), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_124), .Y(n_170) );
OR2x2_ASAP7_75t_L g171 ( .A(n_145), .B(n_93), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_124), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_130), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_130), .Y(n_176) );
INVx5_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_129), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_126), .Y(n_179) );
BUFx10_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
NOR3xp33_ASAP7_75t_L g181 ( .A(n_132), .B(n_141), .C(n_97), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g182 ( .A1(n_168), .A2(n_138), .B1(n_137), .B2(n_140), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_178), .B(n_132), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
OAI221xp5_ASAP7_75t_L g185 ( .A1(n_171), .A2(n_109), .B1(n_115), .B2(n_119), .C(n_95), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_172), .Y(n_186) );
NOR3x1_ASAP7_75t_L g187 ( .A(n_161), .B(n_141), .C(n_115), .Y(n_187) );
NOR3xp33_ASAP7_75t_L g188 ( .A(n_161), .B(n_181), .C(n_171), .Y(n_188) );
NOR2x2_ASAP7_75t_L g189 ( .A(n_168), .B(n_120), .Y(n_189) );
AOI22xp33_ASAP7_75t_SL g190 ( .A1(n_168), .A2(n_138), .B1(n_95), .B2(n_134), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_154), .B(n_90), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_178), .B(n_103), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_169), .B(n_134), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_156), .B(n_140), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_169), .B(n_111), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_147), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_148), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_151), .B(n_168), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_172), .Y(n_199) );
NAND3xp33_ASAP7_75t_L g200 ( .A(n_166), .B(n_108), .C(n_94), .Y(n_200) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_173), .B(n_92), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_159), .A2(n_114), .B(n_108), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_168), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_168), .A2(n_113), .B1(n_94), .B2(n_98), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_154), .B(n_98), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_168), .B(n_112), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
INVx8_ASAP7_75t_L g208 ( .A(n_177), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_147), .Y(n_209) );
AOI221xp5_ASAP7_75t_L g210 ( .A1(n_152), .A2(n_113), .B1(n_114), .B2(n_123), .C(n_118), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_150), .B(n_117), .Y(n_211) );
AOI22xp5_ASAP7_75t_SL g212 ( .A1(n_152), .A2(n_123), .B1(n_104), .B2(n_122), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_173), .B(n_122), .Y(n_213) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_177), .B(n_96), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_153), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_153), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_149), .A2(n_96), .B(n_100), .C(n_105), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_149), .A2(n_157), .B1(n_175), .B2(n_176), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_154), .B(n_100), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_149), .B(n_105), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_154), .A2(n_106), .B1(n_92), .B2(n_127), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_176), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_162), .A2(n_106), .B1(n_128), .B2(n_127), .Y(n_224) );
AO21x1_ASAP7_75t_L g225 ( .A1(n_193), .A2(n_162), .B(n_160), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_SL g226 ( .A1(n_194), .A2(n_160), .B(n_146), .C(n_158), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_190), .B(n_162), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_182), .B(n_162), .Y(n_228) );
NOR2xp67_ASAP7_75t_L g229 ( .A(n_183), .B(n_4), .Y(n_229) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_208), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_198), .B(n_177), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_188), .A2(n_155), .B1(n_158), .B2(n_146), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_192), .B(n_155), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_203), .A2(n_177), .B1(n_180), .B2(n_126), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_185), .A2(n_164), .B(n_165), .C(n_170), .Y(n_235) );
NAND3xp33_ASAP7_75t_L g236 ( .A(n_210), .B(n_177), .C(n_127), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_215), .Y(n_237) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_219), .A2(n_170), .B(n_179), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_197), .B(n_177), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_208), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_195), .B(n_180), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_204), .A2(n_180), .B1(n_144), .B2(n_128), .Y(n_243) );
OR2x6_ASAP7_75t_L g244 ( .A(n_201), .B(n_180), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_193), .B(n_126), .Y(n_245) );
NAND2x1p5_ASAP7_75t_L g246 ( .A(n_199), .B(n_126), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_219), .A2(n_179), .B(n_164), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_191), .A2(n_165), .B(n_167), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_213), .B(n_5), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_216), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_187), .B(n_7), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_218), .A2(n_126), .B1(n_127), .B2(n_128), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_186), .B(n_144), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_191), .A2(n_174), .B(n_167), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_220), .A2(n_174), .B(n_167), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_213), .B(n_8), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_196), .A2(n_144), .B(n_128), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_216), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_226), .A2(n_205), .B(n_186), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_256), .B(n_212), .Y(n_260) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_255), .A2(n_222), .B(n_217), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_230), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_256), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_184), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_251), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_245), .A2(n_205), .B(n_211), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_245), .A2(n_208), .B(n_223), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_230), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_249), .B(n_201), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_238), .A2(n_202), .B(n_224), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_228), .A2(n_208), .B(n_207), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_230), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_225), .A2(n_221), .B(n_200), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_230), .B(n_199), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_240), .Y(n_275) );
NAND3xp33_ASAP7_75t_L g276 ( .A(n_236), .B(n_214), .C(n_206), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_244), .Y(n_277) );
NOR2xp33_ASAP7_75t_SL g278 ( .A(n_240), .B(n_189), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_227), .A2(n_209), .B(n_196), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_233), .B(n_209), .Y(n_280) );
INVx5_ASAP7_75t_L g281 ( .A(n_240), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_264), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_278), .A2(n_229), .B1(n_232), .B2(n_227), .Y(n_283) );
NOR2x1_ASAP7_75t_R g284 ( .A(n_281), .B(n_189), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_260), .B(n_265), .Y(n_285) );
AO31x2_ASAP7_75t_L g286 ( .A1(n_271), .A2(n_252), .A3(n_243), .B(n_250), .Y(n_286) );
AND3x2_ASAP7_75t_L g287 ( .A(n_263), .B(n_258), .C(n_241), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_266), .A2(n_228), .B(n_254), .Y(n_288) );
INVx4_ASAP7_75t_L g289 ( .A(n_281), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_264), .Y(n_290) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_279), .A2(n_257), .B(n_253), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_273), .A2(n_232), .B(n_235), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_279), .A2(n_248), .B(n_246), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_272), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_273), .A2(n_246), .B(n_247), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_261), .A2(n_253), .B(n_231), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_269), .B(n_277), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_280), .B(n_244), .Y(n_298) );
OA21x2_ASAP7_75t_L g299 ( .A1(n_261), .A2(n_231), .B(n_239), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_267), .A2(n_242), .B(n_214), .C(n_240), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_281), .Y(n_301) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_270), .A2(n_242), .B(n_234), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_272), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_276), .A2(n_244), .B(n_144), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_281), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_303), .Y(n_306) );
OR2x6_ASAP7_75t_L g307 ( .A(n_289), .B(n_272), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_292), .A2(n_259), .B(n_270), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_289), .B(n_281), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_282), .B(n_268), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_282), .Y(n_312) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_296), .A2(n_275), .B(n_272), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_284), .B(n_277), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_290), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_290), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_294), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_303), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_296), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_294), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_294), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_294), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_292), .A2(n_274), .B(n_127), .Y(n_326) );
AO31x2_ASAP7_75t_L g327 ( .A1(n_288), .A2(n_144), .A3(n_128), .B(n_275), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_289), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_285), .B(n_262), .Y(n_329) );
BUFx12f_ASAP7_75t_L g330 ( .A(n_289), .Y(n_330) );
CKINVDCx16_ASAP7_75t_R g331 ( .A(n_297), .Y(n_331) );
OR2x6_ASAP7_75t_L g332 ( .A(n_304), .B(n_275), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_299), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_299), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_301), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_301), .B(n_262), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_299), .Y(n_337) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_304), .A2(n_274), .B(n_275), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_305), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_295), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_305), .B(n_274), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_298), .B(n_8), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_299), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_295), .B(n_51), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_335), .B(n_298), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_330), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_342), .B(n_283), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_315), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_310), .B(n_283), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_310), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_328), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_316), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_316), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_330), .Y(n_356) );
NOR2x1_ASAP7_75t_L g357 ( .A(n_328), .B(n_291), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_312), .B(n_302), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_312), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_317), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_342), .B(n_286), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_319), .B(n_286), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_333), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_327), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_331), .B(n_284), .Y(n_367) );
OR2x2_ASAP7_75t_SL g368 ( .A(n_331), .B(n_302), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_306), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_311), .B(n_302), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_311), .B(n_302), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_329), .B(n_287), .Y(n_373) );
INVx5_ASAP7_75t_SL g374 ( .A(n_309), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_327), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_319), .B(n_286), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_327), .Y(n_378) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_339), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_328), .Y(n_380) );
AOI22xp33_ASAP7_75t_SL g381 ( .A1(n_328), .A2(n_291), .B1(n_293), .B2(n_286), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_327), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_306), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_341), .B(n_286), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_334), .Y(n_385) );
OR2x6_ASAP7_75t_L g386 ( .A(n_332), .B(n_293), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_339), .B(n_286), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_334), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_307), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_341), .B(n_9), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_307), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_309), .B(n_300), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_336), .B(n_9), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_337), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_343), .B(n_291), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_343), .B(n_10), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_320), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_309), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_336), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_307), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_309), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_308), .B(n_10), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_307), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_314), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_308), .B(n_11), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_323), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_320), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_323), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_370), .B(n_326), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_370), .B(n_326), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_379), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_372), .B(n_308), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_387), .B(n_340), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_348), .Y(n_414) );
AND2x4_ASAP7_75t_SL g415 ( .A(n_401), .B(n_344), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_387), .B(n_340), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_371), .B(n_399), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_349), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_396), .B(n_338), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_398), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_365), .B(n_338), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_349), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_365), .B(n_338), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_376), .B(n_325), .Y(n_424) );
NOR2x1_ASAP7_75t_L g425 ( .A(n_346), .B(n_344), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_376), .B(n_385), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_385), .B(n_325), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_394), .B(n_313), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_394), .B(n_313), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_369), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_345), .B(n_332), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_396), .B(n_344), .Y(n_432) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_403), .B(n_344), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_393), .B(n_332), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_383), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_398), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_357), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_346), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_345), .B(n_332), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_388), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_393), .B(n_332), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_356), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_353), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_406), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_406), .B(n_324), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_353), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_361), .B(n_324), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_354), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_389), .B(n_322), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_397), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_354), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_356), .B(n_321), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_355), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_389), .B(n_321), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_389), .B(n_318), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_395), .B(n_11), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_390), .B(n_12), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_395), .B(n_12), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_361), .B(n_14), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_360), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_358), .B(n_15), .Y(n_461) );
INVxp67_ASAP7_75t_L g462 ( .A(n_390), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_383), .B(n_16), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_347), .B(n_18), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_408), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_358), .B(n_20), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_408), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_351), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_384), .B(n_21), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_351), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_380), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_397), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_380), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_407), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_347), .B(n_24), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_359), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_359), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_402), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_407), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_402), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_352), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_350), .B(n_25), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_350), .B(n_29), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_374), .B(n_30), .Y(n_484) );
INVxp67_ASAP7_75t_L g485 ( .A(n_367), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_405), .B(n_31), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_373), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_362), .B(n_33), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_362), .B(n_34), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_374), .B(n_35), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_377), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_377), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_456), .B(n_400), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_412), .B(n_357), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_411), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_412), .B(n_366), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_415), .B(n_386), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_417), .B(n_374), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_456), .B(n_458), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_487), .B(n_404), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_430), .Y(n_501) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_433), .B(n_403), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_458), .B(n_400), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_426), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_426), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_413), .B(n_378), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_415), .B(n_386), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_472), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_462), .B(n_391), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_478), .B(n_374), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_438), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_480), .B(n_391), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_442), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_452), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_413), .B(n_378), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_416), .B(n_375), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_435), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_461), .B(n_403), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_414), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_491), .B(n_403), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_416), .B(n_352), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_420), .B(n_352), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_461), .B(n_381), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_420), .B(n_386), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_409), .B(n_363), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_418), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_436), .B(n_386), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_436), .B(n_386), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_492), .B(n_392), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_485), .B(n_368), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_422), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_452), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_459), .B(n_392), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_472), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_465), .B(n_392), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_447), .B(n_368), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_442), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_467), .B(n_382), .Y(n_539) );
NOR2xp33_ASAP7_75t_SL g540 ( .A(n_433), .B(n_382), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_443), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_446), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_425), .B(n_375), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_448), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_451), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_471), .B(n_431), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_453), .B(n_366), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_439), .B(n_364), .Y(n_548) );
NAND2xp33_ASAP7_75t_L g549 ( .A(n_484), .B(n_364), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_474), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_474), .Y(n_551) );
NAND2x1p5_ASAP7_75t_L g552 ( .A(n_486), .B(n_38), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_460), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_409), .B(n_40), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_410), .B(n_42), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_432), .B(n_43), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_486), .B(n_45), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_457), .B(n_48), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_479), .Y(n_559) );
OR2x6_ASAP7_75t_L g560 ( .A(n_473), .B(n_49), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_479), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_424), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_427), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_427), .B(n_50), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_444), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_419), .B(n_52), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_421), .B(n_54), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_444), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_440), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_421), .B(n_56), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_440), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_445), .B(n_60), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_495), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_512), .B(n_463), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_514), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_504), .B(n_423), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_540), .A2(n_434), .B1(n_441), .B2(n_469), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_495), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_546), .B(n_481), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_518), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_518), .Y(n_581) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_531), .A2(n_475), .B(n_464), .C(n_437), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_505), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_538), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_520), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_562), .B(n_428), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_527), .Y(n_587) );
INVx3_ASAP7_75t_L g588 ( .A(n_502), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_532), .Y(n_589) );
CKINVDCx16_ASAP7_75t_R g590 ( .A(n_560), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_541), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g592 ( .A1(n_531), .A2(n_489), .B(n_488), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_558), .B(n_469), .C(n_489), .D(n_488), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_500), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_563), .B(n_428), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_542), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g597 ( .A1(n_560), .A2(n_490), .B(n_466), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_496), .B(n_429), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_496), .B(n_470), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_499), .A2(n_429), .B1(n_482), .B2(n_483), .C(n_466), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_544), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_560), .A2(n_483), .B(n_482), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_526), .B(n_445), .Y(n_603) );
INVx2_ASAP7_75t_SL g604 ( .A(n_515), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_498), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_526), .B(n_477), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_502), .Y(n_607) );
NOR2xp67_ASAP7_75t_L g608 ( .A(n_515), .B(n_476), .Y(n_608) );
INVx3_ASAP7_75t_L g609 ( .A(n_497), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g610 ( .A(n_533), .B(n_455), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_545), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_501), .B(n_468), .Y(n_612) );
OR2x6_ASAP7_75t_L g613 ( .A(n_497), .B(n_455), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_553), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_522), .B(n_454), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_543), .A2(n_454), .B(n_449), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_503), .B(n_449), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_524), .A2(n_449), .B(n_174), .Y(n_618) );
NAND2x1_ASAP7_75t_SL g619 ( .A(n_497), .B(n_61), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_501), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_559), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_537), .B(n_506), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_533), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_539), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_523), .Y(n_625) );
OAI33xp33_ASAP7_75t_L g626 ( .A1(n_510), .A2(n_65), .A3(n_66), .B1(n_67), .B2(n_68), .B3(n_69), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_547), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_494), .A2(n_174), .B1(n_167), .B2(n_73), .C(n_74), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_513), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_516), .B(n_71), .Y(n_630) );
AOI222xp33_ASAP7_75t_L g631 ( .A1(n_594), .A2(n_494), .B1(n_493), .B2(n_534), .C1(n_558), .C2(n_517), .Y(n_631) );
OAI21xp5_ASAP7_75t_SL g632 ( .A1(n_593), .A2(n_552), .B(n_557), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_608), .B(n_508), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_573), .A2(n_552), .B(n_557), .C(n_543), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_598), .B(n_517), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_599), .B(n_548), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_574), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_590), .A2(n_508), .B1(n_519), .B2(n_511), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_578), .B(n_530), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g640 ( .A(n_620), .B(n_549), .C(n_555), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_612), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_593), .A2(n_536), .B(n_554), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_624), .B(n_565), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_627), .B(n_568), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_608), .B(n_508), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_585), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_629), .B(n_569), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_587), .Y(n_648) );
OAI332xp33_ASAP7_75t_L g649 ( .A1(n_584), .A2(n_521), .A3(n_556), .B1(n_566), .B2(n_570), .B3(n_567), .C1(n_571), .C2(n_535), .Y(n_649) );
AND2x4_ASAP7_75t_L g650 ( .A(n_613), .B(n_529), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_602), .A2(n_549), .B(n_525), .Y(n_651) );
NOR2x1_ASAP7_75t_L g652 ( .A(n_588), .B(n_555), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_589), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_583), .B(n_509), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_591), .Y(n_655) );
NOR3xp33_ASAP7_75t_SL g656 ( .A(n_582), .B(n_592), .C(n_626), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_596), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_601), .Y(n_658) );
AOI32xp33_ASAP7_75t_L g659 ( .A1(n_588), .A2(n_528), .A3(n_564), .B1(n_572), .B2(n_507), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_580), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_611), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_581), .B(n_550), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_614), .A2(n_561), .B1(n_551), .B2(n_535), .C(n_509), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_621), .Y(n_664) );
AOI21xp5_ASAP7_75t_SL g665 ( .A1(n_634), .A2(n_618), .B(n_592), .Y(n_665) );
O2A1O1Ixp33_ASAP7_75t_L g666 ( .A1(n_656), .A2(n_575), .B(n_618), .C(n_604), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_642), .A2(n_600), .B1(n_605), .B2(n_607), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_643), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_644), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_632), .A2(n_619), .B(n_607), .C(n_609), .Y(n_670) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_642), .A2(n_597), .B(n_616), .C(n_609), .Y(n_671) );
AOI31xp33_ASAP7_75t_L g672 ( .A1(n_652), .A2(n_623), .A3(n_610), .B(n_577), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_637), .A2(n_595), .B1(n_586), .B2(n_576), .C(n_579), .Y(n_673) );
OAI321xp33_ASAP7_75t_L g674 ( .A1(n_659), .A2(n_577), .A3(n_613), .B1(n_622), .B2(n_630), .C(n_625), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_633), .A2(n_613), .B1(n_603), .B2(n_606), .Y(n_675) );
INVx3_ASAP7_75t_L g676 ( .A(n_633), .Y(n_676) );
OAI211xp5_ASAP7_75t_L g677 ( .A1(n_631), .A2(n_628), .B(n_617), .C(n_615), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_636), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_640), .B(n_645), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_646), .A2(n_77), .B(n_78), .C(n_80), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_651), .B(n_81), .C(n_86), .D(n_663), .Y(n_681) );
AOI222xp33_ASAP7_75t_L g682 ( .A1(n_648), .A2(n_655), .B1(n_661), .B2(n_658), .C1(n_657), .C2(n_653), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_649), .A2(n_647), .B(n_654), .Y(n_683) );
NAND2x1_ASAP7_75t_L g684 ( .A(n_650), .B(n_660), .Y(n_684) );
OAI22xp33_ASAP7_75t_SL g685 ( .A1(n_639), .A2(n_664), .B1(n_635), .B2(n_662), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_642), .B(n_641), .Y(n_686) );
OAI211xp5_ASAP7_75t_L g687 ( .A1(n_632), .A2(n_656), .B(n_642), .C(n_634), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_642), .A2(n_632), .B1(n_656), .B2(n_659), .C(n_638), .Y(n_688) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_687), .B(n_688), .Y(n_689) );
OAI21xp5_ASAP7_75t_L g690 ( .A1(n_666), .A2(n_665), .B(n_674), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_667), .A2(n_679), .B1(n_671), .B2(n_677), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_676), .B(n_678), .Y(n_692) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_681), .B(n_672), .Y(n_693) );
AOI211xp5_ASAP7_75t_SL g694 ( .A1(n_670), .A2(n_685), .B(n_683), .C(n_676), .Y(n_694) );
INVx2_ASAP7_75t_SL g695 ( .A(n_692), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_689), .B(n_682), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_691), .Y(n_697) );
INVx4_ASAP7_75t_L g698 ( .A(n_695), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_697), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_698), .Y(n_700) );
XOR2xp5_ASAP7_75t_L g701 ( .A(n_699), .B(n_696), .Y(n_701) );
BUFx2_ASAP7_75t_L g702 ( .A(n_700), .Y(n_702) );
BUFx2_ASAP7_75t_L g703 ( .A(n_701), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_702), .A2(n_694), .B1(n_690), .B2(n_693), .Y(n_704) );
OR2x6_ASAP7_75t_L g705 ( .A(n_704), .B(n_703), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g706 ( .A1(n_705), .A2(n_679), .B(n_686), .Y(n_706) );
O2A1O1Ixp33_ASAP7_75t_L g707 ( .A1(n_706), .A2(n_680), .B(n_675), .C(n_684), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_668), .B1(n_669), .B2(n_673), .Y(n_708) );
endmodule