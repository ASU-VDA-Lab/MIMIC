module fake_netlist_5_1952_n_2423 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_239, n_175, n_169, n_59, n_26, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2423);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_239;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2423;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2249;
wire n_2180;
wire n_344;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_1079;
wire n_457;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_2400;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_248;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_378;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2371;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2068;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_1178;
wire n_855;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1495;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_2414;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

INVx1_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_115),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_78),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_169),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_141),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_71),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_109),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_128),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_183),
.Y(n_251)
);

BUFx4f_ASAP7_75t_SL g252 ( 
.A(n_93),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_184),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_145),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_206),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_60),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_94),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_102),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_91),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_112),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_40),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_153),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_213),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_24),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_137),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_121),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_152),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_27),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_207),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_14),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_138),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_39),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_170),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_99),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_199),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_35),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_210),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_47),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_209),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_226),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_195),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_192),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_156),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_116),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_149),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_157),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_108),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_54),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_216),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_33),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_35),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_30),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_88),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_84),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_232),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_228),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_90),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_22),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_230),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_119),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_62),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_150),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_50),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_80),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_76),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_235),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_0),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_74),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_107),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_27),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_167),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_36),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_63),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_73),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_241),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_215),
.Y(n_317)
);

BUFx8_ASAP7_75t_SL g318 ( 
.A(n_239),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_161),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_64),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_72),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_102),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_45),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_155),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_11),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_238),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_56),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_189),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_129),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_172),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_134),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_171),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_66),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_68),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_163),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_179),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_85),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_136),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_200),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_100),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_52),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_66),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_78),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_12),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_237),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_234),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_113),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_23),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_188),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_40),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_131),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_132),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_89),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_236),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_180),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_160),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_24),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_182),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_164),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_117),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_178),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_190),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_77),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_65),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_47),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_12),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_181),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_74),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_101),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_73),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_48),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_82),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_61),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_97),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_57),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_22),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_34),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_114),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_29),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_1),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_45),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_49),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_81),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_205),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_62),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_214),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_69),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_146),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_202),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_108),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_14),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_186),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_112),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_223),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_140),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_53),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_176),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_56),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_82),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_75),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_233),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_71),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_130),
.Y(n_403)
);

BUFx5_ASAP7_75t_L g404 ( 
.A(n_75),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_158),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_10),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_7),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_217),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_127),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_218),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_64),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_69),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_42),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_173),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_103),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_77),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_4),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_109),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_7),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_8),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_201),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_148),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_10),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_2),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_80),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_220),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_194),
.Y(n_427)
);

INVxp33_ASAP7_75t_R g428 ( 
.A(n_191),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_104),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_147),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_123),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_84),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_198),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_106),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_31),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_97),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_53),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_48),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_94),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_177),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_83),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_185),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_0),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_79),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_174),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_52),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_23),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_90),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_219),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_212),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_89),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_68),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_19),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_229),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_13),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_8),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_41),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_154),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_107),
.Y(n_459)
);

CKINVDCx14_ASAP7_75t_R g460 ( 
.A(n_57),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_13),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_162),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_30),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_240),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_65),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_18),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_187),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_120),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_144),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_59),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_37),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_159),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_93),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_460),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_258),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_251),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_258),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_264),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_258),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_318),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_292),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_245),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_258),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_258),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_246),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_449),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_254),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_258),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_292),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_295),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_258),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_263),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_258),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_258),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_312),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_256),
.B(n_2),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_266),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_267),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_295),
.Y(n_499)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_311),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_404),
.B(n_3),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_311),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_404),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_367),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_404),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_404),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_312),
.B(n_3),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_270),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_272),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_404),
.B(n_4),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_404),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_276),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_327),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_327),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_404),
.Y(n_515)
);

CKINVDCx14_ASAP7_75t_R g516 ( 
.A(n_401),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_350),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_278),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_350),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_401),
.B(n_5),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_280),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_321),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_256),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_404),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_404),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_281),
.Y(n_526)
);

BUFx2_ASAP7_75t_SL g527 ( 
.A(n_250),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_377),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_271),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_271),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_377),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_282),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_271),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_283),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_294),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_284),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_294),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_285),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_406),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_286),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_294),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_287),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_250),
.B(n_5),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_416),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_406),
.B(n_465),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_253),
.B(n_6),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_416),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_302),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_242),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_302),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_302),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_244),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_253),
.B(n_6),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_340),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_340),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_290),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_296),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_300),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_301),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_307),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_R g561 ( 
.A(n_316),
.B(n_118),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_247),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_340),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_328),
.B(n_9),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_317),
.Y(n_565)
);

INVxp33_ASAP7_75t_SL g566 ( 
.A(n_249),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_324),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_376),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_326),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_330),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_332),
.Y(n_571)
);

CKINVDCx14_ASAP7_75t_R g572 ( 
.A(n_314),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_335),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_261),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_376),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_L g576 ( 
.A(n_289),
.B(n_9),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_336),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_338),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_339),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_376),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_265),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_393),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_347),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_351),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_393),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_242),
.B(n_11),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_393),
.Y(n_587)
);

INVxp33_ASAP7_75t_L g588 ( 
.A(n_257),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_328),
.B(n_15),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_358),
.B(n_15),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_358),
.B(n_16),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_415),
.Y(n_592)
);

BUFx2_ASAP7_75t_SL g593 ( 
.A(n_289),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_355),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_415),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_361),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_415),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_423),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_423),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_423),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g601 ( 
.A(n_367),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_456),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_386),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_388),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_475),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_482),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_475),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_477),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_485),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_545),
.B(n_367),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_504),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_545),
.B(n_406),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_601),
.B(n_389),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_539),
.B(n_465),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_477),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_479),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_487),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_492),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_479),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_483),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_483),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_484),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_476),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_504),
.B(n_392),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_504),
.B(n_405),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_484),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_539),
.B(n_409),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_488),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_488),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_491),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_522),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_593),
.B(n_465),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_491),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_543),
.B(n_410),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_546),
.B(n_553),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_493),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_593),
.B(n_456),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_508),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_509),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_518),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_493),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_494),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_534),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_536),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_542),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_494),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_503),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_564),
.B(n_427),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_557),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_503),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_505),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_505),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_506),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_506),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_511),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_558),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_515),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_559),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_516),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_522),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_560),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_567),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_515),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_589),
.B(n_430),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_529),
.B(n_456),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_524),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_524),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_525),
.Y(n_669)
);

INVxp67_ASAP7_75t_SL g670 ( 
.A(n_523),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_569),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_590),
.B(n_431),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_525),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_478),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_529),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_591),
.B(n_433),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_570),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_527),
.B(n_320),
.Y(n_678)
);

NAND2x1p5_ASAP7_75t_L g679 ( 
.A(n_501),
.B(n_352),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_530),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_571),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_530),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_533),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_573),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_R g685 ( 
.A(n_572),
.B(n_440),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_533),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_501),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_510),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_535),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_579),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_510),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_528),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_496),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_535),
.B(n_352),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_583),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_584),
.Y(n_696)
);

OA21x2_ASAP7_75t_L g697 ( 
.A1(n_537),
.A2(n_259),
.B(n_257),
.Y(n_697)
);

XOR2xp5_ASAP7_75t_L g698 ( 
.A(n_531),
.B(n_260),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_537),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_541),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_R g701 ( 
.A(n_480),
.B(n_454),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_586),
.A2(n_354),
.B(n_352),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_594),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_635),
.B(n_566),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_607),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_611),
.B(n_255),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_615),
.Y(n_707)
);

INVx5_ASAP7_75t_L g708 ( 
.A(n_615),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_605),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_687),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_612),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_687),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_615),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_660),
.B(n_474),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_687),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_607),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_608),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_615),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_611),
.B(n_596),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_608),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_616),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_631),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_616),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_623),
.Y(n_724)
);

AND2x4_ASAP7_75t_L g725 ( 
.A(n_611),
.B(n_255),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_637),
.B(n_495),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_631),
.B(n_531),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_687),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_635),
.A2(n_489),
.B1(n_520),
.B2(n_507),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_613),
.B(n_604),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_611),
.B(n_527),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_661),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_611),
.B(n_474),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_621),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_615),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_661),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_685),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_605),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_687),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_621),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_622),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_637),
.B(n_541),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_615),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_637),
.B(n_548),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_660),
.B(n_544),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_687),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_613),
.B(n_497),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_612),
.B(n_262),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_688),
.B(n_486),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_605),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_612),
.Y(n_751)
);

BUFx4f_ASAP7_75t_L g752 ( 
.A(n_687),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_688),
.B(n_362),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_622),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_685),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_605),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_619),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_630),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_630),
.Y(n_759)
);

AND2x6_ASAP7_75t_L g760 ( 
.A(n_687),
.B(n_688),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_660),
.B(n_544),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_623),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_632),
.B(n_548),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_688),
.B(n_362),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_636),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_610),
.B(n_262),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_691),
.B(n_384),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_634),
.B(n_498),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_610),
.B(n_268),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_636),
.Y(n_770)
);

INVx4_ASAP7_75t_SL g771 ( 
.A(n_615),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_691),
.B(n_384),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_619),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_698),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_619),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_610),
.B(n_268),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_614),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_646),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_606),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_701),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_615),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_692),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_619),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_634),
.B(n_512),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_691),
.B(n_552),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_692),
.B(n_547),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_646),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_628),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_632),
.B(n_550),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_702),
.B(n_274),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_628),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_620),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_632),
.B(n_550),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_658),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_647),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_614),
.B(n_670),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_647),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_614),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_648),
.B(n_354),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_620),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_691),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_702),
.B(n_274),
.Y(n_802)
);

BUFx10_ASAP7_75t_L g803 ( 
.A(n_703),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_620),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_624),
.B(n_562),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_678),
.B(n_547),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_628),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_652),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_652),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_628),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_629),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_653),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_692),
.B(n_574),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_624),
.B(n_581),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_653),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_629),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_693),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_657),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_625),
.B(n_462),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_679),
.A2(n_490),
.B1(n_517),
.B2(n_513),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_648),
.B(n_521),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_665),
.B(n_526),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_697),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_620),
.Y(n_824)
);

INVx1_ASAP7_75t_SL g825 ( 
.A(n_698),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_679),
.A2(n_490),
.B1(n_517),
.B2(n_513),
.Y(n_826)
);

BUFx8_ASAP7_75t_SL g827 ( 
.A(n_674),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_657),
.Y(n_828)
);

NAND2x1p5_ASAP7_75t_L g829 ( 
.A(n_702),
.B(n_297),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_697),
.Y(n_830)
);

BUFx4f_ASAP7_75t_L g831 ( 
.A(n_679),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_625),
.B(n_665),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_672),
.B(n_532),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_670),
.B(n_551),
.Y(n_834)
);

AND2x2_ASAP7_75t_SL g835 ( 
.A(n_672),
.B(n_354),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_666),
.B(n_297),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_676),
.B(n_538),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_697),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_697),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_658),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_693),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_620),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_678),
.B(n_540),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_676),
.B(n_627),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_620),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_627),
.B(n_502),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_620),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_666),
.B(n_694),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_679),
.B(n_468),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_697),
.B(n_514),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_620),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_629),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_609),
.B(n_556),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_626),
.Y(n_854)
);

INVx5_ASAP7_75t_L g855 ( 
.A(n_626),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_626),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_658),
.B(n_472),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_666),
.B(n_551),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_658),
.B(n_394),
.Y(n_859)
);

AND2x6_ASAP7_75t_L g860 ( 
.A(n_658),
.B(n_395),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_694),
.B(n_303),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_667),
.B(n_403),
.Y(n_862)
);

NAND3xp33_ASAP7_75t_L g863 ( 
.A(n_617),
.B(n_499),
.C(n_481),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_697),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_694),
.B(n_303),
.Y(n_865)
);

AND2x2_ASAP7_75t_SL g866 ( 
.A(n_641),
.B(n_395),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_667),
.B(n_329),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_832),
.B(n_667),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_711),
.Y(n_869)
);

OAI21xp33_ASAP7_75t_L g870 ( 
.A1(n_704),
.A2(n_500),
.B(n_586),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_768),
.A2(n_577),
.B1(n_578),
.B2(n_565),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_831),
.A2(n_603),
.B1(n_638),
.B2(n_618),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_796),
.B(n_639),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_844),
.B(n_667),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_752),
.B(n_640),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_823),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_796),
.B(n_519),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_752),
.B(n_643),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_850),
.A2(n_764),
.B(n_767),
.C(n_753),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_823),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_801),
.B(n_667),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_752),
.B(n_644),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_838),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_827),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_726),
.B(n_645),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_831),
.B(n_649),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_711),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_838),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_801),
.B(n_626),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_730),
.B(n_656),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_848),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_839),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_839),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_710),
.B(n_626),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_728),
.B(n_626),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_863),
.B(n_806),
.C(n_784),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_821),
.B(n_659),
.Y(n_897)
);

INVxp67_ASAP7_75t_L g898 ( 
.A(n_722),
.Y(n_898)
);

INVx8_ASAP7_75t_L g899 ( 
.A(n_760),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_848),
.B(n_626),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_777),
.Y(n_901)
);

INVx4_ASAP7_75t_L g902 ( 
.A(n_712),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_822),
.A2(n_663),
.B1(n_671),
.B2(n_662),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_799),
.B(n_626),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_799),
.B(n_650),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_799),
.B(n_650),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_858),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_831),
.A2(n_681),
.B1(n_684),
.B2(n_677),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_835),
.B(n_650),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_830),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_858),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_835),
.B(n_650),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_835),
.B(n_650),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_712),
.B(n_690),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_833),
.B(n_695),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_790),
.A2(n_464),
.B1(n_395),
.B2(n_641),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_837),
.B(n_696),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_722),
.Y(n_918)
);

AO22x1_ASAP7_75t_L g919 ( 
.A1(n_747),
.A2(n_374),
.B1(n_402),
.B2(n_321),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_777),
.B(n_650),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_798),
.B(n_650),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_712),
.B(n_650),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_798),
.B(n_772),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_715),
.B(n_651),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_763),
.B(n_651),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_830),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_L g927 ( 
.A(n_729),
.B(n_549),
.C(n_496),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_715),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_726),
.B(n_588),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_751),
.A2(n_331),
.B1(n_345),
.B2(n_329),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_751),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_763),
.B(n_651),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_789),
.B(n_651),
.Y(n_933)
);

NAND2xp33_ASAP7_75t_L g934 ( 
.A(n_760),
.B(n_864),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_749),
.B(n_428),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_789),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_817),
.B(n_428),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_790),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_793),
.B(n_651),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_715),
.B(n_651),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_780),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_864),
.A2(n_633),
.B(n_629),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_SL g943 ( 
.A1(n_794),
.A2(n_464),
.B(n_345),
.C(n_346),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_727),
.B(n_698),
.Y(n_944)
);

BUFx4f_ASAP7_75t_SL g945 ( 
.A(n_724),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_793),
.B(n_651),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_742),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_817),
.B(n_674),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_850),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_742),
.B(n_651),
.Y(n_950)
);

AOI221xp5_ASAP7_75t_L g951 ( 
.A1(n_820),
.A2(n_826),
.B1(n_424),
.B2(n_436),
.C(n_402),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_744),
.B(n_654),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_744),
.B(n_654),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_760),
.B(n_654),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_785),
.A2(n_464),
.B1(n_346),
.B2(n_349),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_705),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_760),
.B(n_654),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_739),
.B(n_654),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_739),
.B(n_654),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_805),
.A2(n_814),
.B1(n_841),
.B2(n_760),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_760),
.B(n_654),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_760),
.B(n_654),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_790),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_746),
.B(n_655),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_834),
.B(n_523),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_705),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_716),
.B(n_655),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_716),
.B(n_655),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_841),
.B(n_252),
.Y(n_969)
);

NOR3xp33_ASAP7_75t_L g970 ( 
.A(n_745),
.B(n_461),
.C(n_424),
.Y(n_970)
);

AND2x4_ASAP7_75t_SL g971 ( 
.A(n_779),
.B(n_408),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_846),
.B(n_374),
.Y(n_972)
);

NOR3xp33_ASAP7_75t_SL g973 ( 
.A(n_732),
.B(n_273),
.C(n_269),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_717),
.B(n_655),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_790),
.A2(n_641),
.B1(n_664),
.B2(n_642),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_746),
.B(n_655),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_717),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_802),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_720),
.B(n_655),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_802),
.A2(n_576),
.B(n_277),
.C(n_298),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_732),
.B(n_701),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_846),
.B(n_436),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_720),
.B(n_721),
.Y(n_983)
);

AOI21x1_ASAP7_75t_L g984 ( 
.A1(n_857),
.A2(n_664),
.B(n_642),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_L g985 ( 
.A(n_843),
.B(n_576),
.C(n_279),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_721),
.B(n_655),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_727),
.B(n_372),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_813),
.B(n_275),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_723),
.B(n_655),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_748),
.B(n_331),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_723),
.B(n_642),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_734),
.Y(n_992)
);

AND2x2_ASAP7_75t_SL g993 ( 
.A(n_802),
.B(n_866),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_734),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_736),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_740),
.B(n_664),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_813),
.B(n_288),
.Y(n_997)
);

AND2x6_ASAP7_75t_SL g998 ( 
.A(n_853),
.B(n_259),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_740),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_741),
.B(n_668),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_741),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_754),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_754),
.B(n_668),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_802),
.A2(n_668),
.B1(n_669),
.B2(n_633),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_766),
.A2(n_356),
.B1(n_359),
.B2(n_349),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_840),
.A2(n_669),
.B(n_633),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_829),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_758),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_758),
.B(n_633),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_866),
.B(n_243),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_759),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_759),
.B(n_669),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_736),
.B(n_834),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_765),
.B(n_669),
.Y(n_1014)
);

AND2x6_ASAP7_75t_L g1015 ( 
.A(n_766),
.B(n_356),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_765),
.B(n_673),
.Y(n_1016)
);

OR2x6_ASAP7_75t_L g1017 ( 
.A(n_733),
.B(n_359),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_782),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_L g1019 ( 
.A(n_860),
.B(n_243),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_782),
.B(n_314),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_770),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_766),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_780),
.B(n_291),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_770),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_866),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_786),
.B(n_819),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_778),
.B(n_673),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_778),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_787),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_787),
.B(n_673),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_795),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_786),
.B(n_293),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_849),
.B(n_243),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_761),
.Y(n_1034)
);

BUFx8_ASAP7_75t_L g1035 ( 
.A(n_748),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_706),
.B(n_243),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_795),
.B(n_673),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_797),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_860),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_797),
.B(n_397),
.Y(n_1040)
);

AND2x6_ASAP7_75t_SL g1041 ( 
.A(n_762),
.B(n_277),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_891),
.B(n_748),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_888),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_1018),
.Y(n_1044)
);

INVxp67_ASAP7_75t_SL g1045 ( 
.A(n_888),
.Y(n_1045)
);

INVx5_ASAP7_75t_L g1046 ( 
.A(n_899),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_929),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_901),
.B(n_748),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_956),
.Y(n_1049)
);

NOR2x1_ASAP7_75t_L g1050 ( 
.A(n_908),
.B(n_719),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_1013),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_923),
.B(n_766),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_890),
.B(n_769),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_1026),
.B(n_873),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_901),
.B(n_769),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_888),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_885),
.B(n_737),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_R g1058 ( 
.A(n_884),
.B(n_737),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_956),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_877),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_874),
.B(n_769),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_1022),
.B(n_769),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_1022),
.B(n_776),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_877),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_966),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_931),
.B(n_776),
.Y(n_1066)
);

AND3x1_ASAP7_75t_SL g1067 ( 
.A(n_951),
.B(n_306),
.C(n_298),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_868),
.B(n_776),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_966),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_945),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_869),
.B(n_776),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_888),
.Y(n_1072)
);

INVx5_ASAP7_75t_L g1073 ( 
.A(n_899),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_L g1074 ( 
.A(n_875),
.B(n_714),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_992),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_992),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_993),
.B(n_779),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_994),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_972),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_994),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1001),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_993),
.A2(n_836),
.B1(n_865),
.B2(n_861),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_960),
.B(n_808),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_944),
.B(n_774),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_938),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1001),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_935),
.B(n_898),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1021),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_897),
.B(n_755),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_SL g1090 ( 
.A(n_1025),
.B(n_755),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_938),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_887),
.B(n_836),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_949),
.B(n_808),
.Y(n_1093)
);

AND3x2_ASAP7_75t_SL g1094 ( 
.A(n_919),
.B(n_304),
.C(n_299),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_938),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_938),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1021),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_SL g1098 ( 
.A(n_937),
.B(n_308),
.C(n_305),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_SL g1099 ( 
.A(n_948),
.B(n_310),
.C(n_309),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1028),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_949),
.A2(n_836),
.B1(n_865),
.B2(n_861),
.Y(n_1101)
);

BUFx8_ASAP7_75t_L g1102 ( 
.A(n_981),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_977),
.B(n_809),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_999),
.B(n_809),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1028),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_907),
.B(n_836),
.Y(n_1106)
);

INVxp67_ASAP7_75t_SL g1107 ( 
.A(n_883),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_963),
.B(n_812),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1002),
.B(n_812),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1038),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_965),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1008),
.B(n_815),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_911),
.B(n_947),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_935),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1025),
.A2(n_829),
.B1(n_815),
.B2(n_828),
.Y(n_1115)
);

INVx5_ASAP7_75t_L g1116 ( 
.A(n_899),
.Y(n_1116)
);

BUFx3_ASAP7_75t_L g1117 ( 
.A(n_1035),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_936),
.B(n_861),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1038),
.Y(n_1119)
);

OR2x6_ASAP7_75t_L g1120 ( 
.A(n_935),
.B(n_861),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1011),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1024),
.B(n_818),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1029),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_965),
.B(n_779),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1031),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_963),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_963),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_876),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_915),
.B(n_779),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_963),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_983),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_896),
.A2(n_865),
.B1(n_818),
.B2(n_828),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_876),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_880),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_884),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_978),
.B(n_865),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_978),
.Y(n_1137)
);

OR2x2_ASAP7_75t_SL g1138 ( 
.A(n_927),
.B(n_825),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_880),
.B(n_862),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_978),
.Y(n_1140)
);

CKINVDCx16_ASAP7_75t_R g1141 ( 
.A(n_871),
.Y(n_1141)
);

OR2x6_ASAP7_75t_L g1142 ( 
.A(n_935),
.B(n_829),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_R g1143 ( 
.A(n_941),
.B(n_803),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_918),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_892),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_SL g1146 ( 
.A(n_917),
.B(n_344),
.C(n_342),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_892),
.Y(n_1147)
);

NOR3xp33_ASAP7_75t_SL g1148 ( 
.A(n_870),
.B(n_315),
.C(n_313),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_982),
.B(n_803),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_893),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_893),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_883),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1034),
.B(n_803),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_883),
.B(n_859),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_995),
.B(n_706),
.Y(n_1155)
);

BUFx12f_ASAP7_75t_L g1156 ( 
.A(n_1041),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_910),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_1020),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1025),
.B(n_706),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_910),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_987),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_926),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1025),
.B(n_706),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_926),
.B(n_725),
.Y(n_1164)
);

AND2x6_ASAP7_75t_SL g1165 ( 
.A(n_1023),
.B(n_988),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_899),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_879),
.B(n_900),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_950),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_902),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_990),
.B(n_725),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_990),
.B(n_725),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_991),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_990),
.B(n_725),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1017),
.A2(n_731),
.B1(n_860),
.B2(n_803),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_R g1175 ( 
.A(n_941),
.B(n_379),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_997),
.B(n_314),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_R g1177 ( 
.A(n_934),
.B(n_396),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_SL g1178 ( 
.A(n_985),
.B(n_333),
.C(n_323),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_952),
.B(n_713),
.Y(n_1179)
);

BUFx2_ASAP7_75t_L g1180 ( 
.A(n_1035),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_953),
.B(n_713),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_872),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_925),
.B(n_713),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1035),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_996),
.Y(n_1185)
);

AND2x6_ASAP7_75t_L g1186 ( 
.A(n_1007),
.B(n_743),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_902),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1017),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_902),
.B(n_743),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_932),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1000),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1003),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_967),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_968),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_933),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_974),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_979),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1010),
.A2(n_860),
.B1(n_322),
.B2(n_325),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1017),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_SL g1200 ( 
.A(n_886),
.B(n_418),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_986),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1032),
.B(n_314),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1017),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_939),
.B(n_743),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_886),
.B(n_438),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_SL g1206 ( 
.A(n_970),
.B(n_451),
.C(n_447),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_946),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_928),
.B(n_804),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_989),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_928),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1010),
.A2(n_860),
.B1(n_322),
.B2(n_325),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_928),
.B(n_804),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_903),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1009),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1012),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_971),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1039),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1015),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1014),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_971),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_914),
.B(n_397),
.Y(n_1221)
);

OR2x6_ASAP7_75t_L g1222 ( 
.A(n_914),
.B(n_875),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_969),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_916),
.B(n_920),
.Y(n_1224)
);

NOR2xp67_ASAP7_75t_L g1225 ( 
.A(n_878),
.B(n_882),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_921),
.B(n_804),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_878),
.B(n_414),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1016),
.Y(n_1228)
);

AND2x4_ASAP7_75t_L g1229 ( 
.A(n_882),
.B(n_414),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_973),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1039),
.B(n_847),
.Y(n_1231)
);

OR2x2_ASAP7_75t_SL g1232 ( 
.A(n_998),
.B(n_306),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1015),
.Y(n_1233)
);

NOR3xp33_ASAP7_75t_SL g1234 ( 
.A(n_955),
.B(n_337),
.C(n_334),
.Y(n_1234)
);

HB1xp67_ASAP7_75t_L g1235 ( 
.A(n_1040),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1007),
.B(n_847),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1131),
.B(n_1007),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1167),
.A2(n_905),
.B(n_904),
.Y(n_1238)
);

AOI22x1_ASAP7_75t_L g1239 ( 
.A1(n_1215),
.A2(n_1006),
.B1(n_942),
.B2(n_1033),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1157),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1049),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1224),
.A2(n_909),
.B(n_906),
.Y(n_1242)
);

AO21x2_ASAP7_75t_L g1243 ( 
.A1(n_1083),
.A2(n_1033),
.B(n_913),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_1046),
.B(n_1039),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1115),
.A2(n_984),
.B(n_889),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1049),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1044),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_1054),
.B(n_930),
.C(n_1005),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1226),
.A2(n_957),
.B(n_954),
.Y(n_1249)
);

NAND2x1_ASAP7_75t_L g1250 ( 
.A(n_1169),
.B(n_860),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1054),
.B(n_1015),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_SL g1252 ( 
.A1(n_1233),
.A2(n_912),
.B(n_867),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1061),
.A2(n_881),
.B(n_975),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1106),
.B(n_1015),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1069),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1043),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1069),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1053),
.B(n_1039),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1068),
.A2(n_895),
.B(n_894),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1111),
.B(n_980),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1129),
.A2(n_980),
.B(n_1019),
.C(n_407),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1236),
.A2(n_962),
.B(n_961),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1179),
.A2(n_924),
.B(n_922),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1181),
.A2(n_924),
.B(n_922),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1183),
.A2(n_958),
.B(n_940),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1051),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1076),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1084),
.B(n_1027),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1060),
.B(n_1030),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1204),
.A2(n_958),
.B(n_940),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1043),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1079),
.B(n_1015),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1108),
.A2(n_1152),
.B(n_1189),
.Y(n_1273)
);

BUFx10_ASAP7_75t_L g1274 ( 
.A(n_1057),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1080),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1124),
.B(n_1015),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1089),
.B(n_1037),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1108),
.A2(n_964),
.B(n_959),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1233),
.A2(n_1004),
.B(n_422),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1152),
.A2(n_964),
.B(n_959),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1070),
.Y(n_1281)
);

INVxp67_ASAP7_75t_SL g1282 ( 
.A(n_1043),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1089),
.B(n_976),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1080),
.A2(n_1081),
.A3(n_1086),
.B(n_1168),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1169),
.A2(n_1039),
.B(n_976),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1081),
.A2(n_738),
.A3(n_750),
.B(n_709),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_SL g1287 ( 
.A1(n_1082),
.A2(n_422),
.B(n_421),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1187),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1152),
.A2(n_1036),
.B(n_856),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1187),
.A2(n_1019),
.B(n_792),
.Y(n_1290)
);

OAI21xp33_ASAP7_75t_L g1291 ( 
.A1(n_1176),
.A2(n_353),
.B(n_348),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1205),
.A2(n_1146),
.B(n_1206),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_SL g1293 ( 
.A1(n_1166),
.A2(n_1036),
.B(n_718),
.Y(n_1293)
);

AOI221x1_ASAP7_75t_L g1294 ( 
.A1(n_1200),
.A2(n_469),
.B1(n_458),
.B2(n_450),
.C(n_445),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1189),
.A2(n_856),
.B(n_847),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1187),
.A2(n_792),
.B(n_781),
.Y(n_1296)
);

O2A1O1Ixp5_ASAP7_75t_L g1297 ( 
.A1(n_1129),
.A2(n_943),
.B(n_442),
.C(n_445),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1208),
.A2(n_856),
.B(n_738),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1208),
.A2(n_750),
.B(n_709),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1162),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1235),
.B(n_756),
.Y(n_1301)
);

AO21x1_ASAP7_75t_L g1302 ( 
.A1(n_1221),
.A2(n_442),
.B(n_421),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1223),
.B(n_357),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1212),
.A2(n_757),
.B(n_756),
.Y(n_1304)
);

OAI22x1_ASAP7_75t_L g1305 ( 
.A1(n_1205),
.A2(n_407),
.B1(n_372),
.B2(n_343),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1177),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1102),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1159),
.A2(n_458),
.B1(n_469),
.B2(n_450),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1164),
.A2(n_773),
.B(n_757),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1172),
.B(n_773),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1052),
.A2(n_783),
.B(n_775),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1102),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1064),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1210),
.A2(n_792),
.B(n_781),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1212),
.A2(n_783),
.B(n_775),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_SL g1316 ( 
.A(n_1135),
.B(n_408),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1168),
.A2(n_1195),
.B(n_1190),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1210),
.A2(n_845),
.B(n_781),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1190),
.A2(n_791),
.B(n_788),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1210),
.A2(n_845),
.B(n_718),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1106),
.B(n_771),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1154),
.A2(n_791),
.B(n_788),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1086),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1195),
.A2(n_810),
.B(n_807),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1193),
.A2(n_807),
.A3(n_810),
.B(n_852),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1163),
.A2(n_845),
.B(n_718),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1162),
.A2(n_1133),
.B(n_1128),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_SL g1328 ( 
.A(n_1135),
.B(n_408),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1128),
.A2(n_816),
.B(n_811),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1139),
.A2(n_816),
.B(n_811),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1185),
.B(n_852),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1133),
.A2(n_555),
.B(n_554),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_SL g1333 ( 
.A1(n_1207),
.A2(n_343),
.B(n_341),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1134),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1134),
.A2(n_555),
.B(n_554),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1143),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1046),
.A2(n_718),
.B(n_707),
.Y(n_1337)
);

BUFx4f_ASAP7_75t_L g1338 ( 
.A(n_1096),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_1153),
.B(n_122),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1102),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1059),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1147),
.A2(n_568),
.B(n_563),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1101),
.A2(n_800),
.B1(n_707),
.B2(n_718),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1191),
.B(n_860),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1106),
.B(n_771),
.Y(n_1345)
);

NAND2xp33_ASAP7_75t_L g1346 ( 
.A(n_1166),
.B(n_707),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1065),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1101),
.A2(n_800),
.B1(n_707),
.B2(n_854),
.Y(n_1348)
);

NOR4xp25_ASAP7_75t_L g1349 ( 
.A(n_1202),
.B(n_1149),
.C(n_1077),
.D(n_1094),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1075),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1200),
.A2(n_735),
.B1(n_707),
.B2(n_854),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1147),
.A2(n_568),
.B(n_563),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1207),
.A2(n_943),
.B(n_682),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1192),
.B(n_675),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1066),
.A2(n_682),
.B(n_675),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1078),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1151),
.A2(n_580),
.B(n_575),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1046),
.A2(n_800),
.B(n_735),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_SL g1359 ( 
.A1(n_1085),
.A2(n_363),
.B(n_341),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1118),
.B(n_771),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1194),
.A2(n_369),
.A3(n_370),
.B(n_371),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1151),
.A2(n_1050),
.B(n_1088),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1097),
.Y(n_1363)
);

AOI221x1_ASAP7_75t_L g1364 ( 
.A1(n_1221),
.A2(n_448),
.B1(n_363),
.B2(n_369),
.C(n_370),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1046),
.A2(n_800),
.B(n_735),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1100),
.A2(n_580),
.B(n_575),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1073),
.A2(n_800),
.B(n_735),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1105),
.A2(n_1119),
.B(n_1110),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1225),
.B(n_735),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1073),
.A2(n_842),
.B(n_824),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1160),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1145),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1073),
.A2(n_842),
.B(n_824),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1214),
.A2(n_686),
.B(n_683),
.Y(n_1374)
);

O2A1O1Ixp5_ASAP7_75t_L g1375 ( 
.A1(n_1221),
.A2(n_683),
.B(n_686),
.C(n_689),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1073),
.A2(n_842),
.B(n_824),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_SL g1377 ( 
.A1(n_1227),
.A2(n_561),
.B(n_426),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1121),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1057),
.B(n_365),
.C(n_364),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1196),
.A2(n_585),
.B(n_582),
.Y(n_1380)
);

OAI22x1_ASAP7_75t_L g1381 ( 
.A1(n_1213),
.A2(n_1188),
.B1(n_1203),
.B2(n_1199),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1116),
.A2(n_842),
.B(n_824),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1123),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1219),
.B(n_689),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1228),
.B(n_699),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1197),
.A2(n_1209),
.B(n_1201),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1125),
.Y(n_1387)
);

AOI221x1_ASAP7_75t_L g1388 ( 
.A1(n_1227),
.A2(n_463),
.B1(n_457),
.B2(n_448),
.C(n_444),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1113),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1231),
.A2(n_1173),
.B(n_1171),
.Y(n_1390)
);

NAND2xp33_ASAP7_75t_L g1391 ( 
.A(n_1166),
.B(n_824),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1113),
.B(n_699),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1132),
.A2(n_680),
.B(n_708),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1116),
.A2(n_851),
.B(n_842),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1047),
.B(n_582),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1150),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1215),
.A2(n_371),
.A3(n_387),
.B(n_391),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1137),
.A2(n_680),
.B(n_708),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1116),
.A2(n_854),
.B(n_851),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1140),
.A2(n_680),
.B(n_708),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1231),
.A2(n_587),
.B(n_585),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1144),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1103),
.A2(n_592),
.B(n_587),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1266),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1284),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1319),
.A2(n_1109),
.B(n_1104),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1292),
.B(n_1303),
.C(n_1098),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1402),
.B(n_1141),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1252),
.A2(n_1353),
.B(n_1362),
.Y(n_1409)
);

AO222x2_ASAP7_75t_L g1410 ( 
.A1(n_1395),
.A2(n_1094),
.B1(n_1113),
.B2(n_1227),
.C1(n_1229),
.C2(n_1232),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1274),
.B(n_1213),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1284),
.Y(n_1412)
);

NOR2x1_ASAP7_75t_SL g1413 ( 
.A(n_1369),
.B(n_1222),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1247),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1260),
.B(n_1118),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1319),
.A2(n_1122),
.B(n_1112),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1247),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1284),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1336),
.Y(n_1419)
);

OAI21xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1283),
.A2(n_1211),
.B(n_1198),
.Y(n_1420)
);

AO31x2_ASAP7_75t_L g1421 ( 
.A1(n_1302),
.A2(n_1093),
.A3(n_1153),
.B(n_1114),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1324),
.A2(n_1074),
.B(n_1077),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1260),
.B(n_1118),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1240),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1306),
.B(n_1138),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1324),
.A2(n_1126),
.B(n_1095),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1277),
.A2(n_1182),
.B1(n_1158),
.B2(n_1222),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1276),
.B(n_1042),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1248),
.A2(n_1182),
.B1(n_1177),
.B2(n_1229),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1240),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1266),
.Y(n_1431)
);

OAI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1316),
.A2(n_1161),
.B1(n_1087),
.B2(n_1099),
.C(n_1148),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1276),
.B(n_1042),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1306),
.A2(n_1229),
.B1(n_1389),
.B2(n_1042),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1254),
.B(n_1071),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1336),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1258),
.A2(n_1222),
.B(n_1055),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_SL g1438 ( 
.A1(n_1287),
.A2(n_1174),
.B(n_1091),
.Y(n_1438)
);

AOI22x1_ASAP7_75t_L g1439 ( 
.A1(n_1305),
.A2(n_1107),
.B1(n_1055),
.B2(n_1048),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1362),
.A2(n_1126),
.B(n_1095),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1300),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1329),
.A2(n_1126),
.B(n_1095),
.Y(n_1442)
);

AOI221xp5_ASAP7_75t_L g1443 ( 
.A1(n_1305),
.A2(n_1349),
.B1(n_1291),
.B2(n_1328),
.C(n_1381),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1281),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1300),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1395),
.B(n_1048),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1329),
.A2(n_1130),
.B(n_1198),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1268),
.B(n_1165),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1268),
.B(n_1142),
.Y(n_1449)
);

BUFx2_ASAP7_75t_SL g1450 ( 
.A(n_1281),
.Y(n_1450)
);

OAI211xp5_ASAP7_75t_L g1451 ( 
.A1(n_1294),
.A2(n_1175),
.B(n_1143),
.C(n_1230),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1317),
.A2(n_1130),
.B(n_1211),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1259),
.A2(n_1116),
.B(n_1217),
.Y(n_1453)
);

NAND2xp33_ASAP7_75t_SL g1454 ( 
.A(n_1381),
.B(n_1058),
.Y(n_1454)
);

AND2x6_ASAP7_75t_L g1455 ( 
.A(n_1288),
.B(n_1166),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1254),
.B(n_1071),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1334),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1334),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1241),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1317),
.A2(n_1130),
.B(n_1045),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1269),
.B(n_1155),
.Y(n_1461)
);

BUFx12f_ASAP7_75t_L g1462 ( 
.A(n_1307),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1269),
.B(n_1048),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1286),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1262),
.A2(n_595),
.B(n_592),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1372),
.B(n_1055),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1262),
.A2(n_597),
.B(n_595),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1327),
.A2(n_598),
.B(n_597),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1246),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1255),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1403),
.A2(n_599),
.B(n_598),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1245),
.A2(n_1178),
.B(n_1234),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1313),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1403),
.A2(n_600),
.B(n_599),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1327),
.A2(n_602),
.B(n_600),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1251),
.B(n_1142),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1238),
.A2(n_1217),
.B(n_1056),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1286),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1245),
.A2(n_1063),
.B(n_1062),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_SL g1480 ( 
.A1(n_1287),
.A2(n_1091),
.B(n_1085),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1379),
.A2(n_1230),
.B1(n_1090),
.B2(n_1087),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1307),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1286),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1354),
.B(n_1071),
.Y(n_1484)
);

BUFx2_ASAP7_75t_R g1485 ( 
.A(n_1312),
.Y(n_1485)
);

NAND3xp33_ASAP7_75t_L g1486 ( 
.A(n_1364),
.B(n_1142),
.C(n_1087),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1293),
.B(n_1043),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1295),
.A2(n_1380),
.B(n_1249),
.Y(n_1488)
);

OAI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1242),
.A2(n_1063),
.B(n_1062),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1254),
.B(n_1092),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1237),
.A2(n_1170),
.B1(n_1127),
.B2(n_1096),
.Y(n_1491)
);

AO32x2_ASAP7_75t_L g1492 ( 
.A1(n_1308),
.A2(n_1067),
.A3(n_1220),
.B1(n_1090),
.B2(n_1120),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1295),
.A2(n_602),
.B(n_1184),
.Y(n_1493)
);

BUFx12f_ASAP7_75t_L g1494 ( 
.A(n_1312),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1338),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1380),
.A2(n_680),
.B(n_1186),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1378),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1286),
.Y(n_1498)
);

AOI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1258),
.A2(n_1063),
.B(n_1062),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1274),
.A2(n_1216),
.B1(n_1120),
.B2(n_1092),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1288),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1257),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1372),
.B(n_1092),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1272),
.A2(n_1136),
.B1(n_1170),
.B2(n_1120),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1384),
.B(n_1136),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1338),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1340),
.A2(n_1175),
.B1(n_1117),
.B2(n_1180),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1267),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1275),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1321),
.Y(n_1510)
);

AO31x2_ASAP7_75t_L g1511 ( 
.A1(n_1302),
.A2(n_463),
.A3(n_391),
.B(n_400),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1274),
.B(n_1383),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1321),
.B(n_1136),
.Y(n_1513)
);

AO21x2_ASAP7_75t_L g1514 ( 
.A1(n_1261),
.A2(n_1170),
.B(n_400),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1340),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1323),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1387),
.Y(n_1517)
);

AO32x2_ASAP7_75t_L g1518 ( 
.A1(n_1343),
.A2(n_1067),
.A3(n_1186),
.B1(n_1218),
.B2(n_1056),
.Y(n_1518)
);

INVx2_ASAP7_75t_SL g1519 ( 
.A(n_1338),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1321),
.Y(n_1520)
);

NAND2x1_ASAP7_75t_L g1521 ( 
.A(n_1293),
.B(n_1186),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1385),
.B(n_1056),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1401),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1339),
.A2(n_1117),
.B1(n_1156),
.B2(n_1218),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1286),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1366),
.A2(n_420),
.B(n_387),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1301),
.B(n_1056),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1345),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1256),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1392),
.B(n_1072),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1401),
.Y(n_1531)
);

AOI222xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1333),
.A2(n_420),
.B1(n_457),
.B2(n_444),
.C1(n_441),
.C2(n_435),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1249),
.A2(n_1186),
.B(n_435),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1261),
.A2(n_1253),
.B1(n_1374),
.B2(n_1355),
.C(n_1344),
.Y(n_1534)
);

INVx4_ASAP7_75t_L g1535 ( 
.A(n_1256),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1366),
.A2(n_441),
.B(n_432),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1332),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1345),
.B(n_1058),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1332),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1256),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1273),
.A2(n_1186),
.B(n_432),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1390),
.A2(n_1386),
.B(n_1264),
.Y(n_1542)
);

AOI21xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1341),
.A2(n_368),
.B(n_366),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1390),
.A2(n_375),
.B(n_373),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1347),
.A2(n_1127),
.B1(n_1096),
.B2(n_1072),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1335),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1350),
.B(n_1356),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1282),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_SL g1549 ( 
.A1(n_1333),
.A2(n_1127),
.B(n_1096),
.Y(n_1549)
);

OAI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1388),
.A2(n_1156),
.B1(n_1127),
.B2(n_1072),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1335),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1273),
.A2(n_1072),
.B(n_1217),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1396),
.B(n_380),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1363),
.B(n_381),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1396),
.B(n_382),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_L g1556 ( 
.A(n_1375),
.B(n_434),
.C(n_383),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1371),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1393),
.A2(n_771),
.B(n_1217),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1386),
.B(n_1345),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1310),
.B(n_385),
.Y(n_1560)
);

AOI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1369),
.A2(n_854),
.B(n_851),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1398),
.A2(n_851),
.B(n_854),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1256),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1289),
.A2(n_1352),
.B(n_1342),
.Y(n_1564)
);

OAI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1263),
.A2(n_429),
.B(n_390),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1289),
.A2(n_851),
.B(n_855),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1342),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1360),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1331),
.B(n_398),
.Y(n_1569)
);

AO31x2_ASAP7_75t_L g1570 ( 
.A1(n_1348),
.A2(n_16),
.A3(n_17),
.B(n_18),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1360),
.B(n_124),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1352),
.A2(n_708),
.B(n_855),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1297),
.A2(n_437),
.B(n_399),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1357),
.A2(n_708),
.B(n_855),
.Y(n_1574)
);

INVx8_ASAP7_75t_L g1575 ( 
.A(n_1360),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1263),
.A2(n_453),
.B(n_413),
.Y(n_1576)
);

OAI21xp33_ASAP7_75t_L g1577 ( 
.A1(n_1351),
.A2(n_443),
.B(n_473),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1271),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1243),
.B(n_411),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1359),
.A2(n_471),
.B(n_470),
.C(n_466),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_SL g1581 ( 
.A1(n_1279),
.A2(n_231),
.B(n_227),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1346),
.A2(n_855),
.B(n_708),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1400),
.A2(n_243),
.B(n_248),
.Y(n_1583)
);

CKINVDCx11_ASAP7_75t_R g1584 ( 
.A(n_1271),
.Y(n_1584)
);

INVx4_ASAP7_75t_SL g1585 ( 
.A(n_1455),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_1419),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1429),
.A2(n_1239),
.B1(n_1243),
.B2(n_408),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1407),
.A2(n_1243),
.B1(n_426),
.B2(n_417),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1424),
.Y(n_1589)
);

AO21x2_ASAP7_75t_L g1590 ( 
.A1(n_1542),
.A2(n_1311),
.B(n_1309),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1420),
.A2(n_1544),
.B(n_1556),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1513),
.B(n_1271),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1584),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1436),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1547),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1459),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1415),
.B(n_1361),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1424),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1427),
.A2(n_459),
.B1(n_455),
.B2(n_452),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1443),
.A2(n_426),
.B1(n_446),
.B2(n_439),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1461),
.B(n_1361),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_SL g1602 ( 
.A(n_1487),
.B(n_1271),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1449),
.B(n_1361),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1415),
.B(n_1361),
.Y(n_1604)
);

OR2x6_ASAP7_75t_L g1605 ( 
.A(n_1487),
.B(n_1368),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1446),
.B(n_1361),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1410),
.A2(n_426),
.B1(n_412),
.B2(n_419),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1417),
.Y(n_1608)
);

INVxp67_ASAP7_75t_L g1609 ( 
.A(n_1431),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1423),
.B(n_1446),
.Y(n_1610)
);

NAND2xp33_ASAP7_75t_SL g1611 ( 
.A(n_1521),
.B(n_1250),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1430),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1430),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1469),
.Y(n_1614)
);

NAND2xp33_ASAP7_75t_R g1615 ( 
.A(n_1411),
.B(n_1278),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1495),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1445),
.Y(n_1617)
);

AOI222xp33_ASAP7_75t_L g1618 ( 
.A1(n_1448),
.A2(n_425),
.B1(n_1408),
.B2(n_1423),
.C1(n_1517),
.C2(n_1554),
.Y(n_1618)
);

CKINVDCx11_ASAP7_75t_R g1619 ( 
.A(n_1462),
.Y(n_1619)
);

NAND3xp33_ASAP7_75t_SL g1620 ( 
.A(n_1532),
.B(n_1330),
.C(n_1377),
.Y(n_1620)
);

OR2x6_ASAP7_75t_L g1621 ( 
.A(n_1487),
.B(n_1368),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1449),
.B(n_1397),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1445),
.Y(n_1623)
);

O2A1O1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1432),
.A2(n_1346),
.B(n_1391),
.C(n_1322),
.Y(n_1624)
);

OAI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1425),
.A2(n_243),
.B1(n_248),
.B2(n_319),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_SL g1626 ( 
.A(n_1451),
.B(n_1399),
.C(n_1337),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1534),
.A2(n_1391),
.B(n_1290),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1463),
.B(n_1397),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1458),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1414),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1425),
.B(n_1280),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1521),
.A2(n_1285),
.B(n_1320),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1470),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1560),
.B(n_1397),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1575),
.Y(n_1635)
);

CKINVDCx10_ASAP7_75t_R g1636 ( 
.A(n_1485),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1486),
.A2(n_1439),
.B1(n_1577),
.B2(n_1454),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1458),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_SL g1639 ( 
.A(n_1481),
.B(n_1326),
.C(n_1394),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1569),
.B(n_1397),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1557),
.B(n_1397),
.Y(n_1641)
);

AO21x2_ASAP7_75t_L g1642 ( 
.A1(n_1438),
.A2(n_1357),
.B(n_1264),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1512),
.A2(n_1244),
.B1(n_1376),
.B2(n_1373),
.Y(n_1643)
);

AO31x2_ASAP7_75t_L g1644 ( 
.A1(n_1464),
.A2(n_1483),
.A3(n_1498),
.B(n_1478),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_1436),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_SL g1646 ( 
.A1(n_1439),
.A2(n_1450),
.B1(n_1497),
.B2(n_1413),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_SL g1647 ( 
.A(n_1550),
.B(n_1489),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1484),
.A2(n_248),
.B1(n_319),
.B2(n_360),
.Y(n_1648)
);

OAI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1507),
.A2(n_1296),
.B1(n_1314),
.B2(n_1318),
.C(n_378),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1503),
.B(n_1325),
.Y(n_1650)
);

INVx3_ASAP7_75t_L g1651 ( 
.A(n_1495),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1434),
.A2(n_1382),
.B1(n_1370),
.B2(n_1367),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1419),
.Y(n_1653)
);

A2O1A1Ixp33_ASAP7_75t_L g1654 ( 
.A1(n_1571),
.A2(n_1265),
.B(n_1270),
.C(n_1278),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1495),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1428),
.B(n_1325),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1473),
.Y(n_1657)
);

AO21x2_ASAP7_75t_L g1658 ( 
.A1(n_1438),
.A2(n_1270),
.B(n_1265),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1500),
.A2(n_1280),
.B1(n_248),
.B2(n_360),
.Y(n_1659)
);

INVx3_ASAP7_75t_L g1660 ( 
.A(n_1575),
.Y(n_1660)
);

NOR2x1_ASAP7_75t_SL g1661 ( 
.A(n_1476),
.B(n_1325),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1505),
.A2(n_248),
.B1(n_319),
.B2(n_467),
.Y(n_1662)
);

OAI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1524),
.A2(n_1365),
.B1(n_1358),
.B2(n_248),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1565),
.A2(n_1315),
.B(n_1304),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1503),
.B(n_1325),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1428),
.A2(n_319),
.B1(n_360),
.B2(n_378),
.Y(n_1666)
);

AND2x6_ASAP7_75t_L g1667 ( 
.A(n_1559),
.B(n_319),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_SL g1668 ( 
.A(n_1580),
.B(n_17),
.C(n_19),
.Y(n_1668)
);

CKINVDCx8_ASAP7_75t_R g1669 ( 
.A(n_1450),
.Y(n_1669)
);

AOI222xp33_ASAP7_75t_L g1670 ( 
.A1(n_1404),
.A2(n_1433),
.B1(n_1576),
.B2(n_1494),
.C1(n_1462),
.C2(n_1538),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1502),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1513),
.B(n_1325),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1553),
.B(n_1315),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1433),
.B(n_319),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1502),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1435),
.A2(n_360),
.B1(n_378),
.B2(n_467),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1579),
.A2(n_467),
.B1(n_378),
.B2(n_360),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1441),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1513),
.B(n_1299),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1476),
.B(n_1298),
.Y(n_1680)
);

CKINVDCx6p67_ASAP7_75t_R g1681 ( 
.A(n_1494),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1575),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1579),
.A2(n_467),
.B1(n_378),
.B2(n_360),
.Y(n_1683)
);

AOI221x1_ASAP7_75t_L g1684 ( 
.A1(n_1581),
.A2(n_467),
.B1(n_378),
.B2(n_700),
.C(n_1298),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1504),
.A2(n_467),
.B1(n_855),
.B2(n_700),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1466),
.B(n_20),
.Y(n_1686)
);

OAI21x1_ASAP7_75t_L g1687 ( 
.A1(n_1468),
.A2(n_1304),
.B(n_1299),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1466),
.B(n_20),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1508),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1553),
.B(n_21),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1514),
.A2(n_700),
.B1(n_25),
.B2(n_26),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_SL g1692 ( 
.A1(n_1413),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1555),
.B(n_28),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1453),
.A2(n_855),
.B(n_700),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1543),
.B(n_700),
.C(n_29),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1477),
.A2(n_700),
.B(n_225),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1514),
.A2(n_700),
.B1(n_31),
.B2(n_32),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1514),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1508),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1571),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_1700)
);

AOI222xp33_ASAP7_75t_L g1701 ( 
.A1(n_1414),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.C1(n_38),
.C2(n_39),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1435),
.B(n_224),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1444),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1509),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1417),
.A2(n_700),
.B1(n_41),
.B2(n_42),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1457),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1435),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1472),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1472),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1457),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1472),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1482),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1555),
.A2(n_51),
.B1(n_55),
.B2(n_58),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1548),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1456),
.A2(n_1490),
.B1(n_1571),
.B2(n_1482),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1509),
.A2(n_61),
.B1(n_63),
.B2(n_67),
.Y(n_1716)
);

NAND2x1p5_ASAP7_75t_L g1717 ( 
.A(n_1548),
.B(n_222),
.Y(n_1717)
);

OAI21x1_ASAP7_75t_L g1718 ( 
.A1(n_1468),
.A2(n_221),
.B(n_208),
.Y(n_1718)
);

OR2x6_ASAP7_75t_L g1719 ( 
.A(n_1480),
.B(n_1559),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1456),
.B(n_67),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1529),
.A2(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_1721)
);

OAI221xp5_ASAP7_75t_L g1722 ( 
.A1(n_1543),
.A2(n_70),
.B1(n_79),
.B2(n_81),
.C(n_83),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_SL g1723 ( 
.A1(n_1583),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_1723)
);

AOI221xp5_ASAP7_75t_L g1724 ( 
.A1(n_1581),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.C(n_91),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_SL g1725 ( 
.A(n_1529),
.B(n_92),
.C(n_95),
.Y(n_1725)
);

AO221x2_ASAP7_75t_L g1726 ( 
.A1(n_1518),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.C(n_98),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1575),
.Y(n_1727)
);

INVx4_ASAP7_75t_L g1728 ( 
.A(n_1535),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1456),
.B(n_133),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1475),
.A2(n_135),
.B(n_203),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1510),
.B(n_96),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1516),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1522),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1422),
.A2(n_101),
.B(n_103),
.Y(n_1734)
);

OAI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1515),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_1735)
);

AO21x2_ASAP7_75t_L g1736 ( 
.A1(n_1480),
.A2(n_151),
.B(n_196),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1515),
.A2(n_105),
.B1(n_110),
.B2(n_111),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1490),
.A2(n_110),
.B1(n_111),
.B2(n_125),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1490),
.A2(n_126),
.B1(n_139),
.B2(n_142),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1558),
.A2(n_204),
.B(n_165),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1530),
.A2(n_143),
.B1(n_166),
.B2(n_168),
.C(n_175),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1510),
.B(n_193),
.Y(n_1742)
);

AOI21x1_ASAP7_75t_L g1743 ( 
.A1(n_1561),
.A2(n_1437),
.B(n_1499),
.Y(n_1743)
);

AO21x2_ASAP7_75t_L g1744 ( 
.A1(n_1465),
.A2(n_1467),
.B(n_1488),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1510),
.B(n_1520),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1558),
.A2(n_1583),
.B(n_1409),
.Y(n_1746)
);

OAI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1506),
.A2(n_1519),
.B1(n_1527),
.B2(n_1528),
.Y(n_1747)
);

AO31x2_ASAP7_75t_L g1748 ( 
.A1(n_1464),
.A2(n_1478),
.A3(n_1483),
.B(n_1498),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1520),
.B(n_1528),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1573),
.A2(n_1568),
.B1(n_1528),
.B2(n_1520),
.Y(n_1750)
);

AOI21xp33_ASAP7_75t_L g1751 ( 
.A1(n_1491),
.A2(n_1409),
.B(n_1573),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1568),
.B(n_1519),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1412),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1573),
.A2(n_1568),
.B1(n_1583),
.B2(n_1412),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1506),
.B(n_1421),
.Y(n_1755)
);

AO21x2_ASAP7_75t_L g1756 ( 
.A1(n_1465),
.A2(n_1467),
.B(n_1488),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1421),
.B(n_1501),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1573),
.A2(n_1405),
.B1(n_1418),
.B2(n_1409),
.Y(n_1758)
);

AOI21xp33_ASAP7_75t_L g1759 ( 
.A1(n_1479),
.A2(n_1545),
.B(n_1549),
.Y(n_1759)
);

NAND3xp33_ASAP7_75t_SL g1760 ( 
.A(n_1578),
.B(n_1535),
.C(n_1523),
.Y(n_1760)
);

AOI222xp33_ASAP7_75t_L g1761 ( 
.A1(n_1405),
.A2(n_1418),
.B1(n_1525),
.B2(n_1549),
.C1(n_1501),
.C2(n_1455),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1455),
.A2(n_1558),
.B1(n_1535),
.B2(n_1540),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1540),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1563),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1563),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1421),
.B(n_1437),
.Y(n_1766)
);

AND2x4_ASAP7_75t_L g1767 ( 
.A(n_1499),
.B(n_1455),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1523),
.A2(n_1531),
.B1(n_1536),
.B2(n_1526),
.C(n_1551),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1422),
.B(n_1406),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1570),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1479),
.A2(n_1525),
.B1(n_1416),
.B2(n_1406),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1518),
.A2(n_1570),
.B1(n_1492),
.B2(n_1567),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1607),
.A2(n_1531),
.B1(n_1567),
.B2(n_1551),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1610),
.B(n_1421),
.Y(n_1774)
);

OA21x2_ASAP7_75t_L g1775 ( 
.A1(n_1684),
.A2(n_1564),
.B(n_1533),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1607),
.A2(n_1479),
.B1(n_1416),
.B2(n_1562),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_SL g1777 ( 
.A1(n_1618),
.A2(n_1492),
.B1(n_1570),
.B2(n_1518),
.C(n_1421),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1597),
.B(n_1492),
.Y(n_1778)
);

OAI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1600),
.A2(n_1526),
.B1(n_1536),
.B2(n_1546),
.C(n_1539),
.Y(n_1779)
);

AO22x1_ASAP7_75t_L g1780 ( 
.A1(n_1593),
.A2(n_1455),
.B1(n_1570),
.B2(n_1492),
.Y(n_1780)
);

OAI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1707),
.A2(n_1518),
.B1(n_1492),
.B2(n_1570),
.Y(n_1781)
);

AO22x1_ASAP7_75t_L g1782 ( 
.A1(n_1593),
.A2(n_1455),
.B1(n_1537),
.B2(n_1546),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1603),
.B(n_1511),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1600),
.A2(n_1526),
.B1(n_1536),
.B2(n_1539),
.C(n_1537),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1630),
.B(n_1440),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1701),
.A2(n_1562),
.B1(n_1526),
.B2(n_1536),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1726),
.A2(n_1562),
.B1(n_1474),
.B2(n_1471),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1635),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1604),
.B(n_1511),
.Y(n_1789)
);

OAI211xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1599),
.A2(n_1511),
.B(n_1582),
.C(n_1518),
.Y(n_1790)
);

OAI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1735),
.A2(n_1474),
.B1(n_1471),
.B2(n_1561),
.Y(n_1791)
);

OAI222xp33_ASAP7_75t_L g1792 ( 
.A1(n_1700),
.A2(n_1511),
.B1(n_1440),
.B2(n_1452),
.C1(n_1460),
.C2(n_1541),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1726),
.A2(n_1474),
.B1(n_1471),
.B2(n_1452),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1591),
.A2(n_1471),
.B1(n_1474),
.B2(n_1511),
.C(n_1533),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1595),
.B(n_1460),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1657),
.B(n_1426),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1703),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1668),
.A2(n_1493),
.B(n_1541),
.Y(n_1798)
);

OAI22xp33_ASAP7_75t_SL g1799 ( 
.A1(n_1722),
.A2(n_1493),
.B1(n_1426),
.B2(n_1475),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1657),
.B(n_1609),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1700),
.A2(n_1552),
.B1(n_1442),
.B2(n_1447),
.Y(n_1801)
);

BUFx2_ASAP7_75t_L g1802 ( 
.A(n_1630),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1614),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1633),
.Y(n_1804)
);

OAI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1713),
.A2(n_1496),
.B1(n_1552),
.B2(n_1442),
.C(n_1447),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1726),
.A2(n_1564),
.B1(n_1496),
.B2(n_1566),
.Y(n_1806)
);

OAI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1735),
.A2(n_1566),
.B1(n_1574),
.B2(n_1572),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_SL g1808 ( 
.A1(n_1695),
.A2(n_1572),
.B1(n_1574),
.B2(n_1734),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1737),
.A2(n_1713),
.B1(n_1711),
.B2(n_1709),
.C(n_1708),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_SL g1810 ( 
.A1(n_1692),
.A2(n_1711),
.B1(n_1709),
.B2(n_1708),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1720),
.B(n_1674),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1637),
.A2(n_1666),
.B1(n_1715),
.B2(n_1669),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1737),
.A2(n_1733),
.B1(n_1716),
.B2(n_1724),
.C(n_1714),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1635),
.Y(n_1814)
);

OAI211xp5_ASAP7_75t_L g1815 ( 
.A1(n_1716),
.A2(n_1692),
.B(n_1738),
.C(n_1588),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1637),
.A2(n_1666),
.B1(n_1588),
.B2(n_1647),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1725),
.A2(n_1647),
.B1(n_1620),
.B2(n_1691),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1644),
.Y(n_1818)
);

OAI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1627),
.A2(n_1640),
.B(n_1634),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1656),
.B(n_1686),
.Y(n_1820)
);

AO222x2_ASAP7_75t_L g1821 ( 
.A1(n_1636),
.A2(n_1721),
.B1(n_1693),
.B2(n_1690),
.C1(n_1702),
.C2(n_1729),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1609),
.B(n_1688),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1691),
.A2(n_1697),
.B1(n_1723),
.B2(n_1625),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1601),
.B(n_1631),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1625),
.A2(n_1705),
.B1(n_1697),
.B2(n_1739),
.C(n_1772),
.Y(n_1825)
);

AOI22x1_ASAP7_75t_L g1826 ( 
.A1(n_1670),
.A2(n_1717),
.B1(n_1696),
.B2(n_1712),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1723),
.A2(n_1587),
.B1(n_1683),
.B2(n_1677),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1624),
.B(n_1646),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1587),
.A2(n_1677),
.B1(n_1683),
.B2(n_1648),
.Y(n_1829)
);

OAI21x1_ASAP7_75t_L g1830 ( 
.A1(n_1632),
.A2(n_1743),
.B(n_1687),
.Y(n_1830)
);

BUFx2_ASAP7_75t_L g1831 ( 
.A(n_1763),
.Y(n_1831)
);

OAI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1739),
.A2(n_1648),
.B1(n_1662),
.B2(n_1741),
.C(n_1676),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1765),
.Y(n_1833)
);

OR2x6_ASAP7_75t_SL g1834 ( 
.A(n_1594),
.B(n_1645),
.Y(n_1834)
);

AOI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1662),
.A2(n_1772),
.B1(n_1685),
.B2(n_1649),
.C(n_1770),
.Y(n_1835)
);

OAI211xp5_ASAP7_75t_L g1836 ( 
.A1(n_1731),
.A2(n_1659),
.B(n_1646),
.C(n_1606),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1671),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1622),
.A2(n_1639),
.B1(n_1593),
.B2(n_1619),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1675),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1593),
.A2(n_1619),
.B1(n_1702),
.B2(n_1729),
.Y(n_1840)
);

AOI221xp5_ASAP7_75t_L g1841 ( 
.A1(n_1751),
.A2(n_1663),
.B1(n_1641),
.B2(n_1628),
.C(n_1680),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1608),
.A2(n_1586),
.B1(n_1653),
.B2(n_1717),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_R g1843 ( 
.A(n_1615),
.B(n_1616),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1635),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1602),
.A2(n_1654),
.B(n_1643),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1673),
.A2(n_1681),
.B1(n_1672),
.B2(n_1704),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1655),
.A2(n_1616),
.B1(n_1651),
.B2(n_1727),
.Y(n_1847)
);

OAI211xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1755),
.A2(n_1750),
.B(n_1752),
.C(n_1759),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1745),
.B(n_1749),
.Y(n_1849)
);

INVx5_ASAP7_75t_SL g1850 ( 
.A(n_1635),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1682),
.Y(n_1851)
);

AOI221xp5_ASAP7_75t_L g1852 ( 
.A1(n_1680),
.A2(n_1747),
.B1(n_1766),
.B2(n_1750),
.C(n_1698),
.Y(n_1852)
);

OAI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1655),
.A2(n_1651),
.B1(n_1727),
.B2(n_1762),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1689),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1698),
.A2(n_1757),
.B1(n_1754),
.B2(n_1650),
.C(n_1665),
.Y(n_1855)
);

OAI211xp5_ASAP7_75t_L g1856 ( 
.A1(n_1754),
.A2(n_1740),
.B(n_1699),
.C(n_1732),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1589),
.B(n_1612),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1615),
.A2(n_1682),
.B1(n_1660),
.B2(n_1605),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1672),
.A2(n_1742),
.B1(n_1667),
.B2(n_1706),
.Y(n_1859)
);

AOI222xp33_ASAP7_75t_L g1860 ( 
.A1(n_1667),
.A2(n_1742),
.B1(n_1585),
.B2(n_1652),
.C1(n_1678),
.C2(n_1592),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1667),
.A2(n_1736),
.B1(n_1710),
.B2(n_1592),
.Y(n_1861)
);

OAI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1682),
.A2(n_1660),
.B1(n_1605),
.B2(n_1621),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1765),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1758),
.A2(n_1654),
.B1(n_1768),
.B2(n_1771),
.C(n_1760),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1667),
.A2(n_1736),
.B1(n_1679),
.B2(n_1598),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1667),
.A2(n_1679),
.B1(n_1613),
.B2(n_1617),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1626),
.A2(n_1719),
.B1(n_1605),
.B2(n_1621),
.Y(n_1867)
);

OAI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1626),
.A2(n_1664),
.B1(n_1611),
.B2(n_1621),
.C(n_1764),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1719),
.A2(n_1682),
.B1(n_1767),
.B2(n_1728),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_SL g1870 ( 
.A1(n_1767),
.A2(n_1661),
.B1(n_1730),
.B2(n_1718),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1638),
.A2(n_1590),
.B1(n_1623),
.B2(n_1629),
.Y(n_1871)
);

OAI211xp5_ASAP7_75t_L g1872 ( 
.A1(n_1758),
.A2(n_1771),
.B(n_1761),
.C(n_1746),
.Y(n_1872)
);

INVx4_ASAP7_75t_L g1873 ( 
.A(n_1728),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1623),
.B(n_1629),
.Y(n_1874)
);

CKINVDCx5p33_ASAP7_75t_R g1875 ( 
.A(n_1585),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_SL g1876 ( 
.A1(n_1753),
.A2(n_1585),
.B1(n_1611),
.B2(n_1658),
.Y(n_1876)
);

OAI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1769),
.A2(n_1694),
.B1(n_1642),
.B2(n_1590),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1644),
.Y(n_1878)
);

OAI21x1_ASAP7_75t_SL g1879 ( 
.A1(n_1644),
.A2(n_1748),
.B(n_1769),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1744),
.A2(n_1607),
.B1(n_1701),
.B2(n_1726),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1748),
.A2(n_1607),
.B1(n_1182),
.B2(n_1129),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1744),
.A2(n_1756),
.B(n_1748),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_SL g1883 ( 
.A1(n_1756),
.A2(n_1129),
.B1(n_890),
.B2(n_1726),
.Y(n_1883)
);

OAI21xp33_ASAP7_75t_L g1884 ( 
.A1(n_1748),
.A2(n_704),
.B(n_890),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1607),
.A2(n_1701),
.B1(n_1726),
.B2(n_1618),
.Y(n_1885)
);

AO22x2_ASAP7_75t_L g1886 ( 
.A1(n_1770),
.A2(n_1647),
.B1(n_1294),
.B2(n_1486),
.Y(n_1886)
);

OAI221xp5_ASAP7_75t_L g1887 ( 
.A1(n_1607),
.A2(n_890),
.B1(n_1292),
.B2(n_729),
.C(n_915),
.Y(n_1887)
);

OAI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1707),
.A2(n_1735),
.B1(n_1737),
.B2(n_1722),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1618),
.A2(n_890),
.B1(n_915),
.B2(n_897),
.Y(n_1889)
);

BUFx6f_ASAP7_75t_L g1890 ( 
.A(n_1635),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_1669),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1596),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_L g1893 ( 
.A1(n_1607),
.A2(n_1182),
.B1(n_1129),
.B2(n_1429),
.Y(n_1893)
);

OAI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1707),
.A2(n_1735),
.B1(n_1737),
.B2(n_1722),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_SL g1895 ( 
.A1(n_1726),
.A2(n_1129),
.B1(n_890),
.B2(n_1182),
.Y(n_1895)
);

OAI321xp33_ASAP7_75t_L g1896 ( 
.A1(n_1735),
.A2(n_1737),
.A3(n_1709),
.B1(n_1708),
.B2(n_1711),
.C(n_1722),
.Y(n_1896)
);

AO21x2_ASAP7_75t_L g1897 ( 
.A1(n_1591),
.A2(n_1751),
.B(n_1664),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1712),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1607),
.A2(n_1701),
.B1(n_1726),
.B2(n_1618),
.Y(n_1899)
);

O2A1O1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1668),
.A2(n_890),
.B(n_915),
.C(n_897),
.Y(n_1900)
);

AOI221xp5_ASAP7_75t_L g1901 ( 
.A1(n_1607),
.A2(n_729),
.B1(n_704),
.B2(n_919),
.C(n_870),
.Y(n_1901)
);

INVx5_ASAP7_75t_SL g1902 ( 
.A(n_1593),
.Y(n_1902)
);

AND2x2_ASAP7_75t_SL g1903 ( 
.A(n_1708),
.B(n_1129),
.Y(n_1903)
);

AOI31xp67_ASAP7_75t_L g1904 ( 
.A1(n_1768),
.A2(n_1649),
.A3(n_1534),
.B(n_1659),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1607),
.A2(n_1701),
.B1(n_1726),
.B2(n_1618),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1595),
.B(n_1054),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1607),
.A2(n_1182),
.B1(n_1129),
.B2(n_1429),
.Y(n_1907)
);

OAI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1607),
.A2(n_890),
.B1(n_1292),
.B2(n_729),
.C(n_915),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1607),
.A2(n_1182),
.B1(n_1129),
.B2(n_1429),
.Y(n_1909)
);

AOI221xp5_ASAP7_75t_L g1910 ( 
.A1(n_1607),
.A2(n_729),
.B1(n_704),
.B2(n_919),
.C(n_870),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1635),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1596),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_SL g1913 ( 
.A1(n_1726),
.A2(n_1129),
.B1(n_890),
.B2(n_1182),
.Y(n_1913)
);

AOI21xp33_ASAP7_75t_L g1914 ( 
.A1(n_1591),
.A2(n_890),
.B(n_1129),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1603),
.B(n_1622),
.Y(n_1915)
);

OAI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1707),
.A2(n_1735),
.B1(n_1737),
.B2(n_1722),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1607),
.A2(n_729),
.B1(n_704),
.B2(n_919),
.C(n_870),
.Y(n_1917)
);

OAI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1707),
.A2(n_1735),
.B1(n_1737),
.B2(n_1722),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1607),
.A2(n_729),
.B1(n_704),
.B2(n_919),
.C(n_870),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1595),
.B(n_1054),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1607),
.A2(n_1701),
.B1(n_1726),
.B2(n_1618),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1603),
.B(n_1622),
.Y(n_1922)
);

AOI221xp5_ASAP7_75t_L g1923 ( 
.A1(n_1607),
.A2(n_729),
.B1(n_704),
.B2(n_919),
.C(n_870),
.Y(n_1923)
);

OAI211xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1618),
.A2(n_729),
.B(n_1607),
.C(n_1292),
.Y(n_1924)
);

AOI21xp33_ASAP7_75t_L g1925 ( 
.A1(n_1591),
.A2(n_890),
.B(n_1129),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1607),
.A2(n_1701),
.B1(n_1726),
.B2(n_1618),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1607),
.A2(n_1701),
.B1(n_1726),
.B2(n_1618),
.Y(n_1927)
);

OAI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1607),
.A2(n_1182),
.B1(n_1129),
.B2(n_1429),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1595),
.B(n_1054),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1627),
.A2(n_831),
.B(n_1129),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1596),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1607),
.A2(n_1182),
.B1(n_1129),
.B2(n_1429),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1603),
.B(n_1622),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1607),
.A2(n_1701),
.B1(n_1726),
.B2(n_1618),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1596),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1778),
.B(n_1789),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1824),
.B(n_1819),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1774),
.B(n_1878),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1897),
.B(n_1818),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1879),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1915),
.B(n_1922),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1900),
.A2(n_1889),
.B(n_1914),
.Y(n_1942)
);

INVx4_ASAP7_75t_L g1943 ( 
.A(n_1875),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1933),
.B(n_1783),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1803),
.B(n_1804),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1785),
.Y(n_1946)
);

OAI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1887),
.A2(n_1908),
.B1(n_1896),
.B2(n_1809),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1837),
.B(n_1839),
.Y(n_1948)
);

HB1xp67_ASAP7_75t_L g1949 ( 
.A(n_1796),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1793),
.B(n_1852),
.Y(n_1950)
);

INVx3_ASAP7_75t_L g1951 ( 
.A(n_1785),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1854),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1935),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1892),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1871),
.B(n_1780),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1912),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1931),
.B(n_1849),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1795),
.Y(n_1958)
);

OAI21xp5_ASAP7_75t_L g1959 ( 
.A1(n_1925),
.A2(n_1816),
.B(n_1903),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1849),
.B(n_1906),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1830),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1920),
.B(n_1929),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1855),
.B(n_1820),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1775),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1877),
.B(n_1882),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1871),
.B(n_1806),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1841),
.B(n_1883),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1806),
.B(n_1864),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1787),
.B(n_1886),
.Y(n_1969)
);

OA21x2_ASAP7_75t_L g1970 ( 
.A1(n_1787),
.A2(n_1792),
.B(n_1798),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1867),
.B(n_1872),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1886),
.B(n_1874),
.Y(n_1972)
);

CKINVDCx5p33_ASAP7_75t_R g1973 ( 
.A(n_1834),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1924),
.A2(n_1934),
.B1(n_1885),
.B2(n_1905),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1886),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1876),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1885),
.A2(n_1934),
.B1(n_1899),
.B2(n_1905),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1843),
.B(n_1845),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1775),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1775),
.Y(n_1980)
);

HB1xp67_ASAP7_75t_L g1981 ( 
.A(n_1843),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1828),
.B(n_1865),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1857),
.Y(n_1983)
);

INVxp67_ASAP7_75t_SL g1984 ( 
.A(n_1791),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1848),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1899),
.A2(n_1921),
.B1(n_1926),
.B2(n_1927),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1862),
.Y(n_1987)
);

HB1xp67_ASAP7_75t_L g1988 ( 
.A(n_1802),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1828),
.B(n_1865),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1794),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1861),
.B(n_1838),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1862),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1861),
.B(n_1838),
.Y(n_1993)
);

INVxp67_ASAP7_75t_L g1994 ( 
.A(n_1833),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1781),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1781),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1868),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1777),
.B(n_1858),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1846),
.B(n_1895),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1846),
.B(n_1913),
.Y(n_2000)
);

BUFx2_ASAP7_75t_L g2001 ( 
.A(n_1858),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1870),
.B(n_1776),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1776),
.B(n_1811),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1866),
.B(n_1808),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1866),
.B(n_1860),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1825),
.B(n_1859),
.Y(n_2006)
);

INVxp67_ASAP7_75t_SL g2007 ( 
.A(n_1791),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1859),
.B(n_1863),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1801),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1790),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1779),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1880),
.B(n_1822),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1869),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1784),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1880),
.B(n_1835),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1782),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1805),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1903),
.B(n_1786),
.Y(n_2018)
);

AOI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_1901),
.A2(n_1917),
.B1(n_1910),
.B2(n_1923),
.C(n_1919),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1786),
.B(n_1856),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1884),
.B(n_1817),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1800),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1853),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1788),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1807),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1817),
.B(n_1836),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1904),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1807),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1930),
.B(n_1823),
.Y(n_2029)
);

INVx1_ASAP7_75t_SL g2030 ( 
.A(n_1797),
.Y(n_2030)
);

OR2x2_ASAP7_75t_L g2031 ( 
.A(n_1842),
.B(n_1812),
.Y(n_2031)
);

OAI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1977),
.A2(n_1921),
.B1(n_1926),
.B2(n_1927),
.Y(n_2032)
);

AOI211xp5_ASAP7_75t_L g2033 ( 
.A1(n_1947),
.A2(n_1810),
.B(n_1918),
.C(n_1894),
.Y(n_2033)
);

OAI221xp5_ASAP7_75t_L g2034 ( 
.A1(n_1977),
.A2(n_1826),
.B1(n_1815),
.B2(n_1932),
.C(n_1909),
.Y(n_2034)
);

OAI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_1974),
.A2(n_1881),
.B1(n_1773),
.B2(n_1916),
.Y(n_2035)
);

OAI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_1974),
.A2(n_1888),
.B1(n_1894),
.B2(n_1918),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_SL g2037 ( 
.A1(n_1986),
.A2(n_1840),
.B1(n_1907),
.B2(n_1893),
.Y(n_2037)
);

NOR4xp25_ASAP7_75t_SL g2038 ( 
.A(n_2019),
.B(n_1832),
.C(n_1813),
.D(n_1831),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1952),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1952),
.Y(n_2040)
);

CKINVDCx20_ASAP7_75t_R g2041 ( 
.A(n_1973),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1952),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_2024),
.Y(n_2043)
);

OAI211xp5_ASAP7_75t_SL g2044 ( 
.A1(n_2019),
.A2(n_1928),
.B(n_1823),
.C(n_1827),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2022),
.B(n_1916),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1952),
.Y(n_2046)
);

AO21x2_ASAP7_75t_L g2047 ( 
.A1(n_1942),
.A2(n_1888),
.B(n_1847),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1936),
.B(n_1902),
.Y(n_2048)
);

AO21x2_ASAP7_75t_L g2049 ( 
.A1(n_1942),
.A2(n_1799),
.B(n_1829),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1953),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_1944),
.B(n_1902),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1947),
.A2(n_1827),
.B1(n_1829),
.B2(n_1840),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1986),
.A2(n_1891),
.B1(n_1898),
.B2(n_1821),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1953),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2022),
.B(n_1891),
.Y(n_2055)
);

OAI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1959),
.A2(n_1844),
.B(n_1911),
.Y(n_2056)
);

AOI211xp5_ASAP7_75t_SL g2057 ( 
.A1(n_1967),
.A2(n_1844),
.B(n_1911),
.C(n_1850),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1937),
.B(n_1814),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1953),
.Y(n_2059)
);

AOI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_2026),
.A2(n_2015),
.B1(n_1967),
.B2(n_1959),
.Y(n_2060)
);

NAND3xp33_ASAP7_75t_L g2061 ( 
.A(n_2021),
.B(n_1814),
.C(n_1851),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_2015),
.A2(n_2018),
.B1(n_1999),
.B2(n_2000),
.Y(n_2062)
);

AOI21x1_ASAP7_75t_L g2063 ( 
.A1(n_1985),
.A2(n_1850),
.B(n_1873),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1954),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_2015),
.A2(n_1890),
.B1(n_1851),
.B2(n_1814),
.Y(n_2065)
);

AOI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_2026),
.A2(n_1814),
.B1(n_1851),
.B2(n_1890),
.C(n_1873),
.Y(n_2066)
);

AO21x2_ASAP7_75t_L g2067 ( 
.A1(n_1964),
.A2(n_1850),
.B(n_1851),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1954),
.Y(n_2068)
);

OAI22xp5_ASAP7_75t_SL g2069 ( 
.A1(n_2031),
.A2(n_1890),
.B1(n_1976),
.B2(n_1997),
.Y(n_2069)
);

AOI31xp33_ASAP7_75t_L g2070 ( 
.A1(n_2031),
.A2(n_1890),
.A3(n_1971),
.B(n_1997),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1954),
.Y(n_2071)
);

AOI21x1_ASAP7_75t_L g2072 ( 
.A1(n_1985),
.A2(n_2021),
.B(n_2027),
.Y(n_2072)
);

HB1xp67_ASAP7_75t_L g2073 ( 
.A(n_1949),
.Y(n_2073)
);

NAND2xp33_ASAP7_75t_R g2074 ( 
.A(n_1978),
.B(n_2001),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1937),
.B(n_1960),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_1944),
.B(n_1941),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1960),
.B(n_1957),
.Y(n_2077)
);

OAI211xp5_ASAP7_75t_L g2078 ( 
.A1(n_1968),
.A2(n_1950),
.B(n_2031),
.C(n_1975),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_2018),
.A2(n_2000),
.B1(n_1999),
.B2(n_1968),
.Y(n_2079)
);

NOR3xp33_ASAP7_75t_L g2080 ( 
.A(n_1971),
.B(n_1968),
.C(n_2014),
.Y(n_2080)
);

AOI22xp33_ASAP7_75t_L g2081 ( 
.A1(n_2018),
.A2(n_2000),
.B1(n_1999),
.B2(n_1950),
.Y(n_2081)
);

NAND3xp33_ASAP7_75t_SL g2082 ( 
.A(n_1971),
.B(n_2030),
.C(n_1962),
.Y(n_2082)
);

INVx3_ASAP7_75t_SL g2083 ( 
.A(n_2030),
.Y(n_2083)
);

OAI221xp5_ASAP7_75t_L g2084 ( 
.A1(n_2014),
.A2(n_2009),
.B1(n_2007),
.B2(n_1984),
.C(n_1990),
.Y(n_2084)
);

O2A1O1Ixp5_ASAP7_75t_L g2085 ( 
.A1(n_1950),
.A2(n_1982),
.B(n_1989),
.C(n_2009),
.Y(n_2085)
);

AOI322xp5_ASAP7_75t_L g2086 ( 
.A1(n_2012),
.A2(n_2006),
.A3(n_1996),
.B1(n_1995),
.B2(n_1982),
.C1(n_1989),
.C2(n_2029),
.Y(n_2086)
);

AO21x2_ASAP7_75t_L g2087 ( 
.A1(n_1964),
.A2(n_1980),
.B(n_1961),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1972),
.B(n_1938),
.Y(n_2088)
);

AOI221xp5_ASAP7_75t_L g2089 ( 
.A1(n_2010),
.A2(n_1982),
.B1(n_1989),
.B2(n_2012),
.C(n_1996),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2029),
.A2(n_2006),
.B1(n_2012),
.B2(n_1991),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1949),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1956),
.Y(n_2092)
);

OAI22xp5_ASAP7_75t_L g2093 ( 
.A1(n_1998),
.A2(n_1963),
.B1(n_1976),
.B2(n_1981),
.Y(n_2093)
);

INVx5_ASAP7_75t_L g2094 ( 
.A(n_1979),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1972),
.B(n_1938),
.Y(n_2095)
);

AOI211xp5_ASAP7_75t_L g2096 ( 
.A1(n_2002),
.A2(n_1975),
.B(n_2006),
.C(n_1969),
.Y(n_2096)
);

HB1xp67_ASAP7_75t_L g2097 ( 
.A(n_1988),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_1988),
.Y(n_2098)
);

BUFx6f_ASAP7_75t_L g2099 ( 
.A(n_2024),
.Y(n_2099)
);

OAI21x1_ASAP7_75t_SL g2100 ( 
.A1(n_1957),
.A2(n_1948),
.B(n_1945),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_1944),
.B(n_1941),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1941),
.B(n_1983),
.Y(n_2102)
);

NAND3xp33_ASAP7_75t_L g2103 ( 
.A(n_1990),
.B(n_2010),
.C(n_2011),
.Y(n_2103)
);

INVx5_ASAP7_75t_L g2104 ( 
.A(n_2094),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_2076),
.B(n_2025),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2073),
.B(n_2011),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_2094),
.B(n_1946),
.Y(n_2107)
);

NAND2x1_ASAP7_75t_L g2108 ( 
.A(n_2100),
.B(n_1978),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2050),
.Y(n_2109)
);

AOI22xp33_ASAP7_75t_L g2110 ( 
.A1(n_2032),
.A2(n_2029),
.B1(n_2020),
.B2(n_1998),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2091),
.B(n_1990),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2088),
.B(n_2095),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2076),
.B(n_2101),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2087),
.Y(n_2114)
);

NOR3xp33_ASAP7_75t_L g2115 ( 
.A(n_2034),
.B(n_2020),
.C(n_1990),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_R g2116 ( 
.A(n_2041),
.B(n_1943),
.Y(n_2116)
);

BUFx4f_ASAP7_75t_SL g2117 ( 
.A(n_2041),
.Y(n_2117)
);

NAND2x1p5_ASAP7_75t_L g2118 ( 
.A(n_2094),
.B(n_1978),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2101),
.B(n_1951),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2054),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2102),
.B(n_2025),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_2080),
.B(n_2013),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2100),
.B(n_1958),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2087),
.Y(n_2124)
);

BUFx2_ASAP7_75t_L g2125 ( 
.A(n_2067),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2097),
.B(n_2028),
.Y(n_2126)
);

AND2x4_ASAP7_75t_SL g2127 ( 
.A(n_2099),
.B(n_1981),
.Y(n_2127)
);

INVx4_ASAP7_75t_L g2128 ( 
.A(n_2083),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2054),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_2094),
.B(n_1940),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_2060),
.B(n_2075),
.Y(n_2131)
);

AND2x4_ASAP7_75t_L g2132 ( 
.A(n_2094),
.B(n_1940),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2068),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2077),
.B(n_1958),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2068),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2048),
.B(n_1969),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_2099),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_L g2138 ( 
.A(n_2083),
.B(n_1962),
.Y(n_2138)
);

INVx4_ASAP7_75t_L g2139 ( 
.A(n_2099),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2098),
.B(n_2028),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2087),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2040),
.B(n_1995),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2092),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2042),
.B(n_1965),
.Y(n_2144)
);

AND2x2_ASAP7_75t_L g2145 ( 
.A(n_2048),
.B(n_1969),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_2099),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2042),
.B(n_1965),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2046),
.B(n_1965),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_2064),
.B(n_1939),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2096),
.B(n_1984),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2051),
.B(n_1955),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2051),
.B(n_1955),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2071),
.B(n_1955),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2112),
.B(n_2043),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2114),
.Y(n_2155)
);

NAND2x1p5_ASAP7_75t_L g2156 ( 
.A(n_2104),
.B(n_2072),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2112),
.B(n_2043),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2111),
.B(n_2090),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2142),
.Y(n_2159)
);

INVx5_ASAP7_75t_SL g2160 ( 
.A(n_2130),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2142),
.Y(n_2161)
);

BUFx2_ASAP7_75t_L g2162 ( 
.A(n_2118),
.Y(n_2162)
);

NOR2x1_ASAP7_75t_L g2163 ( 
.A(n_2128),
.B(n_2082),
.Y(n_2163)
);

INVx1_ASAP7_75t_SL g2164 ( 
.A(n_2127),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2109),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2109),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2111),
.B(n_2049),
.Y(n_2167)
);

NOR2xp67_ASAP7_75t_L g2168 ( 
.A(n_2104),
.B(n_2078),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2114),
.Y(n_2169)
);

OAI22xp5_ASAP7_75t_L g2170 ( 
.A1(n_2110),
.A2(n_2033),
.B1(n_2052),
.B2(n_2070),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2120),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2114),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2112),
.B(n_2099),
.Y(n_2173)
);

AND2x2_ASAP7_75t_L g2174 ( 
.A(n_2151),
.B(n_2009),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2120),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_2104),
.B(n_2067),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2151),
.B(n_2152),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2123),
.B(n_2049),
.Y(n_2178)
);

NOR2xp33_ASAP7_75t_L g2179 ( 
.A(n_2117),
.B(n_2055),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2124),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2152),
.B(n_2009),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2124),
.Y(n_2182)
);

OR2x2_ASAP7_75t_L g2183 ( 
.A(n_2105),
.B(n_2049),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2105),
.B(n_2007),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2153),
.B(n_2067),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2153),
.B(n_2002),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2129),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_2123),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_L g2189 ( 
.A(n_2106),
.B(n_2086),
.Y(n_2189)
);

OR2x2_ASAP7_75t_L g2190 ( 
.A(n_2113),
.B(n_2039),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2129),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2133),
.Y(n_2192)
);

AOI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2115),
.A2(n_2036),
.B1(n_2037),
.B2(n_2044),
.Y(n_2193)
);

OAI33xp33_ASAP7_75t_L g2194 ( 
.A1(n_2150),
.A2(n_2035),
.A3(n_2093),
.B1(n_2103),
.B2(n_2053),
.B3(n_2045),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2124),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2133),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2135),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2119),
.B(n_2002),
.Y(n_2198)
);

NAND2x1p5_ASAP7_75t_L g2199 ( 
.A(n_2104),
.B(n_2072),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2113),
.B(n_2059),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2141),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2106),
.B(n_2121),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2119),
.B(n_2136),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2135),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2143),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2143),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2160),
.B(n_2136),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2165),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_2168),
.B(n_2104),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_2179),
.Y(n_2210)
);

INVx1_ASAP7_75t_SL g2211 ( 
.A(n_2164),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2165),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2166),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2166),
.Y(n_2214)
);

NAND3xp33_ASAP7_75t_L g2215 ( 
.A(n_2193),
.B(n_2115),
.C(n_2110),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2155),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2171),
.Y(n_2217)
);

OR2x2_ASAP7_75t_L g2218 ( 
.A(n_2202),
.B(n_2121),
.Y(n_2218)
);

NAND2xp33_ASAP7_75t_SL g2219 ( 
.A(n_2170),
.B(n_2116),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2171),
.Y(n_2220)
);

NAND4xp25_ASAP7_75t_L g2221 ( 
.A(n_2193),
.B(n_2085),
.C(n_2062),
.D(n_2079),
.Y(n_2221)
);

NAND4xp25_ASAP7_75t_L g2222 ( 
.A(n_2170),
.B(n_2081),
.C(n_2131),
.D(n_2089),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2189),
.B(n_2131),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2155),
.Y(n_2224)
);

NAND2x1_ASAP7_75t_L g2225 ( 
.A(n_2163),
.B(n_2128),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2189),
.B(n_2150),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2160),
.B(n_2145),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2194),
.A2(n_2047),
.B1(n_2122),
.B2(n_2069),
.Y(n_2228)
);

CKINVDCx16_ASAP7_75t_R g2229 ( 
.A(n_2163),
.Y(n_2229)
);

OAI33xp33_ASAP7_75t_L g2230 ( 
.A1(n_2178),
.A2(n_2134),
.A3(n_2126),
.B1(n_2140),
.B2(n_1994),
.B3(n_2144),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2175),
.Y(n_2231)
);

INVx3_ASAP7_75t_L g2232 ( 
.A(n_2160),
.Y(n_2232)
);

AND2x2_ASAP7_75t_L g2233 ( 
.A(n_2160),
.B(n_2145),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2155),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_2188),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2160),
.B(n_2137),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2175),
.Y(n_2237)
);

NAND3xp33_ASAP7_75t_L g2238 ( 
.A(n_2178),
.B(n_2038),
.C(n_2084),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2177),
.B(n_2137),
.Y(n_2239)
);

INVx1_ASAP7_75t_SL g2240 ( 
.A(n_2164),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_2168),
.B(n_2104),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2169),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2187),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2177),
.B(n_2137),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2198),
.B(n_2146),
.Y(n_2245)
);

NAND2xp33_ASAP7_75t_R g2246 ( 
.A(n_2162),
.B(n_2138),
.Y(n_2246)
);

OR2x2_ASAP7_75t_L g2247 ( 
.A(n_2202),
.B(n_2184),
.Y(n_2247)
);

AOI221xp5_ASAP7_75t_L g2248 ( 
.A1(n_2167),
.A2(n_2138),
.B1(n_2108),
.B2(n_2134),
.C(n_1994),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2187),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2158),
.B(n_2108),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2198),
.B(n_2146),
.Y(n_2251)
);

NOR3xp33_ASAP7_75t_L g2252 ( 
.A(n_2158),
.B(n_2128),
.C(n_2056),
.Y(n_2252)
);

NOR3xp33_ASAP7_75t_SL g2253 ( 
.A(n_2167),
.B(n_2074),
.C(n_2066),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2169),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2186),
.B(n_2146),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2191),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_R g2257 ( 
.A(n_2162),
.B(n_2117),
.Y(n_2257)
);

AOI21xp33_ASAP7_75t_L g2258 ( 
.A1(n_2225),
.A2(n_2183),
.B(n_2128),
.Y(n_2258)
);

NOR2x1_ASAP7_75t_L g2259 ( 
.A(n_2225),
.B(n_2215),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_2255),
.Y(n_2260)
);

OAI21xp33_ASAP7_75t_L g2261 ( 
.A1(n_2222),
.A2(n_2183),
.B(n_1963),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2229),
.B(n_2104),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2223),
.B(n_2174),
.Y(n_2263)
);

OAI32xp33_ASAP7_75t_L g2264 ( 
.A1(n_2229),
.A2(n_2156),
.A3(n_2199),
.B1(n_1998),
.B2(n_2184),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2208),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2208),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2212),
.Y(n_2267)
);

OAI222xp33_ASAP7_75t_L g2268 ( 
.A1(n_2228),
.A2(n_2156),
.B1(n_2199),
.B2(n_2118),
.C1(n_2186),
.C2(n_2185),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2226),
.B(n_2174),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2212),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2219),
.B(n_2118),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2207),
.B(n_2227),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2213),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2211),
.B(n_2240),
.Y(n_2274)
);

OAI21xp33_ASAP7_75t_L g2275 ( 
.A1(n_2238),
.A2(n_2181),
.B(n_2185),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2221),
.B(n_2181),
.Y(n_2276)
);

AOI211xp5_ASAP7_75t_L g2277 ( 
.A1(n_2252),
.A2(n_2020),
.B(n_1993),
.C(n_1991),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2253),
.B(n_2203),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2213),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2214),
.Y(n_2280)
);

OAI21xp33_ASAP7_75t_SL g2281 ( 
.A1(n_2207),
.A2(n_2203),
.B(n_2173),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2214),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2217),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2217),
.Y(n_2284)
);

OAI32xp33_ASAP7_75t_L g2285 ( 
.A1(n_2246),
.A2(n_2156),
.A3(n_2199),
.B1(n_2023),
.B2(n_2118),
.Y(n_2285)
);

OAI221xp5_ASAP7_75t_L g2286 ( 
.A1(n_2248),
.A2(n_2125),
.B1(n_2159),
.B2(n_2161),
.C(n_2200),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2235),
.B(n_2173),
.Y(n_2287)
);

OR2x2_ASAP7_75t_L g2288 ( 
.A(n_2247),
.B(n_2159),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2227),
.B(n_2154),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2220),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2255),
.Y(n_2291)
);

AOI22xp33_ASAP7_75t_L g2292 ( 
.A1(n_2257),
.A2(n_2047),
.B1(n_1993),
.B2(n_1991),
.Y(n_2292)
);

OAI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2210),
.A2(n_2001),
.B1(n_2013),
.B2(n_2023),
.Y(n_2293)
);

AOI21xp5_ASAP7_75t_L g2294 ( 
.A1(n_2230),
.A2(n_2047),
.B(n_2176),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_2210),
.B(n_2176),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2247),
.B(n_2161),
.Y(n_2296)
);

AOI31xp33_ASAP7_75t_L g2297 ( 
.A1(n_2236),
.A2(n_2057),
.A3(n_2061),
.B(n_2176),
.Y(n_2297)
);

OAI22xp5_ASAP7_75t_L g2298 ( 
.A1(n_2250),
.A2(n_2232),
.B1(n_2001),
.B2(n_2233),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_2272),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2259),
.B(n_2245),
.Y(n_2300)
);

OAI21xp5_ASAP7_75t_SL g2301 ( 
.A1(n_2275),
.A2(n_2232),
.B(n_2241),
.Y(n_2301)
);

OAI322xp33_ASAP7_75t_L g2302 ( 
.A1(n_2286),
.A2(n_2218),
.A3(n_2256),
.B1(n_2220),
.B2(n_2249),
.C1(n_2231),
.C2(n_2237),
.Y(n_2302)
);

OAI21xp33_ASAP7_75t_L g2303 ( 
.A1(n_2261),
.A2(n_2233),
.B(n_2218),
.Y(n_2303)
);

OAI221xp5_ASAP7_75t_L g2304 ( 
.A1(n_2277),
.A2(n_2232),
.B1(n_2236),
.B2(n_2251),
.C(n_2245),
.Y(n_2304)
);

OAI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_2292),
.A2(n_2209),
.B1(n_2241),
.B2(n_2244),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_2274),
.B(n_2278),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2276),
.B(n_2251),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2267),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2267),
.Y(n_2309)
);

AOI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2271),
.A2(n_2272),
.B1(n_2298),
.B2(n_2295),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_2289),
.B(n_2239),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2265),
.Y(n_2312)
);

OAI32xp33_ASAP7_75t_L g2313 ( 
.A1(n_2271),
.A2(n_2239),
.A3(n_2244),
.B1(n_2249),
.B2(n_2231),
.Y(n_2313)
);

AOI221xp5_ASAP7_75t_L g2314 ( 
.A1(n_2268),
.A2(n_2256),
.B1(n_2237),
.B2(n_2243),
.C(n_2241),
.Y(n_2314)
);

OAI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2293),
.A2(n_2209),
.B1(n_2241),
.B2(n_2013),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2266),
.Y(n_2316)
);

NOR2xp67_ASAP7_75t_SL g2317 ( 
.A(n_2262),
.B(n_1943),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2260),
.B(n_2291),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_SL g2319 ( 
.A(n_2285),
.B(n_2209),
.Y(n_2319)
);

AOI21xp33_ASAP7_75t_L g2320 ( 
.A1(n_2285),
.A2(n_2262),
.B(n_2295),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2260),
.B(n_2154),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2270),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2273),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2279),
.Y(n_2324)
);

OAI22xp33_ASAP7_75t_L g2325 ( 
.A1(n_2297),
.A2(n_2017),
.B1(n_1970),
.B2(n_1992),
.Y(n_2325)
);

INVx1_ASAP7_75t_SL g2326 ( 
.A(n_2291),
.Y(n_2326)
);

AOI222xp33_ASAP7_75t_L g2327 ( 
.A1(n_2264),
.A2(n_1993),
.B1(n_2004),
.B2(n_2005),
.C1(n_2003),
.C2(n_1966),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2289),
.B(n_2243),
.Y(n_2328)
);

AOI21xp33_ASAP7_75t_L g2329 ( 
.A1(n_2264),
.A2(n_2176),
.B(n_2242),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2311),
.Y(n_2330)
);

INVx1_ASAP7_75t_SL g2331 ( 
.A(n_2299),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2308),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2309),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2306),
.B(n_2263),
.Y(n_2334)
);

NAND2xp33_ASAP7_75t_L g2335 ( 
.A(n_2300),
.B(n_2287),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_2306),
.B(n_2258),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2326),
.B(n_2269),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2307),
.B(n_2294),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2312),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2316),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2328),
.B(n_2281),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2328),
.Y(n_2342)
);

CKINVDCx20_ASAP7_75t_R g2343 ( 
.A(n_2310),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_L g2344 ( 
.A(n_2304),
.B(n_2288),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2303),
.B(n_2280),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2322),
.Y(n_2346)
);

CKINVDCx16_ASAP7_75t_R g2347 ( 
.A(n_2319),
.Y(n_2347)
);

NOR2x1_ASAP7_75t_L g2348 ( 
.A(n_2325),
.B(n_2282),
.Y(n_2348)
);

OAI221xp5_ASAP7_75t_L g2349 ( 
.A1(n_2314),
.A2(n_2296),
.B1(n_2288),
.B2(n_2290),
.C(n_2284),
.Y(n_2349)
);

OA22x2_ASAP7_75t_L g2350 ( 
.A1(n_2301),
.A2(n_2283),
.B1(n_2127),
.B2(n_2139),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2318),
.B(n_2327),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2321),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2323),
.Y(n_2353)
);

OAI21xp33_ASAP7_75t_L g2354 ( 
.A1(n_2314),
.A2(n_2296),
.B(n_2004),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2330),
.B(n_2324),
.Y(n_2355)
);

OR2x2_ASAP7_75t_L g2356 ( 
.A(n_2331),
.B(n_2305),
.Y(n_2356)
);

AOI21xp5_ASAP7_75t_L g2357 ( 
.A1(n_2348),
.A2(n_2320),
.B(n_2302),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2342),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2342),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2330),
.B(n_2325),
.Y(n_2360)
);

AOI22xp5_ASAP7_75t_L g2361 ( 
.A1(n_2343),
.A2(n_2347),
.B1(n_2354),
.B2(n_2336),
.Y(n_2361)
);

A2O1A1Ixp33_ASAP7_75t_L g2362 ( 
.A1(n_2336),
.A2(n_2313),
.B(n_2317),
.C(n_2329),
.Y(n_2362)
);

INVx3_ASAP7_75t_SL g2363 ( 
.A(n_2343),
.Y(n_2363)
);

AOI221xp5_ASAP7_75t_L g2364 ( 
.A1(n_2349),
.A2(n_2315),
.B1(n_2254),
.B2(n_2242),
.C(n_2234),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2334),
.B(n_2190),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2352),
.B(n_2157),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2344),
.B(n_2157),
.Y(n_2367)
);

AOI222xp33_ASAP7_75t_L g2368 ( 
.A1(n_2351),
.A2(n_2125),
.B1(n_2005),
.B2(n_2004),
.C1(n_2216),
.C2(n_2224),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_2350),
.B(n_2127),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2363),
.B(n_2344),
.Y(n_2370)
);

O2A1O1Ixp33_ASAP7_75t_L g2371 ( 
.A1(n_2357),
.A2(n_2345),
.B(n_2335),
.C(n_2338),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2361),
.B(n_2352),
.Y(n_2372)
);

AOI221x1_ASAP7_75t_L g2373 ( 
.A1(n_2358),
.A2(n_2333),
.B1(n_2332),
.B2(n_2346),
.C(n_2340),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_SL g2374 ( 
.A(n_2356),
.B(n_2337),
.Y(n_2374)
);

AOI21xp5_ASAP7_75t_L g2375 ( 
.A1(n_2362),
.A2(n_2341),
.B(n_2350),
.Y(n_2375)
);

O2A1O1Ixp33_ASAP7_75t_L g2376 ( 
.A1(n_2360),
.A2(n_2359),
.B(n_2355),
.C(n_2368),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2368),
.A2(n_2353),
.B(n_2339),
.Y(n_2377)
);

OAI221xp5_ASAP7_75t_L g2378 ( 
.A1(n_2367),
.A2(n_2139),
.B1(n_2234),
.B2(n_2224),
.C(n_2216),
.Y(n_2378)
);

O2A1O1Ixp33_ASAP7_75t_SL g2379 ( 
.A1(n_2369),
.A2(n_2254),
.B(n_2206),
.C(n_2205),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_2365),
.B(n_2190),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2366),
.B(n_2200),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2374),
.B(n_2370),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2375),
.B(n_2364),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2373),
.Y(n_2384)
);

AOI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2372),
.A2(n_2380),
.B1(n_2381),
.B2(n_2377),
.Y(n_2385)
);

OAI211xp5_ASAP7_75t_L g2386 ( 
.A1(n_2371),
.A2(n_2139),
.B(n_1943),
.C(n_2065),
.Y(n_2386)
);

OAI21xp5_ASAP7_75t_SL g2387 ( 
.A1(n_2376),
.A2(n_2005),
.B(n_2063),
.Y(n_2387)
);

AOI221xp5_ASAP7_75t_L g2388 ( 
.A1(n_2379),
.A2(n_2180),
.B1(n_2182),
.B2(n_2169),
.C(n_2201),
.Y(n_2388)
);

NAND2xp33_ASAP7_75t_SL g2389 ( 
.A(n_2378),
.B(n_2139),
.Y(n_2389)
);

NAND3x1_ASAP7_75t_L g2390 ( 
.A(n_2370),
.B(n_2063),
.C(n_2205),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2382),
.Y(n_2391)
);

NAND3xp33_ASAP7_75t_SL g2392 ( 
.A(n_2383),
.B(n_1943),
.C(n_2126),
.Y(n_2392)
);

NOR4xp25_ASAP7_75t_L g2393 ( 
.A(n_2384),
.B(n_2172),
.C(n_2180),
.D(n_2201),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2385),
.Y(n_2394)
);

NAND4xp25_ASAP7_75t_SL g2395 ( 
.A(n_2386),
.B(n_2388),
.C(n_2387),
.D(n_2389),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2390),
.B(n_2191),
.Y(n_2396)
);

OAI211xp5_ASAP7_75t_L g2397 ( 
.A1(n_2383),
.A2(n_1943),
.B(n_2201),
.C(n_2172),
.Y(n_2397)
);

AOI211xp5_ASAP7_75t_L g2398 ( 
.A1(n_2383),
.A2(n_2107),
.B(n_2182),
.C(n_2172),
.Y(n_2398)
);

AOI211x1_ASAP7_75t_L g2399 ( 
.A1(n_2395),
.A2(n_2206),
.B(n_2204),
.C(n_2197),
.Y(n_2399)
);

NOR2x2_ASAP7_75t_L g2400 ( 
.A(n_2394),
.B(n_2180),
.Y(n_2400)
);

NOR3xp33_ASAP7_75t_SL g2401 ( 
.A(n_2392),
.B(n_2058),
.C(n_2197),
.Y(n_2401)
);

NAND5xp2_ASAP7_75t_L g2402 ( 
.A(n_2391),
.B(n_2008),
.C(n_1987),
.D(n_1992),
.E(n_2003),
.Y(n_2402)
);

NAND3xp33_ASAP7_75t_SL g2403 ( 
.A(n_2398),
.B(n_2140),
.C(n_2195),
.Y(n_2403)
);

OAI311xp33_ASAP7_75t_L g2404 ( 
.A1(n_2396),
.A2(n_2147),
.A3(n_2148),
.B1(n_2144),
.C1(n_2149),
.Y(n_2404)
);

OAI21xp5_ASAP7_75t_SL g2405 ( 
.A1(n_2397),
.A2(n_2107),
.B(n_2130),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2400),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_2401),
.B(n_2393),
.Y(n_2407)
);

BUFx2_ASAP7_75t_L g2408 ( 
.A(n_2399),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2403),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2409),
.B(n_2402),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2406),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2411),
.B(n_2407),
.Y(n_2412)
);

OAI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_2410),
.A2(n_2406),
.B1(n_2408),
.B2(n_2407),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2412),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2413),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2412),
.Y(n_2416)
);

AOI222xp33_ASAP7_75t_L g2417 ( 
.A1(n_2415),
.A2(n_2405),
.B1(n_2404),
.B2(n_2182),
.C1(n_2195),
.C2(n_2196),
.Y(n_2417)
);

AOI22xp33_ASAP7_75t_L g2418 ( 
.A1(n_2414),
.A2(n_2195),
.B1(n_2107),
.B2(n_2130),
.Y(n_2418)
);

AOI22xp5_ASAP7_75t_L g2419 ( 
.A1(n_2417),
.A2(n_2416),
.B1(n_2204),
.B2(n_2196),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2418),
.Y(n_2420)
);

NAND3xp33_ASAP7_75t_L g2421 ( 
.A(n_2420),
.B(n_2192),
.C(n_2141),
.Y(n_2421)
);

OAI221xp5_ASAP7_75t_R g2422 ( 
.A1(n_2421),
.A2(n_2419),
.B1(n_2192),
.B2(n_2130),
.C(n_2132),
.Y(n_2422)
);

AOI211xp5_ASAP7_75t_L g2423 ( 
.A1(n_2422),
.A2(n_2141),
.B(n_2107),
.C(n_2016),
.Y(n_2423)
);


endmodule