module fake_netlist_6_2565_n_957 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_957);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_957;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_120),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_32),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_54),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_104),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_141),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_125),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_140),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_99),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_27),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_6),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_95),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_97),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_35),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_115),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_9),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_43),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_175),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_83),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_137),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_142),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_136),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_56),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_18),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_55),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_6),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_29),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_65),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_7),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_3),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_7),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_46),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_144),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_22),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_147),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_89),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_59),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_17),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_91),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

BUFx2_ASAP7_75t_SL g240 ( 
.A(n_117),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_81),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_53),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_45),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_101),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_153),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_44),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_92),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_165),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_42),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_28),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_176),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_8),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_93),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_131),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_114),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_88),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_102),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_34),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_118),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_206),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_188),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_211),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_201),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_221),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_193),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_193),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_211),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_223),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_247),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_0),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_208),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_210),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_198),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_202),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_212),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_189),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_0),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_202),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_205),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_255),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_255),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_198),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_191),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_249),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_224),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_192),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_226),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_197),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_199),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_215),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_227),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_218),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_228),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_200),
.B(n_1),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_237),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_200),
.B(n_1),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_R g312 ( 
.A(n_190),
.B(n_2),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_220),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_198),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g315 ( 
.A(n_216),
.B(n_2),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_276),
.B(n_207),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_275),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_264),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_266),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_216),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_209),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_297),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_301),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_251),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_293),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_294),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_293),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_279),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_288),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

AND2x6_ASAP7_75t_L g337 ( 
.A(n_281),
.B(n_258),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_305),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_268),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_277),
.B(n_222),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_282),
.B(n_190),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_304),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_271),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_267),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_281),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_273),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_267),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_307),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_274),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_265),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_270),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_268),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_285),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_272),
.B(n_263),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_290),
.B(n_195),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_313),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_222),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_302),
.B(n_195),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_310),
.B(n_196),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_309),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_310),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_312),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_R g368 ( 
.A(n_306),
.B(n_234),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_286),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_296),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_306),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_299),
.Y(n_373)
);

OR2x6_ASAP7_75t_L g374 ( 
.A(n_328),
.B(n_284),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_296),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_369),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_235),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_229),
.Y(n_378)
);

NOR3xp33_ASAP7_75t_SL g379 ( 
.A(n_367),
.B(n_244),
.C(n_196),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_338),
.Y(n_380)
);

BUFx4f_ASAP7_75t_L g381 ( 
.A(n_369),
.Y(n_381)
);

BUFx8_ASAP7_75t_SL g382 ( 
.A(n_340),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_320),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_365),
.A2(n_229),
.B1(n_260),
.B2(n_292),
.Y(n_384)
);

OR2x6_ASAP7_75t_L g385 ( 
.A(n_330),
.B(n_240),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_327),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_352),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_358),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_260),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_344),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_347),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_320),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_365),
.B(n_236),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_337),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_203),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_322),
.B(n_238),
.Y(n_399)
);

AND2x2_ASAP7_75t_SL g400 ( 
.A(n_323),
.B(n_204),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_348),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_244),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_337),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_341),
.B(n_213),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_341),
.B(n_214),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_364),
.B(n_308),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_325),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_341),
.B(n_217),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_358),
.B(n_308),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_316),
.Y(n_412)
);

NAND3x1_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_231),
.C(n_225),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_316),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_336),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_359),
.A2(n_295),
.B1(n_294),
.B2(n_253),
.Y(n_416)
);

AND3x2_ASAP7_75t_L g417 ( 
.A(n_333),
.B(n_239),
.C(n_232),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_369),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_SL g419 ( 
.A(n_368),
.B(n_295),
.C(n_287),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_319),
.B(n_241),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_371),
.B(n_253),
.Y(n_421)
);

OR2x6_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_243),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_363),
.B(n_254),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_343),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_319),
.B(n_245),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_363),
.B(n_373),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_369),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_331),
.B(n_256),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_353),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_372),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_370),
.B(n_254),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_370),
.B(n_257),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_317),
.A2(n_257),
.B1(n_242),
.B2(n_250),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_321),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_353),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_327),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_L g437 ( 
.A(n_370),
.B(n_246),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_362),
.A2(n_259),
.B1(n_248),
.B2(n_269),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_355),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_362),
.A2(n_291),
.B1(n_287),
.B2(n_269),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_331),
.B(n_33),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_342),
.B(n_36),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_370),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_327),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_317),
.B(n_342),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_321),
.B(n_291),
.Y(n_446)
);

BUFx4f_ASAP7_75t_L g447 ( 
.A(n_370),
.Y(n_447)
);

INVx4_ASAP7_75t_SL g448 ( 
.A(n_337),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_412),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_375),
.B(n_362),
.Y(n_450)
);

AOI221xp5_ASAP7_75t_L g451 ( 
.A1(n_438),
.A2(n_360),
.B1(n_366),
.B2(n_361),
.C(n_350),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_399),
.B(n_356),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_411),
.Y(n_453)
);

O2A1O1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_378),
.A2(n_355),
.B(n_351),
.C(n_356),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_389),
.B(n_366),
.Y(n_455)
);

OAI22xp33_ASAP7_75t_L g456 ( 
.A1(n_404),
.A2(n_361),
.B1(n_332),
.B2(n_350),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_423),
.B(n_332),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_377),
.B(n_334),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_396),
.B(n_334),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_400),
.B(n_339),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_339),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_378),
.B(n_335),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_390),
.B(n_351),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_390),
.B(n_429),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_430),
.B(n_329),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_426),
.B(n_345),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_335),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_392),
.B(n_327),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_393),
.B(n_346),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_394),
.B(n_406),
.Y(n_471)
);

NOR3xp33_ASAP7_75t_L g472 ( 
.A(n_419),
.B(n_329),
.C(n_372),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_442),
.A2(n_345),
.B1(n_337),
.B2(n_349),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_409),
.B(n_415),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_424),
.B(n_346),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_387),
.B(n_346),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_398),
.B(n_346),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_376),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_418),
.Y(n_479)
);

BUFx8_ASAP7_75t_L g480 ( 
.A(n_382),
.Y(n_480)
);

NAND2x1p5_ASAP7_75t_L g481 ( 
.A(n_397),
.B(n_349),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g482 ( 
.A(n_402),
.B(n_349),
.C(n_354),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_404),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_439),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_384),
.A2(n_433),
.B1(n_385),
.B2(n_410),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_391),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_398),
.B(n_346),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_421),
.B(n_3),
.Y(n_489)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_442),
.A2(n_337),
.B1(n_5),
.B2(n_9),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_442),
.A2(n_337),
.B1(n_5),
.B2(n_10),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_405),
.B(n_337),
.Y(n_492)
);

OAI22xp33_ASAP7_75t_L g493 ( 
.A1(n_405),
.A2(n_4),
.B1(n_10),
.B2(n_11),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_401),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_410),
.B(n_37),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_374),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_431),
.B(n_4),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_436),
.B(n_427),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_397),
.B(n_38),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_408),
.B(n_434),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_432),
.B(n_11),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_442),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_443),
.B(n_39),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_385),
.A2(n_90),
.B1(n_184),
.B2(n_183),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_444),
.B(n_40),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_386),
.B(n_41),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_385),
.A2(n_94),
.B1(n_182),
.B2(n_181),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_420),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_397),
.B(n_403),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_386),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_434),
.B(n_12),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_374),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_397),
.B(n_47),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_386),
.B(n_388),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_416),
.B(n_13),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_379),
.B(n_48),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_403),
.B(n_49),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_430),
.B(n_14),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_388),
.B(n_50),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_440),
.B(n_15),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_374),
.B(n_15),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_388),
.B(n_51),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_428),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_527)
);

AO22x1_ASAP7_75t_L g528 ( 
.A1(n_383),
.A2(n_395),
.B1(n_413),
.B2(n_446),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_381),
.B(n_52),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_428),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_441),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_455),
.B(n_422),
.Y(n_532)
);

A2O1A1Ixp33_ASAP7_75t_L g533 ( 
.A1(n_489),
.A2(n_381),
.B(n_447),
.C(n_441),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_489),
.A2(n_509),
.B(n_519),
.C(n_510),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_451),
.B(n_422),
.C(n_437),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_531),
.B(n_448),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_524),
.B(n_422),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_524),
.A2(n_447),
.B(n_403),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_465),
.A2(n_403),
.B(n_448),
.Y(n_539)
);

NOR3xp33_ASAP7_75t_L g540 ( 
.A(n_457),
.B(n_417),
.C(n_19),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_503),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_480),
.Y(n_542)
);

AOI21x1_ASAP7_75t_L g543 ( 
.A1(n_464),
.A2(n_492),
.B(n_463),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_530),
.A2(n_448),
.B(n_108),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_450),
.B(n_20),
.Y(n_546)
);

NOR2x1_ASAP7_75t_L g547 ( 
.A(n_458),
.B(n_459),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_483),
.B(n_21),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_503),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_449),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_449),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_530),
.A2(n_109),
.B(n_180),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_467),
.B(n_23),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_456),
.B(n_57),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_467),
.B(n_58),
.Y(n_555)
);

NAND2x1p5_ASAP7_75t_L g556 ( 
.A(n_478),
.B(n_60),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_452),
.B(n_24),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_480),
.Y(n_558)
);

NOR2x1_ASAP7_75t_L g559 ( 
.A(n_482),
.B(n_61),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_460),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_501),
.B(n_25),
.Y(n_561)
);

A2O1A1Ixp33_ASAP7_75t_L g562 ( 
.A1(n_498),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_562)
);

A2O1A1Ixp33_ASAP7_75t_L g563 ( 
.A1(n_498),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_531),
.A2(n_499),
.B(n_488),
.Y(n_564)
);

INVx3_ASAP7_75t_SL g565 ( 
.A(n_466),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_471),
.B(n_30),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_490),
.A2(n_30),
.B1(n_31),
.B2(n_62),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_490),
.A2(n_31),
.B1(n_63),
.B2(n_64),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_485),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_477),
.A2(n_66),
.B(n_67),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_486),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_453),
.B(n_71),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_464),
.A2(n_72),
.B(n_73),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_474),
.B(n_468),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_502),
.B(n_74),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_516),
.A2(n_75),
.B(n_76),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_521),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_484),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_514),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_502),
.B(n_77),
.Y(n_581)
);

AO21x1_ASAP7_75t_L g582 ( 
.A1(n_496),
.A2(n_78),
.B(n_79),
.Y(n_582)
);

O2A1O1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_461),
.A2(n_80),
.B(n_82),
.C(n_84),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_461),
.B(n_523),
.Y(n_584)
);

AO21x1_ASAP7_75t_L g585 ( 
.A1(n_454),
.A2(n_85),
.B(n_86),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_517),
.B(n_87),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_484),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_511),
.A2(n_96),
.B(n_98),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_497),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_487),
.A2(n_100),
.B1(n_103),
.B2(n_106),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_513),
.B(n_107),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_511),
.A2(n_110),
.B(n_111),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_525),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_494),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_564),
.A2(n_473),
.B(n_529),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_538),
.A2(n_473),
.B(n_504),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_556),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_580),
.B(n_479),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_570),
.B(n_479),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_547),
.B(n_491),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_543),
.A2(n_506),
.B(n_526),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_534),
.B(n_495),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_538),
.A2(n_522),
.B(n_507),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_551),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_550),
.Y(n_605)
);

OAI21x1_ASAP7_75t_L g606 ( 
.A1(n_544),
.A2(n_469),
.B(n_470),
.Y(n_606)
);

AND3x4_ASAP7_75t_L g607 ( 
.A(n_542),
.B(n_472),
.C(n_518),
.Y(n_607)
);

OAI21x1_ASAP7_75t_L g608 ( 
.A1(n_560),
.A2(n_475),
.B(n_476),
.Y(n_608)
);

AND2x2_ASAP7_75t_SL g609 ( 
.A(n_586),
.B(n_491),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_558),
.Y(n_610)
);

AOI21x1_ASAP7_75t_L g611 ( 
.A1(n_555),
.A2(n_500),
.B(n_520),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_567),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_541),
.A2(n_527),
.B1(n_508),
.B2(n_493),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_579),
.A2(n_512),
.B(n_481),
.Y(n_614)
);

BUFx12f_ASAP7_75t_L g615 ( 
.A(n_532),
.Y(n_615)
);

AO21x2_ASAP7_75t_L g616 ( 
.A1(n_533),
.A2(n_500),
.B(n_520),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_587),
.Y(n_617)
);

NAND2x1_ASAP7_75t_L g618 ( 
.A(n_536),
.B(n_512),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_555),
.A2(n_539),
.B(n_581),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_584),
.B(n_478),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_552),
.A2(n_481),
.B(n_515),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_537),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_576),
.A2(n_515),
.B(n_505),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_574),
.A2(n_571),
.B(n_577),
.Y(n_624)
);

NAND2x1p5_ASAP7_75t_L g625 ( 
.A(n_559),
.B(n_518),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_545),
.B(n_518),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_556),
.B(n_528),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_553),
.B(n_527),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_588),
.A2(n_112),
.B(n_113),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_537),
.A2(n_116),
.B(n_119),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_546),
.A2(n_185),
.B(n_122),
.Y(n_631)
);

AO31x2_ASAP7_75t_L g632 ( 
.A1(n_585),
.A2(n_121),
.A3(n_123),
.B(n_127),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_557),
.B(n_128),
.Y(n_633)
);

A2O1A1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_535),
.A2(n_129),
.B(n_130),
.C(n_133),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_569),
.A2(n_554),
.B(n_591),
.Y(n_635)
);

AOI21x1_ASAP7_75t_SL g636 ( 
.A1(n_566),
.A2(n_134),
.B(n_139),
.Y(n_636)
);

AO31x2_ASAP7_75t_L g637 ( 
.A1(n_582),
.A2(n_143),
.A3(n_148),
.B(n_149),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_565),
.B(n_150),
.Y(n_638)
);

AOI21x1_ASAP7_75t_L g639 ( 
.A1(n_548),
.A2(n_151),
.B(n_154),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_578),
.B(n_155),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_589),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_561),
.B(n_156),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_593),
.Y(n_643)
);

AOI21x1_ASAP7_75t_SL g644 ( 
.A1(n_573),
.A2(n_159),
.B(n_160),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_592),
.A2(n_161),
.B(n_162),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_609),
.B(n_541),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_605),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_615),
.B(n_572),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_594),
.B(n_549),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_610),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_594),
.B(n_549),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_643),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_622),
.B(n_569),
.Y(n_653)
);

BUFx12f_ASAP7_75t_L g654 ( 
.A(n_638),
.Y(n_654)
);

NAND2x1p5_ASAP7_75t_L g655 ( 
.A(n_597),
.B(n_590),
.Y(n_655)
);

O2A1O1Ixp5_ASAP7_75t_L g656 ( 
.A1(n_635),
.A2(n_568),
.B(n_563),
.C(n_562),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_617),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_620),
.B(n_568),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_627),
.B(n_583),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_604),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_598),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_620),
.B(n_599),
.Y(n_662)
);

AOI21xp33_ASAP7_75t_SL g663 ( 
.A1(n_607),
.A2(n_540),
.B(n_164),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_599),
.B(n_163),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_597),
.B(n_628),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_598),
.B(n_536),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_619),
.A2(n_595),
.B(n_623),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_612),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_641),
.B(n_166),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_613),
.A2(n_536),
.B1(n_168),
.B2(n_169),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_596),
.A2(n_536),
.B(n_170),
.Y(n_671)
);

NAND2x1p5_ASAP7_75t_L g672 ( 
.A(n_597),
.B(n_167),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_640),
.B(n_171),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_626),
.B(n_172),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_627),
.B(n_173),
.Y(n_675)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_612),
.Y(n_676)
);

INVx8_ASAP7_75t_L g677 ( 
.A(n_627),
.Y(n_677)
);

AOI21x1_ASAP7_75t_L g678 ( 
.A1(n_611),
.A2(n_177),
.B(n_178),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_642),
.B(n_600),
.Y(n_679)
);

BUFx10_ASAP7_75t_L g680 ( 
.A(n_636),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_642),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_628),
.B(n_625),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_613),
.B(n_602),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_618),
.Y(n_684)
);

AOI222xp33_ASAP7_75t_L g685 ( 
.A1(n_631),
.A2(n_602),
.B1(n_634),
.B2(n_633),
.C1(n_645),
.C2(n_629),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_633),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_608),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_625),
.A2(n_631),
.B1(n_616),
.B2(n_630),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_639),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_616),
.A2(n_630),
.B1(n_624),
.B2(n_603),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_644),
.A2(n_632),
.B1(n_637),
.B2(n_621),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_637),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_606),
.B(n_632),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_632),
.A2(n_637),
.B1(n_614),
.B2(n_601),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_609),
.B(n_594),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_650),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_647),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_695),
.B(n_662),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_657),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_677),
.B(n_659),
.Y(n_700)
);

BUFx8_ASAP7_75t_L g701 ( 
.A(n_654),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_652),
.Y(n_702)
);

OAI22xp33_ASAP7_75t_L g703 ( 
.A1(n_646),
.A2(n_695),
.B1(n_681),
.B2(n_683),
.Y(n_703)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_667),
.A2(n_678),
.B(n_687),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_691),
.A2(n_694),
.B(n_693),
.Y(n_705)
);

BUFx2_ASAP7_75t_R g706 ( 
.A(n_661),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_SL g707 ( 
.A1(n_646),
.A2(n_677),
.B1(n_670),
.B2(n_675),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_660),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_649),
.A2(n_658),
.B1(n_651),
.B2(n_679),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_694),
.A2(n_671),
.B(n_690),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_679),
.B(n_651),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_666),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_668),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_656),
.A2(n_686),
.B(n_688),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_653),
.A2(n_648),
.B1(n_659),
.B2(n_655),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_676),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_653),
.Y(n_717)
);

AOI21x1_ASAP7_75t_L g718 ( 
.A1(n_691),
.A2(n_689),
.B(n_659),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_677),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_682),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_SL g721 ( 
.A1(n_670),
.A2(n_674),
.B1(n_673),
.B2(n_655),
.Y(n_721)
);

NAND2x1p5_ASAP7_75t_L g722 ( 
.A(n_666),
.B(n_664),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_665),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_669),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_672),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_672),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_680),
.Y(n_727)
);

CKINVDCx11_ASAP7_75t_R g728 ( 
.A(n_680),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_684),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_684),
.Y(n_730)
);

AND2x4_ASAP7_75t_L g731 ( 
.A(n_684),
.B(n_692),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_663),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_685),
.B(n_662),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_685),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_646),
.A2(n_609),
.B1(n_613),
.B2(n_549),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_652),
.Y(n_736)
);

BUFx2_ASAP7_75t_R g737 ( 
.A(n_650),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_647),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_684),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_652),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_647),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_647),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_647),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_647),
.Y(n_744)
);

AO21x1_ASAP7_75t_L g745 ( 
.A1(n_683),
.A2(n_549),
.B(n_541),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_647),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_647),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_647),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_683),
.B(n_503),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_647),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_662),
.B(n_648),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_647),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_741),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_733),
.B(n_720),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_704),
.A2(n_710),
.B(n_705),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_704),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_700),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_711),
.B(n_734),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_741),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_742),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_746),
.Y(n_761)
);

AO21x2_ASAP7_75t_L g762 ( 
.A1(n_714),
.A2(n_718),
.B(n_710),
.Y(n_762)
);

AO21x2_ASAP7_75t_L g763 ( 
.A1(n_711),
.A2(n_749),
.B(n_715),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_746),
.Y(n_764)
);

AO21x2_ASAP7_75t_L g765 ( 
.A1(n_749),
.A2(n_745),
.B(n_717),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_731),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_700),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_709),
.B(n_698),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_700),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_747),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_748),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_696),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_734),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_723),
.A2(n_709),
.B(n_748),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_752),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_752),
.Y(n_776)
);

AO21x2_ASAP7_75t_L g777 ( 
.A1(n_703),
.A2(n_744),
.B(n_697),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_700),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_731),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_699),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_738),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_743),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_750),
.Y(n_783)
);

NAND3xp33_ASAP7_75t_L g784 ( 
.A(n_735),
.B(n_721),
.C(n_734),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_734),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_731),
.B(n_725),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_708),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_735),
.B(n_713),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_726),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_716),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_708),
.B(n_751),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_727),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_732),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_739),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_729),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_772),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_792),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_780),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_762),
.B(n_707),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_762),
.B(n_724),
.Y(n_800)
);

OAI33xp33_ASAP7_75t_L g801 ( 
.A1(n_793),
.A2(n_730),
.A3(n_696),
.B1(n_728),
.B2(n_740),
.B3(n_706),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_762),
.B(n_751),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_762),
.B(n_751),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_790),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_762),
.B(n_739),
.Y(n_805)
);

AO31x2_ASAP7_75t_L g806 ( 
.A1(n_756),
.A2(n_712),
.A3(n_728),
.B(n_739),
.Y(n_806)
);

OR2x2_ASAP7_75t_L g807 ( 
.A(n_763),
.B(n_702),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_784),
.A2(n_736),
.B1(n_701),
.B2(n_722),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_780),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_763),
.B(n_719),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_763),
.B(n_719),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_763),
.B(n_722),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_780),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_763),
.B(n_737),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_757),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_765),
.B(n_701),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_780),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_765),
.B(n_701),
.Y(n_818)
);

OA21x2_ASAP7_75t_L g819 ( 
.A1(n_755),
.A2(n_756),
.B(n_774),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_782),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_757),
.Y(n_821)
);

OAI221xp5_ASAP7_75t_SL g822 ( 
.A1(n_808),
.A2(n_784),
.B1(n_758),
.B2(n_785),
.C(n_768),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_797),
.B(n_754),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_801),
.A2(n_773),
.B1(n_785),
.B2(n_778),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_797),
.B(n_754),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_815),
.B(n_754),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_800),
.B(n_758),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_800),
.B(n_758),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_814),
.A2(n_773),
.B1(n_768),
.B2(n_765),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_815),
.B(n_769),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_814),
.A2(n_773),
.B1(n_765),
.B2(n_788),
.Y(n_831)
);

NAND2x1_ASAP7_75t_L g832 ( 
.A(n_800),
.B(n_790),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_801),
.B(n_793),
.C(n_767),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_816),
.B(n_790),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_SL g835 ( 
.A1(n_814),
.A2(n_773),
.B(n_757),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_816),
.B(n_782),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_816),
.B(n_782),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_L g838 ( 
.A(n_807),
.B(n_773),
.C(n_792),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_807),
.B(n_773),
.C(n_769),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_808),
.A2(n_774),
.B(n_767),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_L g841 ( 
.A(n_807),
.B(n_773),
.C(n_791),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_818),
.B(n_782),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_SL g843 ( 
.A1(n_799),
.A2(n_773),
.B1(n_757),
.B2(n_778),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_823),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_843),
.B(n_803),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_827),
.B(n_811),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_826),
.B(n_830),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_828),
.B(n_811),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_831),
.B(n_802),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_825),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_836),
.B(n_818),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_837),
.Y(n_852)
);

NAND2x1_ASAP7_75t_SL g853 ( 
.A(n_835),
.B(n_818),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_842),
.B(n_811),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_834),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_831),
.B(n_802),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_833),
.B(n_765),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_832),
.B(n_802),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_855),
.B(n_841),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_849),
.A2(n_799),
.B1(n_812),
.B2(n_829),
.Y(n_860)
);

NOR2x1_ASAP7_75t_L g861 ( 
.A(n_857),
.B(n_838),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_847),
.B(n_803),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_846),
.Y(n_863)
);

NOR2x1p5_ASAP7_75t_L g864 ( 
.A(n_845),
.B(n_796),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_L g865 ( 
.A(n_844),
.B(n_824),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_851),
.B(n_829),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_850),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_864),
.B(n_858),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_862),
.B(n_858),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_863),
.B(n_847),
.Y(n_870)
);

NAND2x1p5_ASAP7_75t_L g871 ( 
.A(n_861),
.B(n_812),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_867),
.B(n_852),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_863),
.B(n_845),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_859),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_866),
.B(n_856),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_865),
.B(n_856),
.Y(n_876)
);

AOI21xp33_ASAP7_75t_L g877 ( 
.A1(n_860),
.A2(n_849),
.B(n_839),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_872),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_870),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_874),
.B(n_848),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_873),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_876),
.A2(n_799),
.B1(n_840),
.B2(n_812),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_879),
.B(n_868),
.Y(n_883)
);

OAI221xp5_ASAP7_75t_L g884 ( 
.A1(n_882),
.A2(n_876),
.B1(n_877),
.B2(n_871),
.C(n_875),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_881),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_880),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_886),
.B(n_878),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_885),
.Y(n_888)
);

CKINVDCx16_ASAP7_75t_R g889 ( 
.A(n_883),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_883),
.B(n_868),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_889),
.Y(n_891)
);

OAI21xp33_ASAP7_75t_SL g892 ( 
.A1(n_890),
.A2(n_884),
.B(n_877),
.Y(n_892)
);

AOI221xp5_ASAP7_75t_L g893 ( 
.A1(n_888),
.A2(n_882),
.B1(n_871),
.B2(n_822),
.C(n_810),
.Y(n_893)
);

AOI322xp5_ASAP7_75t_L g894 ( 
.A1(n_890),
.A2(n_869),
.A3(n_803),
.B1(n_810),
.B2(n_853),
.C1(n_805),
.C2(n_788),
.Y(n_894)
);

OAI21xp33_ASAP7_75t_SL g895 ( 
.A1(n_887),
.A2(n_848),
.B(n_846),
.Y(n_895)
);

NAND4xp25_ASAP7_75t_L g896 ( 
.A(n_887),
.B(n_810),
.C(n_795),
.D(n_778),
.Y(n_896)
);

AOI21x1_ASAP7_75t_L g897 ( 
.A1(n_888),
.A2(n_795),
.B(n_781),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_889),
.A2(n_777),
.B(n_783),
.Y(n_898)
);

AOI211x1_ASAP7_75t_L g899 ( 
.A1(n_896),
.A2(n_805),
.B(n_781),
.C(n_783),
.Y(n_899)
);

AND3x4_ASAP7_75t_L g900 ( 
.A(n_891),
.B(n_778),
.C(n_821),
.Y(n_900)
);

NAND3xp33_ASAP7_75t_L g901 ( 
.A(n_892),
.B(n_805),
.C(n_789),
.Y(n_901)
);

AOI21xp33_ASAP7_75t_SL g902 ( 
.A1(n_895),
.A2(n_893),
.B(n_894),
.Y(n_902)
);

AOI21xp33_ASAP7_75t_L g903 ( 
.A1(n_898),
.A2(n_777),
.B(n_767),
.Y(n_903)
);

NOR3xp33_ASAP7_75t_L g904 ( 
.A(n_897),
.B(n_789),
.C(n_794),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_891),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_902),
.B(n_854),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_901),
.A2(n_789),
.B(n_821),
.C(n_815),
.Y(n_907)
);

AOI221xp5_ASAP7_75t_L g908 ( 
.A1(n_905),
.A2(n_794),
.B1(n_786),
.B2(n_788),
.C(n_760),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_SL g909 ( 
.A(n_900),
.B(n_770),
.C(n_791),
.Y(n_909)
);

INVxp33_ASAP7_75t_L g910 ( 
.A(n_904),
.Y(n_910)
);

NOR2x1_ASAP7_75t_L g911 ( 
.A(n_899),
.B(n_777),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_903),
.B(n_786),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_905),
.B(n_794),
.C(n_786),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_902),
.A2(n_794),
.B1(n_786),
.B2(n_759),
.C(n_760),
.Y(n_914)
);

NOR3xp33_ASAP7_75t_SL g915 ( 
.A(n_905),
.B(n_787),
.C(n_753),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_915),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_914),
.B(n_806),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_906),
.A2(n_909),
.B1(n_912),
.B2(n_910),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_913),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_908),
.A2(n_786),
.B1(n_777),
.B2(n_791),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_911),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_907),
.B(n_806),
.Y(n_922)
);

NOR2x1p5_ASAP7_75t_L g923 ( 
.A(n_909),
.B(n_821),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_906),
.A2(n_777),
.B1(n_766),
.B2(n_779),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_915),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_911),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_L g927 ( 
.A(n_921),
.B(n_794),
.C(n_753),
.Y(n_927)
);

NAND4xp75_ASAP7_75t_L g928 ( 
.A(n_918),
.B(n_779),
.C(n_819),
.D(n_764),
.Y(n_928)
);

OAI211xp5_ASAP7_75t_L g929 ( 
.A1(n_916),
.A2(n_804),
.B(n_770),
.C(n_775),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_926),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_925),
.A2(n_779),
.B1(n_766),
.B2(n_804),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_919),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_922),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_930),
.Y(n_934)
);

NAND3x1_ASAP7_75t_L g935 ( 
.A(n_932),
.B(n_917),
.C(n_920),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_933),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_L g937 ( 
.A(n_927),
.B(n_924),
.Y(n_937)
);

OR2x2_ASAP7_75t_L g938 ( 
.A(n_931),
.B(n_929),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_928),
.B(n_923),
.Y(n_939)
);

XOR2xp5_ASAP7_75t_L g940 ( 
.A(n_934),
.B(n_787),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_938),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_939),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_936),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_943),
.B(n_935),
.Y(n_944)
);

AOI221xp5_ASAP7_75t_L g945 ( 
.A1(n_941),
.A2(n_937),
.B1(n_759),
.B2(n_775),
.C(n_764),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_944),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_945),
.A2(n_942),
.B(n_940),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_946),
.A2(n_771),
.B1(n_766),
.B2(n_809),
.Y(n_948)
);

XNOR2x1_ASAP7_75t_L g949 ( 
.A(n_947),
.B(n_774),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_946),
.A2(n_771),
.B(n_761),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_SL g951 ( 
.A1(n_948),
.A2(n_766),
.B1(n_809),
.B2(n_820),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_949),
.A2(n_950),
.B(n_755),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_949),
.A2(n_776),
.B(n_761),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_952),
.A2(n_776),
.B(n_761),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_954),
.A2(n_951),
.B1(n_953),
.B2(n_766),
.Y(n_955)
);

AOI221xp5_ASAP7_75t_L g956 ( 
.A1(n_955),
.A2(n_820),
.B1(n_817),
.B2(n_813),
.C(n_798),
.Y(n_956)
);

AOI211xp5_ASAP7_75t_L g957 ( 
.A1(n_956),
.A2(n_798),
.B(n_817),
.C(n_813),
.Y(n_957)
);


endmodule