module real_jpeg_18797_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_469),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_0),
.B(n_470),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_1),
.A2(n_14),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_1),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_1),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_1),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_1),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_1),
.B(n_413),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_2),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_2),
.Y(n_159)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_2),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_3),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_3),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_3),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_3),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_3),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_3),
.B(n_452),
.Y(n_451)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_4),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_4),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_4),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_4),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_4),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_4),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_4),
.B(n_155),
.Y(n_385)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_5),
.Y(n_345)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_5),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_75),
.Y(n_74)
);

NAND2x1p5_ASAP7_75t_L g95 ( 
.A(n_6),
.B(n_71),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_6),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_6),
.B(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_6),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_6),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_6),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_6),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_7),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_7),
.B(n_237),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_7),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_7),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_7),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_7),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_7),
.B(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_8),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_9),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_9),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_9),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_9),
.B(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_9),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_10),
.Y(n_269)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_11),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_12),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_12),
.Y(n_143)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_12),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_13),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_13),
.B(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_13),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_13),
.B(n_361),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_13),
.B(n_165),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_13),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_13),
.B(n_413),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_14),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_14),
.B(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_14),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_14),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_14),
.B(n_450),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_16),
.Y(n_124)
);

BUFx4f_ASAP7_75t_L g210 ( 
.A(n_16),
.Y(n_210)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g302 ( 
.A(n_17),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g454 ( 
.A(n_17),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_436),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2x1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_327),
.Y(n_21)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_223),
.B(n_286),
.C(n_287),
.D(n_326),
.Y(n_22)
);

NAND4xp25_ASAP7_75t_L g327 ( 
.A(n_23),
.B(n_287),
.C(n_328),
.D(n_330),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_176),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_24),
.B(n_176),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_100),
.C(n_146),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_25),
.A2(n_26),
.B1(n_101),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_66),
.Y(n_26)
);

INVxp33_ASAP7_75t_SL g178 ( 
.A(n_27),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_41),
.C(n_49),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_28),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_29),
.B(n_33),
.C(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_30),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_36),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_37),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_37),
.B(n_207),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_38),
.Y(n_248)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_40),
.B(n_207),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_41),
.A2(n_42),
.B1(n_49),
.B2(n_50),
.Y(n_278)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_42),
.A2(n_240),
.B(n_245),
.Y(n_239)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_47),
.Y(n_272)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_48),
.Y(n_244)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.C(n_62),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_51),
.B(n_62),
.Y(n_149)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_56),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_56),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_57),
.B(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_61),
.Y(n_218)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_65),
.Y(n_318)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_65),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_88),
.B1(n_98),
.B2(n_99),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_67),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_67),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B(n_73),
.C(n_85),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_68),
.A2(n_70),
.B1(n_86),
.B2(n_87),
.Y(n_175)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_71),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_72),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_73),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.C(n_81),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_74),
.A2(n_81),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_74),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_74),
.A2(n_164),
.B1(n_251),
.B2(n_261),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_77),
.B(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_81),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_81),
.Y(n_252)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_97),
.Y(n_88)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_92),
.B(n_96),
.C(n_97),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_101),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_114),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_102),
.B(n_128),
.C(n_144),
.Y(n_184)
);

XNOR2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

MAJx2_ASAP7_75t_L g197 ( 
.A(n_103),
.B(n_107),
.C(n_111),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_110),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_111),
.A2(n_447),
.B1(n_448),
.B2(n_449),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_111),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_113),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_128),
.B1(n_144),
.B2(n_145),
.Y(n_114)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_116),
.B(n_120),
.C(n_127),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_117),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_117),
.B(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_125),
.B2(n_127),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_120),
.A2(n_121),
.B1(n_152),
.B2(n_153),
.Y(n_262)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_125),
.A2(n_127),
.B1(n_207),
.B2(n_211),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_125),
.B(n_347),
.Y(n_391)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_126),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_127),
.B(n_202),
.C(n_207),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_127),
.B(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.C(n_140),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_130),
.B1(n_140),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_136),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_135),
.A2(n_136),
.B1(n_320),
.B2(n_325),
.Y(n_319)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_136),
.B(n_316),
.C(n_325),
.Y(n_465)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_139),
.Y(n_401)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_146),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_168),
.C(n_173),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_147),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.C(n_156),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_148),
.B(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_150),
.A2(n_151),
.B1(n_156),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_164),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_157),
.A2(n_164),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_157),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_160),
.B(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_164),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_164),
.A2(n_207),
.B1(n_211),
.B2(n_261),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_164),
.B(n_211),
.C(n_310),
.Y(n_466)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_169),
.B(n_174),
.Y(n_275)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_177),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.C(n_180),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_200),
.B1(n_221),
.B2(n_222),
.Y(n_181)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_199),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_183),
.B(n_186),
.C(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_198),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_188),
.Y(n_198)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_188),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_197),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g298 ( 
.A(n_191),
.B(n_194),
.C(n_197),
.Y(n_298)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_195),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_195),
.B(n_305),
.C(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_200),
.B(n_221),
.C(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_212),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_201),
.B(n_213),
.C(n_214),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.Y(n_201)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_216),
.B(n_220),
.C(n_252),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_218),
.Y(n_367)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

OAI21x1_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_280),
.B(n_285),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_273),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g329 ( 
.A(n_225),
.B(n_273),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_253),
.C(n_257),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_226),
.B(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_238),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_227),
.B(n_239),
.C(n_249),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.C(n_235),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_228),
.B(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_229),
.A2(n_230),
.B1(n_235),
.B2(n_236),
.Y(n_337)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_249),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_253),
.A2(n_254),
.B1(n_257),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_257),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.C(n_263),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_258),
.B(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_262),
.B(n_263),
.Y(n_335)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.C(n_270),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_264),
.B(n_270),
.Y(n_373)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_267),
.B(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_269),
.Y(n_364)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx8_ASAP7_75t_L g450 ( 
.A(n_272),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_277),
.C(n_279),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NOR2x1_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_290),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_291),
.B(n_294),
.C(n_307),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_307),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_306),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_295),
.B(n_298),
.C(n_299),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

AO22x1_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_300),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_301),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_303),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_308),
.B(n_314),
.C(n_315),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_311),
.B(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_320),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_353),
.B(n_435),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_350),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_332),
.B(n_350),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.C(n_338),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_333),
.A2(n_334),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_336),
.B(n_338),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.C(n_346),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_339),
.A2(n_340),
.B1(n_341),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_339),
.Y(n_358)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_346),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_348),
.Y(n_428)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

AOI21x1_ASAP7_75t_SL g353 ( 
.A1(n_354),
.A2(n_377),
.B(n_434),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_374),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_355),
.B(n_374),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_359),
.C(n_372),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_372),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_365),
.C(n_368),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_360),
.B(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_368),
.Y(n_382)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI21x1_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_394),
.B(n_433),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_392),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_379),
.B(n_392),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.C(n_390),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_380),
.A2(n_381),
.B1(n_404),
.B2(n_406),
.Y(n_403)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_390),
.B1(n_391),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_383),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_384),
.A2(n_385),
.B1(n_386),
.B2(n_387),
.Y(n_397)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_407),
.B(n_432),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_403),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_396),
.B(n_403),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.C(n_402),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_416),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_398),
.A2(n_399),
.B1(n_402),
.B2(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_402),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_404),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_418),
.B(n_431),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_415),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_409),
.B(n_415),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_412),
.Y(n_424)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_419),
.A2(n_425),
.B(n_430),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_424),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_420),
.B(n_424),
.Y(n_430)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_429),
.Y(n_425)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_468),
.Y(n_436)
);

OR2x6_ASAP7_75t_SL g437 ( 
.A(n_438),
.B(n_467),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_438),
.B(n_467),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_458),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_456),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_451),
.B2(n_455),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_451),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_453),
.Y(n_452)
);

INVx8_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_464),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);


endmodule