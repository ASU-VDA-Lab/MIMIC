module fake_jpeg_21801_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_1),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_17),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_35),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_29),
.C(n_17),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_26),
.C(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_42),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_2),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_43),
.Y(n_46)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

NOR4xp25_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_22),
.C(n_11),
.D(n_13),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_27),
.A3(n_30),
.B1(n_15),
.B2(n_14),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_58),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_23),
.B1(n_18),
.B2(n_25),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_62),
.B1(n_30),
.B2(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_22),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_31),
.B(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_70),
.B(n_14),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_32),
.B(n_28),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_19),
.B1(n_23),
.B2(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_23),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_68),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_26),
.B(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_27),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_3),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_53),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_73),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_36),
.B1(n_33),
.B2(n_34),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_90),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_70),
.C(n_56),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_82),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_88),
.Y(n_105)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_15),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_38),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_91),
.A2(n_65),
.B(n_48),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_96),
.B(n_93),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_46),
.B(n_47),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_100),
.C(n_103),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_57),
.C(n_67),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_101),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_84),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_57),
.C(n_67),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_67),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_80),
.C(n_81),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_80),
.Y(n_118)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_118),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_74),
.B1(n_76),
.B2(n_71),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_108),
.B(n_105),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_108),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_81),
.C(n_86),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.C(n_121),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_81),
.C(n_86),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_87),
.C(n_89),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_96),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_64),
.B1(n_77),
.B2(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_124),
.B(n_125),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_61),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_104),
.B1(n_102),
.B2(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_136),
.C(n_137),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_109),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_120),
.C(n_119),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_108),
.C(n_111),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_115),
.B(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_139),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_126),
.CI(n_113),
.CON(n_139),
.SN(n_139)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_142),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_116),
.C(n_117),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_132),
.Y(n_149)
);

AO221x1_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_83),
.B1(n_112),
.B2(n_77),
.C(n_64),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_145),
.B(n_127),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_146),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_151),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_135),
.A3(n_139),
.B1(n_132),
.B2(n_136),
.C1(n_141),
.C2(n_142),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_156),
.B(n_157),
.Y(n_158)
);

NAND4xp25_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_3),
.C(n_6),
.D(n_7),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_150),
.A2(n_146),
.B1(n_140),
.B2(n_8),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_9),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.C1(n_6),
.C2(n_7),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_152),
.B(n_6),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_154),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_156),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_158),
.Y(n_164)
);


endmodule