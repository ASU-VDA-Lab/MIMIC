module fake_netlist_1_5312_n_32 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2xp33_ASAP7_75t_L g12 ( .A(n_0), .B(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_10), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_11), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_4), .B(n_5), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
A2O1A1Ixp33_ASAP7_75t_L g18 ( .A1(n_14), .A2(n_0), .B(n_1), .C(n_2), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_14), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
AOI22xp33_ASAP7_75t_SL g21 ( .A1(n_20), .A2(n_16), .B1(n_13), .B2(n_12), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
BUFx10_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
NAND3xp33_ASAP7_75t_SL g26 ( .A(n_24), .B(n_18), .C(n_13), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
XNOR2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_23), .Y(n_28) );
NAND2xp33_ASAP7_75t_R g29 ( .A(n_28), .B(n_1), .Y(n_29) );
AND4x1_ASAP7_75t_L g30 ( .A(n_27), .B(n_18), .C(n_3), .D(n_4), .Y(n_30) );
AOI22xp5_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_2), .B1(n_5), .B2(n_15), .Y(n_31) );
AOI22xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_30), .B1(n_7), .B2(n_9), .Y(n_32) );
endmodule