module fake_jpeg_16356_n_303 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_288;
wire n_284;
wire n_272;
wire n_234;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_11),
.B(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx2_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12f_ASAP7_75t_SL g40 ( 
.A(n_20),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_40),
.B(n_39),
.Y(n_88)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_2),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_48),
.B(n_58),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_59),
.Y(n_81)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_62),
.Y(n_89)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_2),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_24),
.B(n_0),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_30),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_69),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_14),
.B(n_5),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_0),
.C(n_1),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_15),
.C(n_26),
.Y(n_107)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_75),
.B(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_30),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_83),
.B(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_23),
.B1(n_31),
.B2(n_14),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_87),
.A2(n_93),
.B1(n_102),
.B2(n_104),
.Y(n_143)
);

OR2x2_ASAP7_75t_SL g152 ( 
.A(n_88),
.B(n_109),
.Y(n_152)
);

CKINVDCx12_ASAP7_75t_R g92 ( 
.A(n_40),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_99),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_31),
.B1(n_23),
.B2(n_26),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_37),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_SL g97 ( 
.A(n_44),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_54),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_37),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_101),
.B(n_106),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_35),
.B1(n_21),
.B2(n_29),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_55),
.A2(n_29),
.B1(n_21),
.B2(n_34),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_50),
.B(n_34),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_46),
.B(n_15),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_47),
.B(n_17),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_41),
.A2(n_71),
.B1(n_49),
.B2(n_57),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_63),
.B(n_67),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_60),
.A2(n_9),
.A3(n_10),
.B1(n_12),
.B2(n_0),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_63),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_51),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_119)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_56),
.B(n_12),
.Y(n_120)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_88),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_122),
.A2(n_123),
.B(n_150),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_66),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_79),
.C(n_85),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_125),
.A2(n_74),
.B1(n_100),
.B2(n_94),
.Y(n_180)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_68),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_128),
.B(n_142),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_133),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_134),
.Y(n_173)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_80),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_146),
.Y(n_169)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g141 ( 
.A(n_105),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_141),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_101),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_91),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_144),
.B(n_148),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_104),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_108),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_81),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_154),
.Y(n_170)
);

OR2x4_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_119),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_157),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_84),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_86),
.B(n_74),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_159),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_116),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_130),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_79),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_117),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_177),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_162),
.A2(n_117),
.B1(n_105),
.B2(n_98),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_187),
.B1(n_188),
.B2(n_193),
.Y(n_200)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_157),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_85),
.B1(n_94),
.B2(n_95),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_185),
.B1(n_160),
.B2(n_140),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_103),
.B1(n_123),
.B2(n_150),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_125),
.A2(n_103),
.B1(n_151),
.B2(n_145),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_143),
.A2(n_129),
.B1(n_153),
.B2(n_126),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_196),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_191),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_124),
.B(n_129),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_134),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_143),
.A2(n_129),
.B1(n_152),
.B2(n_124),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g195 ( 
.A1(n_131),
.A2(n_155),
.A3(n_152),
.B1(n_121),
.B2(n_127),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_130),
.A3(n_149),
.B1(n_175),
.B2(n_163),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_199),
.A2(n_206),
.B1(n_183),
.B2(n_215),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_205),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_215),
.B(n_217),
.Y(n_229)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_207),
.B(n_211),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_137),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_210),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_163),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_218),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_171),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_164),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_220),
.A2(n_183),
.B1(n_190),
.B2(n_173),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_166),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_222),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_224),
.B(n_240),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_174),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_235),
.C(n_200),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_182),
.B1(n_173),
.B2(n_176),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_243),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_215),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_230),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_196),
.B(n_184),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_203),
.B(n_209),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_179),
.B1(n_177),
.B2(n_166),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_184),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_236),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_229),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_255),
.C(n_259),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_249),
.Y(n_269)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_221),
.B(n_206),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_252),
.A2(n_257),
.B1(n_217),
.B2(n_239),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_208),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_200),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_256),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_244),
.B(n_238),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_201),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_232),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

AO221x1_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_202),
.B1(n_205),
.B2(n_225),
.C(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_241),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_248),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_259),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_227),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_255),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_217),
.B1(n_241),
.B2(n_206),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_253),
.B1(n_257),
.B2(n_245),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_252),
.B(n_253),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_272),
.B(n_248),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_239),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_246),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_277),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_270),
.B(n_269),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_281),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_280),
.A2(n_271),
.B(n_260),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_246),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_280),
.B(n_268),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_279),
.A2(n_251),
.B1(n_256),
.B2(n_264),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_286),
.A2(n_279),
.B1(n_249),
.B2(n_242),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_242),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_292),
.C(n_293),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_288),
.A2(n_263),
.A3(n_266),
.B1(n_281),
.B2(n_282),
.C1(n_273),
.C2(n_249),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_295),
.B(n_289),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_273),
.B1(n_234),
.B2(n_204),
.Y(n_295)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_234),
.C(n_287),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_297),
.A2(n_285),
.B(n_290),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_SL g301 ( 
.A1(n_300),
.A2(n_298),
.B(n_233),
.C(n_212),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_299),
.B1(n_198),
.B2(n_219),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_179),
.Y(n_303)
);


endmodule