module real_jpeg_4419_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_0),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_0),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_0),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_0),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_0),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_0),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_0),
.B(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_1),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_2),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_2),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_2),
.B(n_229),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_2),
.B(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_2),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_2),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_2),
.B(n_126),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_3),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_3),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_3),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_4),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_4),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_4),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_5),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_5),
.Y(n_191)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_5),
.Y(n_223)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_5),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_6),
.B(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_6),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_6),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_6),
.B(n_300),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_6),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_6),
.B(n_42),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_6),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_6),
.B(n_400),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_7),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_7),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_7),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_7),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_7),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_7),
.B(n_229),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_7),
.B(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_7),
.B(n_231),
.Y(n_401)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_8),
.Y(n_129)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_9),
.Y(n_488)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_10),
.Y(n_284)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_12),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_12),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_12),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_12),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_12),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_12),
.B(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_13),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_13),
.Y(n_316)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_15),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_15),
.B(n_105),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_15),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_15),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_15),
.B(n_124),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_15),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_15),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_16),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_16),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_16),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_16),
.B(n_226),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_16),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_16),
.B(n_361),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_17),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_17),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_17),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_17),
.B(n_117),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_17),
.B(n_318),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_17),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_17),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_18),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_18),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_18),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_18),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_18),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g277 ( 
.A(n_18),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_18),
.B(n_361),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_18),
.B(n_408),
.Y(n_407)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_486),
.B(n_489),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_193),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_192),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_159),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_25),
.B(n_159),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_118),
.B2(n_158),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_82),
.C(n_99),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_28),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_50),
.C(n_68),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_29),
.B(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_30),
.B(n_38),
.C(n_44),
.Y(n_130)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_34),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_35),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_44),
.B2(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_37),
.A2(n_38),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_37),
.B(n_122),
.C(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_43),
.Y(n_278)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_43),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_44),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_44),
.B(n_102),
.C(n_106),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_44),
.A2(n_49),
.B1(n_106),
.B2(n_107),
.Y(n_168)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_48),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_50),
.B(n_68),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.C(n_61),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_51),
.B(n_61),
.Y(n_175)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_53),
.Y(n_213)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_53),
.Y(n_346)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_54),
.Y(n_153)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_55),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_56),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_60),
.Y(n_232)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_65),
.Y(n_210)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_65),
.Y(n_403)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_67),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_67),
.Y(n_328)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_67),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g492 ( 
.A(n_68),
.Y(n_492)
);

FAx1_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_75),
.CI(n_79),
.CON(n_68),
.SN(n_68)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_69),
.B(n_75),
.C(n_79),
.Y(n_131)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx8_ASAP7_75t_L g400 ( 
.A(n_73),
.Y(n_400)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_74),
.Y(n_381)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_78),
.Y(n_281)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_82),
.A2(n_99),
.B1(n_100),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_83),
.B(n_89),
.C(n_98),
.Y(n_142)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_94),
.B2(n_98),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_97),
.Y(n_260)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.C(n_115),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_101),
.B(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_102),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_106),
.A2(n_107),
.B1(n_171),
.B2(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_107),
.B(n_170),
.C(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_109),
.A2(n_110),
.B1(n_115),
.B2(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_115),
.A2(n_116),
.B1(n_189),
.B2(n_190),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_179),
.C(n_189),
.Y(n_178)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_117),
.Y(n_235)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_132),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_130),
.C(n_131),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_123),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_129),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_131),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_143),
.B2(n_157),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_155),
.B2(n_156),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_149),
.B1(n_150),
.B2(n_154),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_160),
.B(n_163),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_165),
.B(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_176),
.C(n_178),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_166),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.C(n_174),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_167),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_169),
.B(n_174),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_215),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_171),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_173),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_173),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_176),
.B(n_178),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.C(n_186),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_186),
.Y(n_201)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_188),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AO21x1_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_479),
.B(n_484),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_286),
.B(n_478),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_241),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_197),
.B(n_241),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_236),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_198),
.B(n_237),
.C(n_239),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_217),
.C(n_219),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_199),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.C(n_214),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_200),
.B(n_464),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_202),
.A2(n_203),
.B1(n_214),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.C(n_211),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_204),
.B(n_211),
.Y(n_454)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_207),
.B(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_214),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_219),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.C(n_233),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.C(n_228),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_221),
.B(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_228),
.Y(n_253)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_230),
.B(n_233),
.Y(n_270)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_248),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_243),
.B(n_246),
.Y(n_474)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_248),
.B(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_268),
.C(n_271),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_250),
.B(n_467),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_261),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_251),
.A2(n_252),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_254),
.A2(n_255),
.B(n_257),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_254),
.B(n_261),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.C(n_266),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_422)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_266),
.B(n_422),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_267),
.B(n_358),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_268),
.A2(n_269),
.B1(n_271),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_271),
.Y(n_468)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_282),
.C(n_285),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_273),
.B(n_456),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.C(n_279),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_274),
.B(n_434),
.Y(n_433)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_277),
.A2(n_279),
.B1(n_280),
.B2(n_435),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_277),
.Y(n_435)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_282),
.B(n_285),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_284),
.Y(n_358)
);

AOI21x1_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_472),
.B(n_477),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_459),
.B(n_471),
.Y(n_287)
);

AOI21x1_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_441),
.B(n_458),
.Y(n_288)
);

OAI21x1_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_415),
.B(n_440),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_385),
.B(n_414),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_350),
.B(n_384),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_330),
.B(n_349),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_307),
.B(n_329),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_304),
.B(n_306),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_302),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_302),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_299),
.Y(n_308)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_309),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_320),
.B2(n_321),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_323),
.C(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_317),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_348),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_348),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_340),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_339),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_339),
.C(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_338),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_338),
.Y(n_355)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_340),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_368),
.C(n_369),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_347),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_347),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_351),
.B(n_353),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_366),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_354),
.B(n_367),
.C(n_370),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_357),
.C(n_359),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_362),
.B1(n_363),
.B2(n_365),
.Y(n_359)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_360),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_365),
.Y(n_395)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_SL g409 ( 
.A(n_364),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_375),
.Y(n_370)
);

MAJx2_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_379),
.C(n_382),
.Y(n_412)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_379),
.B1(n_382),
.B2(n_383),
.Y(n_375)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_376),
.Y(n_382)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_378),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_379),
.Y(n_383)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_413),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_413),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_397),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_396),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_396),
.C(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_395),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.Y(n_389)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_429),
.C(n_430),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_397),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_404),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_398),
.B(n_406),
.C(n_411),
.Y(n_418)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_398),
.Y(n_494)
);

FAx1_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_401),
.CI(n_402),
.CON(n_398),
.SN(n_398)
);

MAJx2_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_401),
.C(n_402),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_406),
.B1(n_411),
.B2(n_412),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_410),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_410),
.Y(n_425)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_438),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_438),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_427),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_419),
.C(n_427),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_423),
.B2(n_424),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_450),
.C(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_425),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_431),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_432),
.C(n_437),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_433),
.B1(n_436),
.B2(n_437),
.Y(n_431)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_432),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_433),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_457),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_457),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_448),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_447),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_447),
.C(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_445),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_452),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_449),
.B(n_453),
.C(n_455),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_469),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_460),
.B(n_469),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_461),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_466),
.C(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_473),
.B(n_475),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_475),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_483),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_483),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx13_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_488),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);


endmodule