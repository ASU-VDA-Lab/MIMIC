module fake_jpeg_27683_n_297 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_297);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_297;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_24),
.B1(n_22),
.B2(n_27),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_50),
.B1(n_34),
.B2(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_45),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_51),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_25),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_38),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_24),
.B1(n_22),
.B2(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_59),
.B(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_67),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_87),
.B1(n_29),
.B2(n_28),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_84),
.Y(n_112)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_82),
.Y(n_103)
);

AOI32xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_45),
.A3(n_37),
.B1(n_26),
.B2(n_40),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_83),
.B(n_85),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_17),
.B1(n_21),
.B2(n_18),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_80),
.A2(n_29),
.B1(n_28),
.B2(n_30),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_35),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_100),
.Y(n_129)
);

XOR2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_26),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_26),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_30),
.B(n_32),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_31),
.B(n_33),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_102),
.B1(n_108),
.B2(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_19),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_77),
.B1(n_33),
.B2(n_21),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_71),
.A2(n_16),
.B1(n_32),
.B2(n_31),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_16),
.B1(n_31),
.B2(n_29),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_131),
.B1(n_92),
.B2(n_91),
.Y(n_149)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_57),
.B1(n_68),
.B2(n_67),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_118),
.A2(n_125),
.B1(n_127),
.B2(n_134),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_65),
.B1(n_67),
.B2(n_87),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_119),
.A2(n_141),
.B1(n_94),
.B2(n_110),
.Y(n_157)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_124),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_128),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_67),
.B(n_65),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_92),
.B1(n_91),
.B2(n_88),
.Y(n_144)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_76),
.B1(n_84),
.B2(n_82),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_61),
.B1(n_77),
.B2(n_64),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_98),
.B(n_107),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_128),
.B(n_123),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_86),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_138),
.Y(n_150)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_0),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_40),
.B1(n_17),
.B2(n_21),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_136),
.C(n_114),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_105),
.C(n_100),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_21),
.B1(n_17),
.B2(n_26),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_112),
.B(n_26),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_89),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_97),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_101),
.A2(n_88),
.B1(n_114),
.B2(n_106),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_19),
.B1(n_25),
.B2(n_20),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_144),
.A2(n_153),
.B(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_162),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_131),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_166),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_157),
.B1(n_133),
.B2(n_117),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_118),
.A2(n_124),
.B1(n_139),
.B2(n_143),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_94),
.B1(n_110),
.B2(n_2),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_160),
.B1(n_165),
.B2(n_5),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_25),
.C(n_18),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_164),
.C(n_134),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_19),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_25),
.C(n_19),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_120),
.A2(n_25),
.B1(n_20),
.B2(n_9),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_169),
.B1(n_137),
.B2(n_138),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_123),
.A2(n_20),
.B1(n_8),
.B2(n_9),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_0),
.Y(n_192)
);

AO22x1_ASAP7_75t_SL g173 ( 
.A1(n_123),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_173)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_135),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_188),
.C(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_195),
.B1(n_201),
.B2(n_152),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_130),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_184),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_193),
.B1(n_199),
.B2(n_169),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_191),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_186),
.A2(n_146),
.B(n_167),
.Y(n_208)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_192),
.Y(n_213)
);

AOI22x1_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_146),
.B(n_8),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_15),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_11),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_197),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_155),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_11),
.B1(n_13),
.B2(n_7),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_154),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_207),
.A2(n_219),
.B1(n_193),
.B2(n_194),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_211),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_163),
.B1(n_171),
.B2(n_170),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_216),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_163),
.B1(n_145),
.B2(n_152),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_150),
.B1(n_165),
.B2(n_173),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_221),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_144),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_200),
.B(n_189),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_144),
.B1(n_172),
.B2(n_173),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_150),
.B1(n_162),
.B2(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_192),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_187),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_176),
.C(n_188),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_220),
.C(n_196),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_214),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_227),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_222),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_180),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_228),
.B(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_233),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_175),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_209),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_200),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_186),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_215),
.B1(n_211),
.B2(n_195),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_240),
.A2(n_223),
.B1(n_187),
.B2(n_220),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_177),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_208),
.Y(n_249)
);

AOI21x1_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_218),
.B(n_209),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_249),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_218),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_253),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_219),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_207),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_238),
.C(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_235),
.B1(n_238),
.B2(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_261),
.B1(n_242),
.B2(n_232),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_265),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_235),
.B1(n_226),
.B2(n_240),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_237),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_246),
.A2(n_178),
.B1(n_232),
.B2(n_211),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_250),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_254),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_271),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_252),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_276),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_253),
.C(n_251),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_274),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_SL g275 ( 
.A(n_267),
.B(n_248),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_258),
.B(n_265),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_264),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_10),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_277),
.B(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_191),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_259),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_270),
.B(n_272),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_285),
.B(n_288),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_287),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_282),
.A2(n_273),
.B1(n_259),
.B2(n_7),
.Y(n_287)
);

A2O1A1O1Ixp25_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_282),
.B(n_278),
.C(n_10),
.D(n_12),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_289),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_290),
.C(n_12),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_293),
.B(n_13),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_15),
.C(n_5),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_6),
.C(n_15),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_6),
.Y(n_297)
);


endmodule