module fake_jpeg_16975_n_302 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_36),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_25),
.B1(n_32),
.B2(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_32),
.B1(n_18),
.B2(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_17),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_33),
.B1(n_40),
.B2(n_32),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_43),
.B1(n_18),
.B2(n_32),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_23),
.B1(n_47),
.B2(n_28),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_71),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_35),
.CI(n_40),
.CON(n_68),
.SN(n_68)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_68),
.B(n_35),
.Y(n_102)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_44),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_83),
.B(n_71),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_79),
.B1(n_81),
.B2(n_26),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_24),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_17),
.B1(n_20),
.B2(n_28),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_23),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_23),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_97),
.B(n_113),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_33),
.B1(n_57),
.B2(n_58),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_105),
.B1(n_78),
.B2(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_52),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_90),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_93),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_66),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_94),
.A2(n_78),
.B1(n_44),
.B2(n_33),
.Y(n_131)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_35),
.C(n_41),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_101),
.C(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_35),
.C(n_49),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_112),
.Y(n_126)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_35),
.C(n_49),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_24),
.B1(n_26),
.B2(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_111),
.Y(n_136)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_83),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_23),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_125),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_80),
.B1(n_85),
.B2(n_76),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_119),
.B1(n_122),
.B2(n_135),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_88),
.A2(n_70),
.B1(n_72),
.B2(n_20),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_124),
.B1(n_131),
.B2(n_113),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_83),
.B1(n_85),
.B2(n_76),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_68),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_129),
.C(n_139),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_89),
.A2(n_70),
.B1(n_72),
.B2(n_17),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_68),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_86),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_138),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_60),
.B1(n_62),
.B2(n_33),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_52),
.B1(n_84),
.B2(n_59),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_35),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_21),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_167),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_107),
.B1(n_108),
.B2(n_113),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_148),
.B1(n_149),
.B2(n_165),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_123),
.C(n_129),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_154),
.C(n_157),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_101),
.B1(n_98),
.B2(n_91),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_103),
.B1(n_91),
.B2(n_92),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_151),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_156),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_109),
.C(n_96),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_100),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_162),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_110),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_0),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_164),
.B(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_30),
.B(n_21),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_96),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_163),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_30),
.B(n_29),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_29),
.B1(n_30),
.B2(n_12),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_125),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_169),
.B(n_186),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_170),
.A2(n_185),
.B(n_164),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_117),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_179),
.C(n_180),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_173),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_176),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_165),
.B1(n_141),
.B2(n_161),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_114),
.C(n_69),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_118),
.Y(n_180)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_21),
.A3(n_27),
.B1(n_22),
.B2(n_69),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_38),
.Y(n_210)
);

INVxp33_ASAP7_75t_SL g185 ( 
.A(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_27),
.Y(n_186)
);

BUFx2_ASAP7_75t_SL g192 ( 
.A(n_146),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_158),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_154),
.C(n_157),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_198),
.C(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_148),
.C(n_160),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_145),
.C(n_152),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_175),
.A2(n_156),
.B1(n_144),
.B2(n_162),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_204),
.B1(n_207),
.B2(n_216),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_215),
.B(n_217),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_143),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_205),
.C(n_206),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_188),
.B1(n_173),
.B2(n_179),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_149),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_163),
.C(n_140),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_158),
.B1(n_150),
.B2(n_11),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_69),
.C(n_27),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_212),
.C(n_213),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_38),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_38),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_21),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_182),
.B1(n_191),
.B2(n_183),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_186),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_222),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_221),
.B(n_226),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_189),
.B(n_193),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_170),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_187),
.C(n_184),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_234),
.C(n_194),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_183),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_233),
.Y(n_238)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_178),
.C(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_237),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_203),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_223),
.B1(n_227),
.B2(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_244),
.C(n_247),
.Y(n_253)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_206),
.C(n_212),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_11),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_210),
.C(n_27),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_229),
.B(n_8),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_248),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_231),
.B1(n_234),
.B2(n_224),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_8),
.B1(n_15),
.B2(n_13),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_228),
.A2(n_13),
.B(n_12),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_13),
.Y(n_265)
);

AOI21x1_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_249),
.B(n_241),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_265),
.B(n_10),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_224),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_260),
.C(n_262),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_222),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_238),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_2),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_230),
.C(n_236),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_246),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_270),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_247),
.C(n_243),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_262),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_252),
.B1(n_3),
.B2(n_4),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_269),
.A2(n_272),
.B1(n_276),
.B2(n_273),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_275),
.B(n_6),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_256),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_4),
.B(n_5),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_4),
.B(n_5),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_5),
.B(n_6),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_258),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_278),
.B(n_279),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_254),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_253),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_282),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_257),
.B(n_7),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_285),
.A2(n_6),
.B(n_7),
.C(n_268),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_291),
.B(n_292),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_280),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_266),
.B(n_267),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_266),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_295),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_6),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_286),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_296),
.A2(n_288),
.B(n_7),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_297),
.B1(n_21),
.B2(n_38),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_38),
.Y(n_300)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_300),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_38),
.Y(n_302)
);


endmodule