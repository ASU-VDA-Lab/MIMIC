module fake_netlist_6_4365_n_2208 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_2208);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2208;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_907;
wire n_1446;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_824;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_1843;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_2101;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_697;
wire n_890;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_1765;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_2069;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1951;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_956;
wire n_960;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_2016;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_1270;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_1667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2200;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_962;
wire n_1041;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_1222;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_879;
wire n_959;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2154;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1373;
wire n_1292;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_1678;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_1170;
wire n_1629;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2116;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1612;
wire n_1240;

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_116),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_642),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_665),
.Y(n_695)
);

BUFx5_ASAP7_75t_L g696 ( 
.A(n_243),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_417),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_393),
.Y(n_698)
);

CKINVDCx16_ASAP7_75t_R g699 ( 
.A(n_565),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_35),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_335),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_128),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_539),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_92),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_635),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_667),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_277),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_334),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_20),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_196),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_641),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_367),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_436),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_458),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_620),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_581),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_202),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_636),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_604),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_646),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_657),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_655),
.Y(n_722)
);

CKINVDCx20_ASAP7_75t_R g723 ( 
.A(n_612),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_652),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_597),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_378),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_543),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_640),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_605),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_663),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_149),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_174),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_297),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_593),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_633),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_625),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_638),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_84),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_282),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_586),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_388),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_649),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_256),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_618),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_402),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_587),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_584),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_13),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_131),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_266),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_384),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_606),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_204),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_221),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_227),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_329),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_217),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_510),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_181),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_32),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_566),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_576),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_595),
.Y(n_763)
);

BUFx10_ASAP7_75t_L g764 ( 
.A(n_656),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_421),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_481),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_127),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_639),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_634),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_219),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_574),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_564),
.Y(n_772)
);

BUFx2_ASAP7_75t_SL g773 ( 
.A(n_648),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_598),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_632),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_216),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_209),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_589),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_112),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_591),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_644),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_18),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_619),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_689),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_659),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_508),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_178),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_590),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_600),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_658),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_452),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_19),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_107),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_37),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_60),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_88),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_76),
.Y(n_797)
);

CKINVDCx16_ASAP7_75t_R g798 ( 
.A(n_575),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_439),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_446),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_650),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_346),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_666),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_553),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_611),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_503),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_447),
.Y(n_807)
);

CKINVDCx16_ASAP7_75t_R g808 ( 
.A(n_582),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_499),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_32),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_501),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_563),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_52),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_373),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_171),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_261),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_214),
.Y(n_817)
);

CKINVDCx16_ASAP7_75t_R g818 ( 
.A(n_181),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_637),
.Y(n_819)
);

CKINVDCx16_ASAP7_75t_R g820 ( 
.A(n_427),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_399),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_10),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_408),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_616),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_614),
.Y(n_825)
);

INVxp33_ASAP7_75t_R g826 ( 
.A(n_471),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_187),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_493),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_505),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_71),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_49),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_613),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_592),
.Y(n_833)
);

BUFx10_ASAP7_75t_L g834 ( 
.A(n_470),
.Y(n_834)
);

CKINVDCx16_ASAP7_75t_R g835 ( 
.A(n_607),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_201),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_186),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_429),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_496),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_599),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_536),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_621),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_573),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_257),
.Y(n_844)
);

BUFx5_ASAP7_75t_L g845 ( 
.A(n_74),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_480),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_434),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_561),
.Y(n_848)
);

CKINVDCx16_ASAP7_75t_R g849 ( 
.A(n_654),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_643),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_661),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_38),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_630),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_622),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_428),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_424),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_178),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_603),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_522),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_671),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_594),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_285),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_175),
.Y(n_863)
);

BUFx5_ASAP7_75t_L g864 ( 
.A(n_500),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_372),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_347),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_631),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_114),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_380),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_80),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_664),
.Y(n_871)
);

BUFx5_ASAP7_75t_L g872 ( 
.A(n_438),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_492),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_645),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_624),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_363),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_487),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_265),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_577),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_125),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_610),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_601),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_98),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_407),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_628),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_662),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_660),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_141),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_546),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_544),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_440),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_415),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_362),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_43),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_52),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_426),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_216),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_99),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_596),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_530),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_580),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_268),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_413),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_484),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_552),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_545),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_64),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_219),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_670),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_617),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_163),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_627),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_401),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_623),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_571),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_588),
.Y(n_916)
);

BUFx2_ASAP7_75t_SL g917 ( 
.A(n_579),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_228),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_262),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_158),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_122),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_337),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_158),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_668),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_247),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_228),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_684),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_531),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_629),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_653),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_329),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_524),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_687),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_651),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_609),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_669),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_182),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_159),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_475),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_585),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_677),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_244),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_148),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_283),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_615),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_83),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_147),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_491),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_578),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_680),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_81),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_231),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_263),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_271),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_672),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_608),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_210),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_420),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_626),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_583),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_443),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_55),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_331),
.Y(n_963)
);

BUFx5_ASAP7_75t_L g964 ( 
.A(n_312),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_99),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_65),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_279),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_122),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_567),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_602),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_647),
.Y(n_971)
);

BUFx2_ASAP7_75t_SL g972 ( 
.A(n_694),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_698),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_696),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_795),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_696),
.Y(n_976)
);

INVxp33_ASAP7_75t_SL g977 ( 
.A(n_794),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_703),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_790),
.B(n_1),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_715),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_711),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_827),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_696),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_713),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_696),
.Y(n_985)
);

CKINVDCx14_ASAP7_75t_R g986 ( 
.A(n_862),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_696),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_716),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_845),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_718),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_719),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_722),
.Y(n_992)
);

CKINVDCx20_ASAP7_75t_R g993 ( 
.A(n_723),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_740),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_724),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_845),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_845),
.Y(n_997)
);

INVxp67_ASAP7_75t_SL g998 ( 
.A(n_875),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_725),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_845),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_982),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_982),
.Y(n_1002)
);

NAND2x1p5_ASAP7_75t_L g1003 ( 
.A(n_979),
.B(n_799),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_1000),
.Y(n_1004)
);

NAND2xp33_ASAP7_75t_SL g1005 ( 
.A(n_975),
.B(n_827),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_986),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_974),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_973),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_976),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_983),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_985),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_987),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_978),
.B(n_828),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_975),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_989),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_977),
.B(n_699),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_998),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_981),
.B(n_901),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_984),
.B(n_960),
.Y(n_1019)
);

AND2x6_ASAP7_75t_L g1020 ( 
.A(n_996),
.B(n_842),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_997),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_988),
.B(n_806),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_990),
.B(n_856),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_991),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_SL g1025 ( 
.A1(n_980),
.A2(n_754),
.B1(n_810),
.B2(n_749),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_992),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_995),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_999),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_SL g1029 ( 
.A(n_972),
.B(n_798),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_993),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_1024),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1015),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_1015),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1007),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_1021),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1009),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_1027),
.B(n_758),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_1004),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_1014),
.Y(n_1039)
);

AND2x2_ASAP7_75t_SL g1040 ( 
.A(n_1029),
.B(n_693),
.Y(n_1040)
);

INVx3_ASAP7_75t_SL g1041 ( 
.A(n_1024),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_1010),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1011),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1012),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_1019),
.B(n_808),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_1023),
.B(n_820),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1017),
.B(n_818),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1001),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1022),
.B(n_701),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_1013),
.B(n_835),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_1026),
.B(n_763),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_1008),
.B(n_1028),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1002),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_1006),
.B(n_778),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1020),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1020),
.Y(n_1056)
);

INVxp33_ASAP7_75t_L g1057 ( 
.A(n_1025),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1018),
.B(n_812),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_1020),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1005),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1003),
.B(n_849),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_1030),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_1016),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1027),
.B(n_879),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1007),
.B(n_777),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_1024),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1004),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_1024),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_1015),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_1023),
.Y(n_1070)
);

CKINVDCx6p67_ASAP7_75t_R g1071 ( 
.A(n_1006),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1019),
.B(n_994),
.Y(n_1072)
);

OAI221xp5_ASAP7_75t_L g1073 ( 
.A1(n_1050),
.A2(n_831),
.B1(n_837),
.B2(n_815),
.C(n_753),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1041),
.B(n_1049),
.Y(n_1074)
);

AO22x2_ASAP7_75t_L g1075 ( 
.A1(n_1046),
.A2(n_946),
.B1(n_866),
.B2(n_863),
.Y(n_1075)
);

AND2x6_ASAP7_75t_L g1076 ( 
.A(n_1056),
.B(n_695),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1034),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1045),
.B(n_705),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_1068),
.B(n_824),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1058),
.A2(n_903),
.B1(n_932),
.B2(n_900),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1034),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1036),
.B(n_706),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_1039),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_1049),
.Y(n_1084)
);

AO22x2_ASAP7_75t_L g1085 ( 
.A1(n_1047),
.A2(n_702),
.B1(n_739),
.B2(n_731),
.Y(n_1085)
);

OAI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_1043),
.A2(n_966),
.B1(n_732),
.B2(n_738),
.C(n_709),
.Y(n_1086)
);

AO22x2_ASAP7_75t_L g1087 ( 
.A1(n_1047),
.A2(n_802),
.B1(n_743),
.B2(n_748),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_1071),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1044),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1067),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_1031),
.B(n_1069),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1038),
.B(n_714),
.Y(n_1092)
);

AO22x2_ASAP7_75t_L g1093 ( 
.A1(n_1060),
.A2(n_792),
.B1(n_793),
.B2(n_787),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_1065),
.Y(n_1094)
);

BUFx8_ASAP7_75t_L g1095 ( 
.A(n_1054),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1038),
.B(n_720),
.Y(n_1096)
);

AO22x2_ASAP7_75t_L g1097 ( 
.A1(n_1061),
.A2(n_830),
.B1(n_893),
.B2(n_868),
.Y(n_1097)
);

AO22x2_ASAP7_75t_L g1098 ( 
.A1(n_1057),
.A2(n_925),
.B1(n_926),
.B2(n_920),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_1065),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1048),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1053),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_1051),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1042),
.Y(n_1103)
);

NAND2x1p5_ASAP7_75t_L g1104 ( 
.A(n_1033),
.B(n_912),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1035),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1040),
.B(n_940),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1035),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1032),
.Y(n_1108)
);

AO22x2_ASAP7_75t_L g1109 ( 
.A1(n_1070),
.A2(n_943),
.B1(n_947),
.B2(n_942),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1072),
.B(n_721),
.Y(n_1110)
);

OAI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_1063),
.A2(n_962),
.B1(n_918),
.B2(n_954),
.C(n_796),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1033),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1069),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1037),
.A2(n_869),
.B1(n_729),
.B2(n_734),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1062),
.B(n_923),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1055),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1056),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1064),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1052),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_1059),
.B(n_697),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1034),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1067),
.Y(n_1122)
);

BUFx8_ASAP7_75t_L g1123 ( 
.A(n_1054),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1034),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1039),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1045),
.B(n_727),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_1041),
.Y(n_1127)
);

OAI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1050),
.A2(n_708),
.B1(n_969),
.B2(n_882),
.C(n_769),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1050),
.A2(n_728),
.B1(n_730),
.B2(n_726),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1067),
.Y(n_1130)
);

OAI221xp5_ASAP7_75t_L g1131 ( 
.A1(n_1050),
.A2(n_877),
.B1(n_927),
.B2(n_811),
.C(n_765),
.Y(n_1131)
);

AO22x2_ASAP7_75t_L g1132 ( 
.A1(n_1046),
.A2(n_826),
.B1(n_768),
.B2(n_771),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1034),
.Y(n_1133)
);

BUFx8_ASAP7_75t_L g1134 ( 
.A(n_1054),
.Y(n_1134)
);

AND2x2_ASAP7_75t_SL g1135 ( 
.A(n_1040),
.B(n_827),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1034),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1054),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1034),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_SL g1139 ( 
.A(n_1041),
.B(n_844),
.Y(n_1139)
);

AO22x2_ASAP7_75t_L g1140 ( 
.A1(n_1046),
.A2(n_783),
.B1(n_788),
.B2(n_735),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1050),
.A2(n_774),
.B1(n_784),
.B2(n_736),
.Y(n_1141)
);

AND2x4_ASAP7_75t_L g1142 ( 
.A(n_1031),
.B(n_801),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1050),
.B(n_700),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1045),
.B(n_803),
.Y(n_1144)
);

NAND2x1p5_ASAP7_75t_L g1145 ( 
.A(n_1066),
.B(n_814),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1045),
.B(n_821),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1045),
.B(n_829),
.Y(n_1147)
);

AO22x2_ASAP7_75t_L g1148 ( 
.A1(n_1046),
.A2(n_838),
.B1(n_841),
.B2(n_839),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1034),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1041),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_1039),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1034),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1039),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1045),
.B(n_847),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1045),
.B(n_850),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1034),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1041),
.B(n_878),
.Y(n_1157)
);

AO22x2_ASAP7_75t_L g1158 ( 
.A1(n_1046),
.A2(n_855),
.B1(n_860),
.B2(n_859),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1034),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1045),
.B(n_867),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1067),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1067),
.Y(n_1162)
);

AO22x2_ASAP7_75t_L g1163 ( 
.A1(n_1046),
.A2(n_873),
.B1(n_889),
.B2(n_874),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1034),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1050),
.A2(n_741),
.B1(n_742),
.B2(n_737),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1034),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1034),
.Y(n_1167)
);

NAND2x1p5_ASAP7_75t_L g1168 ( 
.A(n_1066),
.B(n_892),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1034),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1050),
.A2(n_745),
.B1(n_746),
.B2(n_744),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1135),
.B(n_747),
.Y(n_1171)
);

NAND2xp33_ASAP7_75t_SL g1172 ( 
.A(n_1150),
.B(n_883),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1083),
.B(n_751),
.Y(n_1173)
);

NAND2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1127),
.B(n_1119),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1105),
.B(n_899),
.Y(n_1175)
);

NAND2xp33_ASAP7_75t_SL g1176 ( 
.A(n_1074),
.B(n_752),
.Y(n_1176)
);

NAND2xp33_ASAP7_75t_SL g1177 ( 
.A(n_1110),
.B(n_761),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1143),
.B(n_904),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1084),
.B(n_762),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1078),
.B(n_909),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1103),
.B(n_913),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1126),
.B(n_766),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1144),
.B(n_772),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1146),
.B(n_1147),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1118),
.B(n_775),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1154),
.B(n_780),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1155),
.B(n_781),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1160),
.B(n_785),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1077),
.B(n_1081),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1094),
.B(n_786),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1099),
.B(n_789),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1139),
.B(n_791),
.Y(n_1192)
);

NAND2xp33_ASAP7_75t_SL g1193 ( 
.A(n_1106),
.B(n_800),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1121),
.B(n_916),
.Y(n_1194)
);

NAND2xp33_ASAP7_75t_SL g1195 ( 
.A(n_1137),
.B(n_1088),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1151),
.B(n_804),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1107),
.B(n_924),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1124),
.B(n_805),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1133),
.B(n_807),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1136),
.B(n_809),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1138),
.B(n_819),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1149),
.B(n_823),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1152),
.B(n_825),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1156),
.B(n_930),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1159),
.B(n_833),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1164),
.B(n_840),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1166),
.B(n_843),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1167),
.B(n_846),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_1169),
.B(n_848),
.Y(n_1209)
);

NAND2xp33_ASAP7_75t_SL g1210 ( 
.A(n_1114),
.B(n_851),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1089),
.B(n_853),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1080),
.B(n_854),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1117),
.B(n_935),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1125),
.B(n_858),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_SL g1215 ( 
.A(n_1153),
.B(n_861),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1100),
.B(n_936),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1129),
.B(n_865),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1090),
.B(n_945),
.Y(n_1218)
);

NAND2xp33_ASAP7_75t_SL g1219 ( 
.A(n_1157),
.B(n_1112),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1115),
.B(n_704),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_1165),
.B(n_871),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1122),
.B(n_959),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_SL g1223 ( 
.A(n_1113),
.B(n_881),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1130),
.B(n_832),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1170),
.B(n_885),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1102),
.B(n_886),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1161),
.B(n_887),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1162),
.B(n_890),
.Y(n_1228)
);

XNOR2xp5_ASAP7_75t_L g1229 ( 
.A(n_1132),
.B(n_891),
.Y(n_1229)
);

NAND2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1142),
.B(n_896),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1120),
.B(n_905),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1092),
.B(n_906),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1116),
.B(n_884),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1096),
.B(n_910),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1101),
.B(n_914),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1082),
.B(n_915),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1108),
.B(n_928),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1141),
.B(n_929),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1091),
.B(n_1145),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1168),
.B(n_933),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1076),
.B(n_934),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1079),
.B(n_939),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1076),
.B(n_941),
.Y(n_1243)
);

NAND2xp33_ASAP7_75t_SL g1244 ( 
.A(n_1140),
.B(n_948),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1095),
.B(n_1123),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1076),
.B(n_949),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1134),
.B(n_950),
.Y(n_1247)
);

NAND2xp33_ASAP7_75t_SL g1248 ( 
.A(n_1148),
.B(n_955),
.Y(n_1248)
);

NAND2xp33_ASAP7_75t_SL g1249 ( 
.A(n_1158),
.B(n_956),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1104),
.B(n_958),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1163),
.B(n_371),
.Y(n_1251)
);

XNOR2x2_ASAP7_75t_L g1252 ( 
.A(n_1128),
.B(n_0),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1131),
.B(n_961),
.Y(n_1253)
);

NAND2xp33_ASAP7_75t_SL g1254 ( 
.A(n_1075),
.B(n_970),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1097),
.B(n_971),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1098),
.B(n_764),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1109),
.B(n_773),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1085),
.B(n_917),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1073),
.B(n_764),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1087),
.B(n_834),
.Y(n_1260)
);

NAND2xp33_ASAP7_75t_SL g1261 ( 
.A(n_1093),
.B(n_707),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1111),
.B(n_834),
.Y(n_1262)
);

NAND2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1093),
.B(n_710),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_SL g1264 ( 
.A(n_1086),
.B(n_712),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1135),
.B(n_842),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1143),
.B(n_964),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1135),
.B(n_864),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1074),
.B(n_717),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1135),
.B(n_864),
.Y(n_1269)
);

NAND2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1150),
.B(n_733),
.Y(n_1270)
);

AND2x2_ASAP7_75t_SL g1271 ( 
.A(n_1135),
.B(n_919),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1074),
.B(n_750),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_SL g1273 ( 
.A(n_1135),
.B(n_864),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1135),
.B(n_864),
.Y(n_1274)
);

NAND2xp33_ASAP7_75t_SL g1275 ( 
.A(n_1150),
.B(n_755),
.Y(n_1275)
);

NAND2xp33_ASAP7_75t_SL g1276 ( 
.A(n_1150),
.B(n_756),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1135),
.B(n_872),
.Y(n_1277)
);

NAND2xp33_ASAP7_75t_SL g1278 ( 
.A(n_1150),
.B(n_757),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1135),
.B(n_872),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1135),
.B(n_872),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1135),
.B(n_872),
.Y(n_1281)
);

NAND2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1150),
.B(n_759),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1135),
.B(n_872),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_SL g1284 ( 
.A(n_1135),
.B(n_919),
.Y(n_1284)
);

NAND2xp33_ASAP7_75t_SL g1285 ( 
.A(n_1150),
.B(n_760),
.Y(n_1285)
);

NAND2xp33_ASAP7_75t_SL g1286 ( 
.A(n_1150),
.B(n_767),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_1135),
.B(n_919),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1135),
.B(n_964),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1135),
.B(n_964),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1074),
.B(n_770),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1135),
.B(n_964),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1135),
.B(n_776),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1143),
.B(n_779),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1135),
.B(n_782),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1143),
.B(n_797),
.Y(n_1295)
);

NAND2xp33_ASAP7_75t_SL g1296 ( 
.A(n_1150),
.B(n_813),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_SL g1297 ( 
.A(n_1150),
.B(n_816),
.Y(n_1297)
);

NAND2xp33_ASAP7_75t_SL g1298 ( 
.A(n_1150),
.B(n_817),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1135),
.B(n_822),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1143),
.B(n_836),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1135),
.B(n_852),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1143),
.B(n_857),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1143),
.B(n_870),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1135),
.B(n_876),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1135),
.B(n_880),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1135),
.B(n_888),
.Y(n_1306)
);

AND2x2_ASAP7_75t_SL g1307 ( 
.A(n_1135),
.B(n_0),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1135),
.B(n_894),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_SL g1309 ( 
.A(n_1135),
.B(n_895),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1143),
.B(n_897),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1135),
.B(n_898),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1074),
.B(n_902),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_SL g1313 ( 
.A(n_1135),
.B(n_907),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1135),
.B(n_908),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1143),
.B(n_911),
.Y(n_1315)
);

NAND2xp33_ASAP7_75t_SL g1316 ( 
.A(n_1150),
.B(n_921),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1135),
.B(n_922),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1135),
.B(n_931),
.Y(n_1318)
);

NAND2xp33_ASAP7_75t_SL g1319 ( 
.A(n_1150),
.B(n_937),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1184),
.A2(n_944),
.B(n_938),
.Y(n_1320)
);

OAI22x1_ASAP7_75t_L g1321 ( 
.A1(n_1229),
.A2(n_952),
.B1(n_953),
.B2(n_951),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1189),
.A2(n_375),
.B(n_374),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1245),
.B(n_1),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1271),
.B(n_957),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1172),
.Y(n_1325)
);

NOR2x1_ASAP7_75t_SL g1326 ( 
.A(n_1231),
.B(n_376),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1315),
.B(n_963),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1293),
.B(n_965),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1295),
.B(n_967),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1178),
.A2(n_379),
.B(n_377),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1307),
.A2(n_968),
.B1(n_4),
.B2(n_2),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1300),
.B(n_2),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1302),
.B(n_3),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1268),
.B(n_3),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1303),
.B(n_4),
.Y(n_1335)
);

O2A1O1Ixp5_ASAP7_75t_L g1336 ( 
.A1(n_1266),
.A2(n_686),
.B(n_688),
.C(n_685),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1233),
.A2(n_382),
.B(n_381),
.Y(n_1337)
);

INVx4_ASAP7_75t_L g1338 ( 
.A(n_1197),
.Y(n_1338)
);

AO32x2_ASAP7_75t_L g1339 ( 
.A1(n_1252),
.A2(n_7),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1218),
.Y(n_1340)
);

NAND3x1_ASAP7_75t_L g1341 ( 
.A(n_1258),
.B(n_5),
.C(n_6),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1179),
.A2(n_385),
.B(n_383),
.Y(n_1342)
);

AO21x1_ASAP7_75t_L g1343 ( 
.A1(n_1310),
.A2(n_8),
.B(n_9),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1222),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1194),
.Y(n_1345)
);

OAI22x1_ASAP7_75t_L g1346 ( 
.A1(n_1251),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1204),
.Y(n_1347)
);

NAND3xp33_ASAP7_75t_L g1348 ( 
.A(n_1210),
.B(n_12),
.C(n_13),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1213),
.A2(n_387),
.B(n_386),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1198),
.A2(n_390),
.B(n_389),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1180),
.B(n_12),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1272),
.B(n_14),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1224),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1199),
.A2(n_392),
.B(n_391),
.Y(n_1354)
);

AO21x2_ASAP7_75t_L g1355 ( 
.A1(n_1182),
.A2(n_395),
.B(n_394),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1227),
.A2(n_397),
.B(n_396),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1292),
.B(n_14),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1175),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1228),
.A2(n_400),
.B(n_398),
.Y(n_1359)
);

AO21x1_ASAP7_75t_L g1360 ( 
.A1(n_1254),
.A2(n_1248),
.B(n_1244),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1220),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1251),
.A2(n_1265),
.B(n_1239),
.Y(n_1362)
);

A2O1A1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1288),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1200),
.A2(n_404),
.B(n_403),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1201),
.A2(n_1203),
.B(n_1202),
.Y(n_1365)
);

AO31x2_ASAP7_75t_L g1366 ( 
.A1(n_1257),
.A2(n_691),
.A3(n_692),
.B(n_690),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1290),
.B(n_1312),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1181),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1216),
.B(n_15),
.Y(n_1369)
);

AO31x2_ASAP7_75t_L g1370 ( 
.A1(n_1241),
.A2(n_406),
.A3(n_409),
.B(n_405),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1205),
.A2(n_411),
.B(n_410),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1216),
.B(n_16),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1174),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1175),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1289),
.B(n_17),
.Y(n_1375)
);

AO21x1_ASAP7_75t_L g1376 ( 
.A1(n_1249),
.A2(n_18),
.B(n_19),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1206),
.A2(n_414),
.B(n_412),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1207),
.A2(n_418),
.B(n_416),
.Y(n_1378)
);

NAND2x1_ASAP7_75t_L g1379 ( 
.A(n_1197),
.B(n_419),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_L g1380 ( 
.A(n_1243),
.B(n_422),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1208),
.A2(n_1209),
.B(n_1211),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1291),
.B(n_20),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1246),
.A2(n_425),
.B(n_423),
.Y(n_1383)
);

AO31x2_ASAP7_75t_L g1384 ( 
.A1(n_1235),
.A2(n_678),
.A3(n_679),
.B(n_676),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1171),
.A2(n_431),
.B1(n_432),
.B2(n_430),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1237),
.A2(n_435),
.B(n_433),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1195),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1267),
.A2(n_441),
.B(n_437),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1219),
.B(n_442),
.Y(n_1389)
);

NOR2xp67_ASAP7_75t_L g1390 ( 
.A(n_1242),
.B(n_444),
.Y(n_1390)
);

OR2x6_ASAP7_75t_L g1391 ( 
.A(n_1256),
.B(n_21),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1215),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1269),
.A2(n_448),
.B(n_445),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1183),
.B(n_21),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1190),
.A2(n_450),
.B(n_449),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1191),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1186),
.A2(n_453),
.B(n_451),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1273),
.A2(n_455),
.B(n_454),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1226),
.B(n_456),
.Y(n_1399)
);

O2A1O1Ixp5_ASAP7_75t_L g1400 ( 
.A1(n_1274),
.A2(n_682),
.B(n_683),
.C(n_681),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1294),
.B(n_22),
.C(n_23),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1277),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1187),
.B(n_22),
.Y(n_1403)
);

AO22x2_ASAP7_75t_L g1404 ( 
.A1(n_1260),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1193),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1279),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1280),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1232),
.A2(n_1234),
.B(n_1236),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1188),
.B(n_27),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1281),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1255),
.Y(n_1411)
);

AOI211x1_ASAP7_75t_L g1412 ( 
.A1(n_1283),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1412)
);

AOI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1238),
.A2(n_1221),
.B(n_1217),
.Y(n_1413)
);

AO31x2_ASAP7_75t_L g1414 ( 
.A1(n_1177),
.A2(n_674),
.A3(n_675),
.B(n_673),
.Y(n_1414)
);

NOR3xp33_ASAP7_75t_SL g1415 ( 
.A(n_1261),
.B(n_29),
.C(n_30),
.Y(n_1415)
);

OR2x6_ASAP7_75t_L g1416 ( 
.A(n_1247),
.B(n_1284),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1196),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1287),
.A2(n_34),
.B(n_31),
.C(n_33),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1240),
.A2(n_459),
.B(n_457),
.Y(n_1419)
);

XOR2xp5_ASAP7_75t_L g1420 ( 
.A(n_1212),
.B(n_460),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1225),
.A2(n_462),
.B(n_461),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1319),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1299),
.B(n_31),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1253),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1301),
.B(n_463),
.Y(n_1425)
);

BUFx12f_ASAP7_75t_L g1426 ( 
.A(n_1270),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1176),
.A2(n_465),
.B(n_464),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1304),
.B(n_33),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1262),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1214),
.A2(n_1306),
.B(n_1305),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1308),
.B(n_34),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1318),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1432)
);

INVxp67_ASAP7_75t_SL g1433 ( 
.A(n_1368),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1360),
.A2(n_1263),
.A3(n_1311),
.B(n_1309),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1327),
.B(n_1314),
.Y(n_1435)
);

INVxp33_ASAP7_75t_L g1436 ( 
.A(n_1367),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1337),
.A2(n_1250),
.B(n_1192),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1361),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1345),
.A2(n_1230),
.B(n_1313),
.Y(n_1439)
);

AOI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1357),
.A2(n_1264),
.B1(n_1259),
.B2(n_1317),
.C(n_1276),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1334),
.B(n_1173),
.Y(n_1441)
);

OAI22x1_ASAP7_75t_L g1442 ( 
.A1(n_1428),
.A2(n_1275),
.B1(n_1278),
.B2(n_1282),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1358),
.B(n_36),
.Y(n_1443)
);

INVx4_ASAP7_75t_L g1444 ( 
.A(n_1338),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1413),
.A2(n_1223),
.B(n_1185),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1393),
.A2(n_467),
.B(n_466),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1347),
.Y(n_1447)
);

INVx6_ASAP7_75t_L g1448 ( 
.A(n_1426),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1411),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1407),
.A2(n_1286),
.B1(n_1296),
.B2(n_1285),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1398),
.A2(n_469),
.B(n_468),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1371),
.A2(n_473),
.B(n_472),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1374),
.Y(n_1453)
);

CKINVDCx16_ASAP7_75t_R g1454 ( 
.A(n_1325),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1335),
.A2(n_1298),
.B(n_1297),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1373),
.B(n_38),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1377),
.A2(n_476),
.B(n_474),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1320),
.B(n_39),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1378),
.A2(n_478),
.B(n_477),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1381),
.A2(n_1316),
.B(n_482),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1328),
.B(n_39),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1387),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1340),
.B(n_40),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_SL g1464 ( 
.A1(n_1326),
.A2(n_1376),
.B(n_1343),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1332),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1344),
.Y(n_1466)
);

AO21x2_ASAP7_75t_L g1467 ( 
.A1(n_1389),
.A2(n_483),
.B(n_479),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1353),
.Y(n_1468)
);

BUFx2_ASAP7_75t_L g1469 ( 
.A(n_1417),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1369),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1329),
.B(n_41),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1423),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_L g1473 ( 
.A1(n_1321),
.A2(n_1401),
.B1(n_1331),
.B2(n_1432),
.C(n_1346),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1356),
.A2(n_486),
.B(n_485),
.Y(n_1474)
);

CKINVDCx12_ASAP7_75t_R g1475 ( 
.A(n_1416),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1372),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1402),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1333),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1359),
.A2(n_489),
.B(n_488),
.Y(n_1479)
);

NAND2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1379),
.B(n_497),
.Y(n_1480)
);

BUFx4_ASAP7_75t_SL g1481 ( 
.A(n_1323),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1362),
.A2(n_494),
.B(n_490),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_SL g1483 ( 
.A1(n_1363),
.A2(n_498),
.B(n_502),
.C(n_495),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1386),
.A2(n_506),
.B(n_504),
.Y(n_1484)
);

BUFx4f_ASAP7_75t_L g1485 ( 
.A(n_1416),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1349),
.A2(n_509),
.B(n_507),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1410),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1323),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1352),
.B(n_44),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1399),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1396),
.Y(n_1491)
);

AO31x2_ASAP7_75t_L g1492 ( 
.A1(n_1405),
.A2(n_512),
.A3(n_513),
.B(n_511),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_L g1493 ( 
.A(n_1415),
.B(n_1348),
.C(n_1431),
.Y(n_1493)
);

AOI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1408),
.A2(n_515),
.B(n_514),
.Y(n_1494)
);

AOI21xp33_ASAP7_75t_L g1495 ( 
.A1(n_1424),
.A2(n_45),
.B(n_46),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1391),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1383),
.A2(n_517),
.B(n_516),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1392),
.B(n_45),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1420),
.A2(n_1391),
.B1(n_1324),
.B2(n_1394),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1404),
.B(n_46),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1429),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1351),
.B(n_47),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1422),
.B(n_47),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1430),
.B(n_518),
.Y(n_1504)
);

A2O1A1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1365),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_1505)
);

OAI22x1_ASAP7_75t_L g1506 ( 
.A1(n_1425),
.A2(n_51),
.B1(n_53),
.B2(n_50),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1403),
.Y(n_1507)
);

A2O1A1Ixp33_ASAP7_75t_L g1508 ( 
.A1(n_1409),
.A2(n_53),
.B(n_48),
.C(n_51),
.Y(n_1508)
);

BUFx2_ASAP7_75t_SL g1509 ( 
.A(n_1390),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_R g1510 ( 
.A1(n_1385),
.A2(n_54),
.B(n_55),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1380),
.A2(n_520),
.B(n_519),
.Y(n_1511)
);

INVx4_ASAP7_75t_SL g1512 ( 
.A(n_1414),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1375),
.B(n_54),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1382),
.A2(n_1406),
.B1(n_1404),
.B2(n_1388),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1355),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1419),
.A2(n_523),
.B(n_521),
.Y(n_1516)
);

O2A1O1Ixp33_ASAP7_75t_L g1517 ( 
.A1(n_1418),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1427),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1400),
.A2(n_526),
.B(n_525),
.Y(n_1519)
);

INVx5_ASAP7_75t_L g1520 ( 
.A(n_1341),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1339),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1421),
.A2(n_1342),
.B1(n_1395),
.B2(n_1330),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1397),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1523)
);

AOI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1322),
.A2(n_1354),
.B(n_1350),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_SL g1525 ( 
.A1(n_1364),
.A2(n_528),
.B(n_527),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1339),
.A2(n_1412),
.B1(n_62),
.B2(n_59),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1366),
.Y(n_1527)
);

BUFx4f_ASAP7_75t_L g1528 ( 
.A(n_1414),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1384),
.A2(n_532),
.B(n_529),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1366),
.B(n_61),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1384),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1370),
.A2(n_65),
.B1(n_62),
.B2(n_63),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1345),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1336),
.A2(n_534),
.B(n_533),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1327),
.B(n_66),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1327),
.A2(n_537),
.B(n_535),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1327),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1358),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1361),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1327),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1334),
.B(n_69),
.Y(n_1541)
);

INVx6_ASAP7_75t_L g1542 ( 
.A(n_1426),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1337),
.A2(n_540),
.B(n_538),
.Y(n_1543)
);

OA21x2_ASAP7_75t_L g1544 ( 
.A1(n_1336),
.A2(n_542),
.B(n_541),
.Y(n_1544)
);

CKINVDCx20_ASAP7_75t_R g1545 ( 
.A(n_1325),
.Y(n_1545)
);

AOI21xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1331),
.A2(n_70),
.B(n_71),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1327),
.A2(n_73),
.B(n_70),
.C(n_72),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1337),
.A2(n_548),
.B(n_547),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1368),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1360),
.A2(n_550),
.B(n_549),
.Y(n_1550)
);

AOI222xp33_ASAP7_75t_L g1551 ( 
.A1(n_1331),
.A2(n_74),
.B1(n_76),
.B2(n_72),
.C1(n_73),
.C2(n_75),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1361),
.Y(n_1552)
);

OAI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1327),
.A2(n_78),
.B1(n_75),
.B2(n_77),
.Y(n_1553)
);

NAND2x1p5_ASAP7_75t_L g1554 ( 
.A(n_1338),
.B(n_555),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_L g1555 ( 
.A(n_1361),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1462),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1435),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.C(n_81),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1527),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1531),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1468),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1447),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1436),
.B(n_79),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1535),
.B(n_551),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1555),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1555),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1533),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1466),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1489),
.B(n_82),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1539),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1477),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1487),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1543),
.A2(n_1548),
.B(n_1486),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1501),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1448),
.B(n_554),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1538),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1514),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1454),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1453),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1493),
.A2(n_85),
.B(n_86),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1469),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1476),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1463),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1470),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1491),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1507),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1541),
.B(n_86),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1549),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1502),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1472),
.B(n_1449),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1521),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1441),
.B(n_87),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1497),
.A2(n_557),
.B(n_556),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1438),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1521),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1448),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1542),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1461),
.B(n_87),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1542),
.B(n_558),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1552),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1443),
.B(n_88),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1485),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1494),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1471),
.Y(n_1603)
);

CKINVDCx16_ASAP7_75t_R g1604 ( 
.A(n_1545),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1481),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1504),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1512),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1490),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1433),
.B(n_89),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1464),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1512),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1446),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1451),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1474),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1456),
.B(n_89),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1524),
.A2(n_1479),
.B(n_1457),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1490),
.B(n_1444),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1458),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1513),
.B(n_90),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1473),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1530),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1506),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1551),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1526),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1440),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1452),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1509),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1459),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1528),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1496),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1582),
.B(n_1500),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1580),
.B(n_1520),
.Y(n_1632)
);

INVx3_ASAP7_75t_L g1633 ( 
.A(n_1564),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1556),
.Y(n_1634)
);

NAND2xp33_ASAP7_75t_R g1635 ( 
.A(n_1577),
.B(n_1488),
.Y(n_1635)
);

NAND2xp33_ASAP7_75t_R g1636 ( 
.A(n_1605),
.B(n_1503),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_R g1637 ( 
.A(n_1604),
.B(n_1475),
.Y(n_1637)
);

CKINVDCx11_ASAP7_75t_R g1638 ( 
.A(n_1595),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1591),
.B(n_1520),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1585),
.B(n_1498),
.Y(n_1640)
);

XNOR2xp5_ASAP7_75t_L g1641 ( 
.A(n_1601),
.B(n_1596),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1588),
.B(n_1499),
.Y(n_1642)
);

NAND2xp33_ASAP7_75t_R g1643 ( 
.A(n_1574),
.B(n_1546),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1565),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1581),
.B(n_1603),
.Y(n_1645)
);

BUFx10_ASAP7_75t_L g1646 ( 
.A(n_1617),
.Y(n_1646)
);

NAND2xp33_ASAP7_75t_R g1647 ( 
.A(n_1574),
.B(n_1536),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_R g1648 ( 
.A(n_1608),
.B(n_1515),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1618),
.B(n_1583),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1606),
.B(n_1434),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_R g1651 ( 
.A(n_1569),
.B(n_1511),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1630),
.B(n_1455),
.Y(n_1652)
);

NAND2xp33_ASAP7_75t_SL g1653 ( 
.A(n_1623),
.B(n_1442),
.Y(n_1653)
);

NAND2xp33_ASAP7_75t_R g1654 ( 
.A(n_1598),
.B(n_1534),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1558),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_R g1656 ( 
.A(n_1629),
.B(n_1478),
.Y(n_1656)
);

NAND2xp33_ASAP7_75t_R g1657 ( 
.A(n_1598),
.B(n_1544),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1593),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1587),
.B(n_1561),
.Y(n_1659)
);

OR2x6_ASAP7_75t_L g1660 ( 
.A(n_1629),
.B(n_1554),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1566),
.B(n_1465),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1560),
.B(n_1495),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1589),
.B(n_1450),
.Y(n_1663)
);

NAND2xp33_ASAP7_75t_R g1664 ( 
.A(n_1617),
.B(n_1439),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1564),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1573),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1584),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1599),
.B(n_1508),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_R g1669 ( 
.A(n_1627),
.B(n_1537),
.Y(n_1669)
);

INVx2_ASAP7_75t_SL g1670 ( 
.A(n_1578),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1570),
.B(n_1492),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1567),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_R g1673 ( 
.A(n_1621),
.B(n_1510),
.Y(n_1673)
);

OR2x4_ASAP7_75t_L g1674 ( 
.A(n_1622),
.B(n_1553),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1634),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1655),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1663),
.B(n_1562),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1667),
.B(n_1590),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1653),
.A2(n_1579),
.B1(n_1557),
.B2(n_1576),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1670),
.B(n_1594),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1659),
.B(n_1631),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1649),
.B(n_1559),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1672),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1658),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1645),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1642),
.B(n_1559),
.Y(n_1686)
);

NOR2x1_ASAP7_75t_SL g1687 ( 
.A(n_1660),
.B(n_1607),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1666),
.Y(n_1688)
);

NOR2x1p5_ASAP7_75t_L g1689 ( 
.A(n_1662),
.B(n_1619),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1671),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1652),
.B(n_1571),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1638),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1639),
.B(n_1568),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1650),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1668),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1648),
.B(n_1615),
.Y(n_1696)
);

OR2x6_ASAP7_75t_SL g1697 ( 
.A(n_1661),
.B(n_1597),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1632),
.B(n_1586),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1640),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1633),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1674),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1646),
.B(n_1600),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1673),
.B(n_1563),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1656),
.A2(n_1624),
.B1(n_1625),
.B2(n_1620),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1637),
.B(n_1610),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1665),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1669),
.B(n_1575),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1644),
.B(n_1560),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1641),
.B(n_1609),
.Y(n_1709)
);

INVxp67_ASAP7_75t_SL g1710 ( 
.A(n_1664),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1651),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1660),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1636),
.B(n_1607),
.Y(n_1713)
);

BUFx2_ASAP7_75t_SL g1714 ( 
.A(n_1635),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1654),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1647),
.B(n_1611),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1657),
.B(n_1611),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1643),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1676),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_SL g1720 ( 
.A(n_1715),
.B(n_1460),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1691),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1716),
.B(n_1677),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1679),
.A2(n_1540),
.B1(n_1547),
.B2(n_1523),
.C(n_1505),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1683),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1705),
.B(n_1492),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1681),
.B(n_1602),
.Y(n_1726)
);

OR2x6_ASAP7_75t_L g1727 ( 
.A(n_1714),
.B(n_1482),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1692),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1717),
.B(n_1675),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1717),
.B(n_1529),
.Y(n_1730)
);

AOI221xp5_ASAP7_75t_L g1731 ( 
.A1(n_1704),
.A2(n_1518),
.B1(n_1532),
.B2(n_1517),
.C(n_1483),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1682),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1685),
.B(n_1445),
.Y(n_1733)
);

INVxp67_ASAP7_75t_SL g1734 ( 
.A(n_1686),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1688),
.Y(n_1735)
);

OAI33xp33_ASAP7_75t_L g1736 ( 
.A1(n_1701),
.A2(n_1703),
.A3(n_1718),
.B1(n_1711),
.B2(n_1712),
.B3(n_1699),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1708),
.B(n_1710),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1707),
.B(n_1522),
.C(n_1519),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1696),
.B(n_1550),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1680),
.Y(n_1740)
);

NOR3xp33_ASAP7_75t_SL g1741 ( 
.A(n_1694),
.B(n_1525),
.C(n_95),
.Y(n_1741)
);

OAI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1684),
.A2(n_1480),
.B1(n_1613),
.B2(n_1614),
.C(n_1612),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1690),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_1697),
.B(n_96),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1678),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_L g1746 ( 
.A(n_1695),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1706),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1689),
.A2(n_1467),
.B1(n_1437),
.B2(n_1626),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1700),
.B(n_1628),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1702),
.B(n_97),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1693),
.B(n_1616),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1698),
.B(n_1592),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1687),
.A2(n_1572),
.B1(n_1516),
.B2(n_1484),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1709),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1714),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1676),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1713),
.B(n_100),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1676),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1717),
.B(n_101),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1683),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1717),
.B(n_102),
.Y(n_1761)
);

BUFx2_ASAP7_75t_SL g1762 ( 
.A(n_1717),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1713),
.B(n_103),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1713),
.B(n_103),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1683),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1683),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_R g1767 ( 
.A(n_1692),
.B(n_104),
.Y(n_1767)
);

OAI31xp33_ASAP7_75t_L g1768 ( 
.A1(n_1679),
.A2(n_106),
.A3(n_104),
.B(n_105),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1683),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1715),
.B(n_108),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1679),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1676),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1713),
.B(n_109),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1713),
.B(n_110),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1722),
.B(n_111),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1734),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1762),
.B(n_113),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1721),
.B(n_114),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1745),
.B(n_115),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1737),
.B(n_115),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1724),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1740),
.B(n_1760),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1755),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1746),
.Y(n_1784)
);

OR2x6_ASAP7_75t_L g1785 ( 
.A(n_1727),
.B(n_117),
.Y(n_1785)
);

NAND2x1_ASAP7_75t_L g1786 ( 
.A(n_1751),
.B(n_117),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1719),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1754),
.B(n_1743),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1735),
.B(n_118),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1765),
.B(n_118),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1766),
.B(n_119),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1769),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1747),
.B(n_120),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1730),
.B(n_120),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1725),
.B(n_121),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1756),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1726),
.B(n_123),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1728),
.B(n_124),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1767),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1733),
.B(n_125),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1758),
.B(n_126),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1772),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1749),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1744),
.B(n_1750),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1739),
.B(n_126),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1752),
.B(n_127),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1757),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1768),
.B(n_128),
.C(n_129),
.Y(n_1808)
);

AND2x4_ASAP7_75t_SL g1809 ( 
.A(n_1759),
.B(n_559),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1759),
.B(n_129),
.Y(n_1810)
);

NAND2x1p5_ASAP7_75t_L g1811 ( 
.A(n_1761),
.B(n_560),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1761),
.B(n_130),
.Y(n_1812)
);

NOR2x1p5_ASAP7_75t_L g1813 ( 
.A(n_1770),
.B(n_131),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1738),
.B(n_132),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1727),
.B(n_132),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1763),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1764),
.B(n_1773),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1720),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1742),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1774),
.B(n_133),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1731),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1736),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1748),
.B(n_135),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1741),
.B(n_136),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1753),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1723),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1771),
.B(n_136),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1724),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1719),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1721),
.B(n_137),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1721),
.B(n_138),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1719),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1732),
.B(n_139),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1729),
.B(n_139),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1729),
.B(n_140),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1729),
.B(n_140),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1719),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1729),
.B(n_141),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1719),
.Y(n_1839)
);

INVxp67_ASAP7_75t_SL g1840 ( 
.A(n_1732),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_SL g1841 ( 
.A(n_1762),
.B(n_142),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1782),
.Y(n_1842)
);

INVx4_ASAP7_75t_L g1843 ( 
.A(n_1836),
.Y(n_1843)
);

INVx2_ASAP7_75t_SL g1844 ( 
.A(n_1784),
.Y(n_1844)
);

NOR4xp25_ASAP7_75t_SL g1845 ( 
.A(n_1776),
.B(n_1825),
.C(n_1840),
.D(n_1814),
.Y(n_1845)
);

OAI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1821),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1819),
.B(n_144),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1822),
.B(n_146),
.Y(n_1848)
);

INVx3_ASAP7_75t_L g1849 ( 
.A(n_1783),
.Y(n_1849)
);

INVxp33_ASAP7_75t_SL g1850 ( 
.A(n_1799),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1788),
.B(n_147),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1803),
.B(n_150),
.Y(n_1852)
);

AO221x2_ASAP7_75t_L g1853 ( 
.A1(n_1817),
.A2(n_153),
.B1(n_155),
.B2(n_152),
.C(n_154),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1800),
.B(n_151),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1787),
.Y(n_1855)
);

NAND2xp33_ASAP7_75t_SL g1856 ( 
.A(n_1813),
.B(n_153),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1815),
.Y(n_1857)
);

NOR2x1_ASAP7_75t_L g1858 ( 
.A(n_1777),
.B(n_156),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_SL g1859 ( 
.A(n_1826),
.B(n_157),
.Y(n_1859)
);

OAI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1785),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.Y(n_1860)
);

AO221x2_ASAP7_75t_L g1861 ( 
.A1(n_1808),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.C(n_163),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1805),
.B(n_162),
.Y(n_1862)
);

NOR2x1_ASAP7_75t_L g1863 ( 
.A(n_1818),
.B(n_164),
.Y(n_1863)
);

AO221x2_ASAP7_75t_L g1864 ( 
.A1(n_1780),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_167),
.Y(n_1864)
);

NOR2x1_ASAP7_75t_L g1865 ( 
.A(n_1778),
.B(n_165),
.Y(n_1865)
);

INVxp33_ASAP7_75t_SL g1866 ( 
.A(n_1807),
.Y(n_1866)
);

OAI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1785),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_1867)
);

OAI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1804),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.C(n_171),
.Y(n_1868)
);

AO221x2_ASAP7_75t_L g1869 ( 
.A1(n_1830),
.A2(n_172),
.B1(n_174),
.B2(n_170),
.C(n_173),
.Y(n_1869)
);

OAI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1786),
.A2(n_1806),
.B1(n_1816),
.B2(n_1831),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1781),
.B(n_172),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1796),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1792),
.B(n_1828),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1802),
.Y(n_1874)
);

AO221x2_ASAP7_75t_L g1875 ( 
.A1(n_1789),
.A2(n_1793),
.B1(n_1797),
.B2(n_1832),
.C(n_1829),
.Y(n_1875)
);

OAI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1824),
.A2(n_1811),
.B1(n_1791),
.B2(n_1790),
.C(n_1827),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1836),
.B(n_176),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1833),
.A2(n_1823),
.B1(n_1794),
.B2(n_1837),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1839),
.B(n_176),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1794),
.B(n_177),
.Y(n_1880)
);

NOR2x1_ASAP7_75t_L g1881 ( 
.A(n_1801),
.B(n_179),
.Y(n_1881)
);

NOR2x1_ASAP7_75t_L g1882 ( 
.A(n_1801),
.B(n_179),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1820),
.B(n_180),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1795),
.B(n_180),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_R g1885 ( 
.A(n_1810),
.B(n_182),
.Y(n_1885)
);

OAI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1775),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_SL g1887 ( 
.A(n_1812),
.B(n_183),
.Y(n_1887)
);

AO221x2_ASAP7_75t_L g1888 ( 
.A1(n_1841),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.C(n_188),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1834),
.B(n_189),
.Y(n_1889)
);

AO221x2_ASAP7_75t_L g1890 ( 
.A1(n_1835),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.C(n_193),
.Y(n_1890)
);

NAND2xp33_ASAP7_75t_SL g1891 ( 
.A(n_1838),
.B(n_191),
.Y(n_1891)
);

AOI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1809),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_1892)
);

OAI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1779),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.C(n_198),
.Y(n_1893)
);

NOR2xp67_ASAP7_75t_L g1894 ( 
.A(n_1798),
.B(n_195),
.Y(n_1894)
);

OAI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1821),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_1895)
);

INVxp67_ASAP7_75t_L g1896 ( 
.A(n_1819),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1783),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1784),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1826),
.B(n_199),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1819),
.B(n_200),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1808),
.A2(n_206),
.B1(n_203),
.B2(n_205),
.Y(n_1901)
);

OAI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1821),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.C(n_208),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1819),
.B(n_207),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1787),
.Y(n_1904)
);

AO221x2_ASAP7_75t_L g1905 ( 
.A1(n_1822),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.C(n_211),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1821),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1819),
.B(n_215),
.Y(n_1907)
);

INVxp33_ASAP7_75t_SL g1908 ( 
.A(n_1799),
.Y(n_1908)
);

NOR2x1_ASAP7_75t_L g1909 ( 
.A(n_1822),
.B(n_215),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_SL g1910 ( 
.A(n_1783),
.B(n_217),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1819),
.B(n_218),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1783),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1822),
.B(n_218),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1819),
.B(n_220),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_R g1915 ( 
.A(n_1799),
.B(n_222),
.Y(n_1915)
);

AO221x2_ASAP7_75t_L g1916 ( 
.A1(n_1822),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.C(n_226),
.Y(n_1916)
);

AOI221x1_ASAP7_75t_SL g1917 ( 
.A1(n_1826),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.C(n_226),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1819),
.B(n_227),
.Y(n_1918)
);

OAI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1821),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1819),
.B(n_229),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1857),
.B(n_230),
.Y(n_1921)
);

NAND2x1_ASAP7_75t_L g1922 ( 
.A(n_1849),
.B(n_1844),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1897),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1842),
.B(n_232),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_1912),
.Y(n_1925)
);

INVx1_ASAP7_75t_SL g1926 ( 
.A(n_1915),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1898),
.B(n_233),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1872),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1874),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1904),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1875),
.B(n_233),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_R g1932 ( 
.A(n_1856),
.B(n_234),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1873),
.Y(n_1933)
);

INVx1_ASAP7_75t_SL g1934 ( 
.A(n_1850),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1861),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1909),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1843),
.B(n_236),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1913),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1908),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1861),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1851),
.B(n_238),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1871),
.Y(n_1942)
);

AOI22x1_ASAP7_75t_L g1943 ( 
.A1(n_1880),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1902),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1870),
.B(n_242),
.Y(n_1945)
);

OR2x6_ASAP7_75t_L g1946 ( 
.A(n_1881),
.B(n_244),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1866),
.Y(n_1947)
);

INVxp67_ASAP7_75t_L g1948 ( 
.A(n_1863),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1852),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1879),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1848),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1847),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1858),
.B(n_245),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1900),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1903),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1882),
.B(n_246),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1907),
.Y(n_1957)
);

OR2x2_ASAP7_75t_L g1958 ( 
.A(n_1878),
.B(n_246),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1911),
.B(n_247),
.Y(n_1959)
);

AND2x4_ASAP7_75t_L g1960 ( 
.A(n_1894),
.B(n_248),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1914),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1885),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1865),
.Y(n_1963)
);

INVx3_ASAP7_75t_L g1964 ( 
.A(n_1888),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1920),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1918),
.B(n_248),
.Y(n_1966)
);

NAND2x1_ASAP7_75t_SL g1967 ( 
.A(n_1877),
.B(n_249),
.Y(n_1967)
);

NAND2x1_ASAP7_75t_L g1968 ( 
.A(n_1854),
.B(n_249),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1876),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1862),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_SL g1971 ( 
.A(n_1859),
.B(n_250),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_R g1972 ( 
.A(n_1891),
.B(n_250),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_SL g1973 ( 
.A1(n_1853),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1910),
.Y(n_1974)
);

BUFx2_ASAP7_75t_L g1975 ( 
.A(n_1884),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1883),
.B(n_254),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1905),
.Y(n_1977)
);

AND2x4_ASAP7_75t_SL g1978 ( 
.A(n_1892),
.B(n_255),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1889),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1899),
.B(n_255),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_L g1981 ( 
.A(n_1887),
.B(n_258),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1864),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1864),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1916),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1901),
.B(n_259),
.Y(n_1985)
);

INVxp67_ASAP7_75t_L g1986 ( 
.A(n_1893),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1890),
.B(n_259),
.Y(n_1987)
);

INVx1_ASAP7_75t_SL g1988 ( 
.A(n_1869),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1886),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1868),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1917),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1860),
.B(n_260),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1867),
.B(n_260),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1846),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1919),
.B(n_261),
.Y(n_1995)
);

INVx3_ASAP7_75t_L g1996 ( 
.A(n_1895),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1906),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1896),
.B(n_262),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1855),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1857),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1855),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1845),
.A2(n_264),
.B(n_266),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1857),
.B(n_267),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1861),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1857),
.B(n_269),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1855),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1857),
.B(n_270),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1896),
.B(n_270),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1855),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_1897),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1857),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1896),
.B(n_272),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1857),
.B(n_272),
.Y(n_2013)
);

INVx1_ASAP7_75t_SL g2014 ( 
.A(n_1897),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1896),
.B(n_273),
.Y(n_2015)
);

NOR2x1_ASAP7_75t_L g2016 ( 
.A(n_1863),
.B(n_274),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1857),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1855),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1857),
.B(n_275),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1857),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1896),
.B(n_276),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1896),
.B(n_278),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1896),
.B(n_278),
.Y(n_2023)
);

INVx3_ASAP7_75t_L g2024 ( 
.A(n_1843),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1857),
.B(n_279),
.Y(n_2025)
);

INVx1_ASAP7_75t_SL g2026 ( 
.A(n_1897),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1857),
.B(n_280),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1857),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1857),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1896),
.B(n_281),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_1934),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1963),
.B(n_284),
.Y(n_2032)
);

INVxp33_ASAP7_75t_L g2033 ( 
.A(n_1947),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1930),
.Y(n_2034)
);

INVx1_ASAP7_75t_SL g2035 ( 
.A(n_1939),
.Y(n_2035)
);

OAI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_2002),
.A2(n_286),
.B(n_287),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_2024),
.B(n_2000),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1928),
.Y(n_2038)
);

OAI21xp33_ASAP7_75t_SL g2039 ( 
.A1(n_1931),
.A2(n_288),
.B(n_289),
.Y(n_2039)
);

AOI322xp5_ASAP7_75t_L g2040 ( 
.A1(n_1988),
.A2(n_293),
.A3(n_292),
.B1(n_290),
.B2(n_288),
.C1(n_289),
.C2(n_291),
.Y(n_2040)
);

AOI221xp5_ASAP7_75t_L g2041 ( 
.A1(n_1986),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.C(n_293),
.Y(n_2041)
);

OAI221xp5_ASAP7_75t_SL g2042 ( 
.A1(n_1935),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.C(n_297),
.Y(n_2042)
);

NAND3xp33_ASAP7_75t_L g2043 ( 
.A(n_1936),
.B(n_294),
.C(n_295),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1938),
.B(n_298),
.Y(n_2044)
);

AOI21xp33_ASAP7_75t_SL g2045 ( 
.A1(n_1984),
.A2(n_299),
.B(n_300),
.Y(n_2045)
);

INVx3_ASAP7_75t_L g2046 ( 
.A(n_1922),
.Y(n_2046)
);

AOI221xp5_ASAP7_75t_L g2047 ( 
.A1(n_1996),
.A2(n_1964),
.B1(n_1983),
.B2(n_1991),
.C(n_1990),
.Y(n_2047)
);

OAI21xp33_ASAP7_75t_L g2048 ( 
.A1(n_1973),
.A2(n_301),
.B(n_302),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1945),
.A2(n_1948),
.B(n_2016),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1977),
.B(n_301),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1929),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1982),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1999),
.Y(n_2053)
);

OAI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_1940),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2011),
.B(n_2017),
.Y(n_2055)
);

O2A1O1Ixp33_ASAP7_75t_L g2056 ( 
.A1(n_1946),
.A2(n_309),
.B(n_307),
.C(n_308),
.Y(n_2056)
);

OAI322xp33_ASAP7_75t_L g2057 ( 
.A1(n_1995),
.A2(n_309),
.A3(n_310),
.B1(n_311),
.B2(n_312),
.C1(n_313),
.C2(n_314),
.Y(n_2057)
);

OR2x2_ASAP7_75t_L g2058 ( 
.A(n_2020),
.B(n_310),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1965),
.B(n_311),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2028),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1952),
.B(n_313),
.Y(n_2061)
);

AOI221xp5_ASAP7_75t_L g2062 ( 
.A1(n_1997),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.C(n_317),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1954),
.B(n_1955),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2001),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1971),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1946),
.A2(n_318),
.B(n_319),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_2029),
.B(n_320),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2006),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2009),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1957),
.B(n_321),
.Y(n_2070)
);

O2A1O1Ixp33_ASAP7_75t_L g2071 ( 
.A1(n_1958),
.A2(n_323),
.B(n_321),
.C(n_322),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_1951),
.B(n_322),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1961),
.B(n_323),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1923),
.B(n_324),
.Y(n_2074)
);

OAI21xp5_ASAP7_75t_L g2075 ( 
.A1(n_1981),
.A2(n_325),
.B(n_326),
.Y(n_2075)
);

OAI21xp33_ASAP7_75t_L g2076 ( 
.A1(n_1944),
.A2(n_327),
.B(n_328),
.Y(n_2076)
);

OAI322xp33_ASAP7_75t_L g2077 ( 
.A1(n_1992),
.A2(n_328),
.A3(n_330),
.B1(n_331),
.B2(n_332),
.C1(n_333),
.C2(n_334),
.Y(n_2077)
);

OAI21xp33_ASAP7_75t_L g2078 ( 
.A1(n_2004),
.A2(n_336),
.B(n_337),
.Y(n_2078)
);

OAI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1987),
.A2(n_336),
.B(n_338),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1975),
.B(n_338),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_1969),
.B(n_339),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_1933),
.B(n_339),
.Y(n_2082)
);

AOI22xp5_ASAP7_75t_L g2083 ( 
.A1(n_1994),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_2083)
);

NAND2x1_ASAP7_75t_L g2084 ( 
.A(n_2018),
.B(n_343),
.Y(n_2084)
);

AOI322xp5_ASAP7_75t_L g2085 ( 
.A1(n_1989),
.A2(n_344),
.A3(n_345),
.B1(n_346),
.B2(n_347),
.C1(n_348),
.C2(n_349),
.Y(n_2085)
);

OAI211xp5_ASAP7_75t_L g2086 ( 
.A1(n_1972),
.A2(n_348),
.B(n_344),
.C(n_345),
.Y(n_2086)
);

AOI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_1985),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_2087)
);

AOI211xp5_ASAP7_75t_L g2088 ( 
.A1(n_1932),
.A2(n_1985),
.B(n_1980),
.C(n_1993),
.Y(n_2088)
);

A2O1A1Ixp33_ASAP7_75t_L g2089 ( 
.A1(n_1956),
.A2(n_353),
.B(n_350),
.C(n_351),
.Y(n_2089)
);

AOI21x1_ASAP7_75t_L g2090 ( 
.A1(n_1998),
.A2(n_353),
.B(n_354),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_1962),
.B(n_1926),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1925),
.B(n_2010),
.Y(n_2092)
);

AOI21xp33_ASAP7_75t_SL g2093 ( 
.A1(n_1974),
.A2(n_354),
.B(n_355),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_2014),
.B(n_355),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_2026),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_1950),
.B(n_356),
.Y(n_2096)
);

OAI21xp33_ASAP7_75t_L g2097 ( 
.A1(n_1942),
.A2(n_356),
.B(n_357),
.Y(n_2097)
);

AOI21xp33_ASAP7_75t_L g2098 ( 
.A1(n_1968),
.A2(n_1970),
.B(n_1949),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1979),
.B(n_357),
.Y(n_2099)
);

OAI221xp5_ASAP7_75t_L g2100 ( 
.A1(n_2008),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.C(n_361),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2015),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1937),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2022),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1924),
.Y(n_2104)
);

AOI221x1_ASAP7_75t_SL g2105 ( 
.A1(n_1959),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.C(n_367),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2023),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1927),
.B(n_1921),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2012),
.B(n_368),
.Y(n_2108)
);

HB1xp67_ASAP7_75t_L g2109 ( 
.A(n_2003),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2005),
.B(n_368),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2007),
.B(n_369),
.Y(n_2111)
);

HB1xp67_ASAP7_75t_SL g2112 ( 
.A(n_2105),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2031),
.B(n_1960),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_2033),
.B(n_1966),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_2109),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2035),
.B(n_1953),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2037),
.B(n_2013),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2049),
.B(n_2025),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2046),
.Y(n_2119)
);

NOR2xp33_ASAP7_75t_L g2120 ( 
.A(n_2095),
.B(n_2092),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2039),
.B(n_2047),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2102),
.B(n_2021),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2104),
.B(n_2030),
.Y(n_2123)
);

INVxp67_ASAP7_75t_SL g2124 ( 
.A(n_2084),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2055),
.B(n_2019),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2101),
.B(n_1976),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2103),
.B(n_2106),
.Y(n_2127)
);

INVx1_ASAP7_75t_SL g2128 ( 
.A(n_2107),
.Y(n_2128)
);

BUFx2_ASAP7_75t_L g2129 ( 
.A(n_2046),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2081),
.B(n_2027),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2038),
.Y(n_2131)
);

NAND2x1_ASAP7_75t_L g2132 ( 
.A(n_2034),
.B(n_1941),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2051),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2060),
.B(n_1978),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2088),
.B(n_1967),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2053),
.Y(n_2136)
);

INVx1_ASAP7_75t_SL g2137 ( 
.A(n_2058),
.Y(n_2137)
);

NOR2xp67_ASAP7_75t_SL g2138 ( 
.A(n_2086),
.B(n_1943),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2064),
.Y(n_2139)
);

NOR2x1_ASAP7_75t_L g2140 ( 
.A(n_2043),
.B(n_370),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2091),
.B(n_370),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_SL g2142 ( 
.A(n_2048),
.B(n_562),
.Y(n_2142)
);

NAND2x1_ASAP7_75t_L g2143 ( 
.A(n_2068),
.B(n_568),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2069),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_2074),
.Y(n_2145)
);

OR2x2_ASAP7_75t_L g2146 ( 
.A(n_2063),
.B(n_569),
.Y(n_2146)
);

INVx2_ASAP7_75t_SL g2147 ( 
.A(n_2067),
.Y(n_2147)
);

NOR2x1_ASAP7_75t_L g2148 ( 
.A(n_2082),
.B(n_570),
.Y(n_2148)
);

INVx1_ASAP7_75t_SL g2149 ( 
.A(n_2080),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2098),
.B(n_572),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2115),
.Y(n_2151)
);

BUFx12f_ASAP7_75t_L g2152 ( 
.A(n_2141),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2127),
.Y(n_2153)
);

INVx2_ASAP7_75t_SL g2154 ( 
.A(n_2129),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_2125),
.Y(n_2155)
);

HB1xp67_ASAP7_75t_L g2156 ( 
.A(n_2113),
.Y(n_2156)
);

INVx3_ASAP7_75t_L g2157 ( 
.A(n_2119),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2117),
.Y(n_2158)
);

BUFx2_ASAP7_75t_L g2159 ( 
.A(n_2124),
.Y(n_2159)
);

INVx1_ASAP7_75t_SL g2160 ( 
.A(n_2128),
.Y(n_2160)
);

INVxp67_ASAP7_75t_L g2161 ( 
.A(n_2120),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2131),
.Y(n_2162)
);

HB1xp67_ASAP7_75t_L g2163 ( 
.A(n_2132),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2133),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2136),
.Y(n_2165)
);

INVx1_ASAP7_75t_SL g2166 ( 
.A(n_2145),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2139),
.Y(n_2167)
);

XNOR2xp5_ASAP7_75t_L g2168 ( 
.A(n_2112),
.B(n_2054),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_2116),
.B(n_2032),
.Y(n_2169)
);

BUFx2_ASAP7_75t_L g2170 ( 
.A(n_2134),
.Y(n_2170)
);

INVxp67_ASAP7_75t_SL g2171 ( 
.A(n_2148),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2144),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2143),
.Y(n_2173)
);

AOI221x1_ASAP7_75t_SL g2174 ( 
.A1(n_2151),
.A2(n_2121),
.B1(n_2135),
.B2(n_2114),
.C(n_2118),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_2159),
.B(n_2138),
.Y(n_2175)
);

OAI211xp5_ASAP7_75t_L g2176 ( 
.A1(n_2171),
.A2(n_2040),
.B(n_2085),
.C(n_2045),
.Y(n_2176)
);

OAI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_2168),
.A2(n_2140),
.B(n_2066),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2154),
.B(n_2147),
.Y(n_2178)
);

NAND3xp33_ASAP7_75t_SL g2179 ( 
.A(n_2160),
.B(n_2142),
.C(n_2036),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2161),
.A2(n_2137),
.B1(n_2078),
.B2(n_2149),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_2170),
.A2(n_2079),
.B1(n_2076),
.B2(n_2041),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_SL g2182 ( 
.A1(n_2173),
.A2(n_2056),
.B(n_2071),
.Y(n_2182)
);

NAND4xp25_ASAP7_75t_L g2183 ( 
.A(n_2166),
.B(n_2126),
.C(n_2122),
.D(n_2123),
.Y(n_2183)
);

NAND4xp75_ASAP7_75t_L g2184 ( 
.A(n_2153),
.B(n_2062),
.C(n_2075),
.D(n_2065),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2156),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2157),
.B(n_2130),
.Y(n_2186)
);

NOR3xp33_ASAP7_75t_L g2187 ( 
.A(n_2169),
.B(n_2100),
.C(n_2057),
.Y(n_2187)
);

AOI211xp5_ASAP7_75t_SL g2188 ( 
.A1(n_2176),
.A2(n_2163),
.B(n_2077),
.C(n_2042),
.Y(n_2188)
);

O2A1O1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_2177),
.A2(n_2089),
.B(n_2044),
.C(n_2093),
.Y(n_2189)
);

AOI22xp33_ASAP7_75t_SL g2190 ( 
.A1(n_2175),
.A2(n_2152),
.B1(n_2158),
.B2(n_2155),
.Y(n_2190)
);

OAI221xp5_ASAP7_75t_L g2191 ( 
.A1(n_2174),
.A2(n_2083),
.B1(n_2087),
.B2(n_2150),
.C(n_2097),
.Y(n_2191)
);

NAND4xp25_ASAP7_75t_L g2192 ( 
.A(n_2183),
.B(n_2164),
.C(n_2165),
.D(n_2162),
.Y(n_2192)
);

NOR2xp67_ASAP7_75t_L g2193 ( 
.A(n_2192),
.B(n_2185),
.Y(n_2193)
);

NOR2x1_ASAP7_75t_L g2194 ( 
.A(n_2189),
.B(n_2182),
.Y(n_2194)
);

NOR2xp67_ASAP7_75t_L g2195 ( 
.A(n_2191),
.B(n_2178),
.Y(n_2195)
);

NOR3xp33_ASAP7_75t_L g2196 ( 
.A(n_2190),
.B(n_2186),
.C(n_2187),
.Y(n_2196)
);

NAND2xp33_ASAP7_75t_L g2197 ( 
.A(n_2194),
.B(n_2184),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_R g2198 ( 
.A(n_2193),
.B(n_2090),
.Y(n_2198)
);

AOI21xp5_ASAP7_75t_L g2199 ( 
.A1(n_2197),
.A2(n_2179),
.B(n_2188),
.Y(n_2199)
);

OAI221xp5_ASAP7_75t_L g2200 ( 
.A1(n_2198),
.A2(n_2181),
.B1(n_2196),
.B2(n_2195),
.C(n_2180),
.Y(n_2200)
);

XOR2xp5_ASAP7_75t_L g2201 ( 
.A(n_2199),
.B(n_2108),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2201),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2202),
.A2(n_2200),
.B1(n_2167),
.B2(n_2172),
.Y(n_2203)
);

XNOR2xp5_ASAP7_75t_L g2204 ( 
.A(n_2203),
.B(n_2050),
.Y(n_2204)
);

AOI222xp33_ASAP7_75t_L g2205 ( 
.A1(n_2204),
.A2(n_2094),
.B1(n_2073),
.B2(n_2061),
.C1(n_2070),
.C2(n_2099),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2205),
.Y(n_2206)
);

AOI221xp5_ASAP7_75t_L g2207 ( 
.A1(n_2206),
.A2(n_2052),
.B1(n_2111),
.B2(n_2110),
.C(n_2059),
.Y(n_2207)
);

AOI211xp5_ASAP7_75t_L g2208 ( 
.A1(n_2207),
.A2(n_2146),
.B(n_2096),
.C(n_2072),
.Y(n_2208)
);


endmodule