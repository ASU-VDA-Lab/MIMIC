module fake_jpeg_20261_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_44),
.Y(n_46)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_27),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_54),
.Y(n_96)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_40),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_27),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_27),
.Y(n_55)
);

AO21x1_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_43),
.B(n_40),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_27),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_57),
.B(n_62),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_40),
.Y(n_72)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_27),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_42),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_74),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_47),
.B(n_62),
.C(n_57),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_69),
.B(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_81),
.Y(n_118)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

OR2x2_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_20),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_78),
.B(n_88),
.C(n_91),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_82),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_20),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_85),
.Y(n_126)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_46),
.B(n_42),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_40),
.C(n_60),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_46),
.B(n_26),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_39),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_134)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

OR2x4_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_34),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_101),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_56),
.A2(n_23),
.B1(n_19),
.B2(n_43),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_23),
.B1(n_43),
.B2(n_21),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_40),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_52),
.A2(n_43),
.B1(n_44),
.B2(n_39),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_105),
.A2(n_108),
.B1(n_64),
.B2(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_44),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_107),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_60),
.B(n_17),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_44),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_42),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_122),
.B1(n_131),
.B2(n_82),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_33),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_73),
.B(n_33),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_61),
.B1(n_18),
.B2(n_34),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_78),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_135),
.B1(n_79),
.B2(n_84),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_133),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_73),
.B(n_28),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_136),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_32),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_17),
.A3(n_28),
.B1(n_35),
.B2(n_22),
.Y(n_137)
);

AOI32xp33_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_105),
.A3(n_100),
.B1(n_81),
.B2(n_90),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_89),
.B(n_103),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_139),
.A2(n_150),
.B(n_155),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_106),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_141),
.Y(n_200)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_166),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_153),
.B1(n_158),
.B2(n_161),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_89),
.B(n_87),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_146),
.A2(n_160),
.B(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_149),
.B(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_105),
.B1(n_98),
.B2(n_101),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_105),
.B(n_98),
.C(n_16),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_84),
.B1(n_79),
.B2(n_86),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_167),
.B1(n_71),
.B2(n_16),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_112),
.A2(n_79),
.B1(n_84),
.B2(n_77),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_121),
.B(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_159),
.B(n_169),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_17),
.C(n_35),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_35),
.B1(n_25),
.B2(n_22),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_0),
.B(n_1),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_104),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_165),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_35),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_129),
.C(n_122),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_136),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_110),
.B1(n_137),
.B2(n_126),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_110),
.A2(n_22),
.B1(n_25),
.B2(n_16),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_126),
.B(n_11),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_118),
.B(n_93),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_184),
.C(n_195),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_131),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_187),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_130),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_180),
.B(n_14),
.Y(n_216)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_164),
.C(n_156),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_135),
.B1(n_109),
.B2(n_127),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_185),
.A2(n_188),
.B1(n_194),
.B2(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_109),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_138),
.B1(n_123),
.B2(n_104),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_138),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_199),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_123),
.B1(n_80),
.B2(n_11),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_25),
.C(n_22),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_201),
.B1(n_0),
.B2(n_2),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_25),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_167),
.A2(n_71),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

AND2x4_ASAP7_75t_SL g202 ( 
.A(n_150),
.B(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_202),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_142),
.B1(n_149),
.B2(n_145),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_206),
.B1(n_212),
.B2(n_197),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_162),
.B1(n_168),
.B2(n_145),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_223),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_166),
.B1(n_143),
.B2(n_147),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_211),
.A2(n_195),
.B1(n_172),
.B2(n_186),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_14),
.Y(n_214)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_0),
.B(n_1),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_215),
.A2(n_229),
.B(n_196),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_218),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_184),
.B(n_14),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_220),
.A2(n_194),
.B1(n_171),
.B2(n_188),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_13),
.C(n_12),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_216),
.C(n_215),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_187),
.B(n_2),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_13),
.Y(n_224)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_175),
.B(n_12),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_226),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_192),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_228),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_176),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_8),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_226),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_237),
.B1(n_246),
.B2(n_204),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_198),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_238),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_202),
.B1(n_193),
.B2(n_201),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_218),
.Y(n_238)
);

NAND2x1_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_202),
.Y(n_240)
);

AOI21x1_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_199),
.B(n_191),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_198),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_250),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_222),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_190),
.C(n_180),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_248),
.C(n_223),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_209),
.A2(n_219),
.B1(n_213),
.B2(n_205),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_174),
.C(n_185),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_249),
.A2(n_219),
.B1(n_209),
.B2(n_177),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_174),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_247),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_253),
.A2(n_254),
.B1(n_261),
.B2(n_265),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_221),
.B1(n_208),
.B2(n_179),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_241),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_255),
.B(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_233),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_221),
.B1(n_177),
.B2(n_204),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_263),
.B1(n_230),
.B2(n_242),
.Y(n_272)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_229),
.CI(n_225),
.CON(n_264),
.SN(n_264)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_267),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

AOI22x1_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_171),
.B1(n_220),
.B2(n_191),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_270),
.B1(n_10),
.B2(n_4),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_277),
.B1(n_268),
.B2(n_253),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_238),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_278),
.Y(n_296)
);

NAND5xp2_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_245),
.C(n_234),
.D(n_237),
.E(n_250),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_236),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_280),
.C(n_269),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_233),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_252),
.A2(n_239),
.B(n_224),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_282),
.A2(n_258),
.B(n_264),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_244),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_254),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_290),
.Y(n_303)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_261),
.C(n_264),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_293),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_291),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_274),
.B1(n_271),
.B2(n_276),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_294),
.B1(n_283),
.B2(n_10),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_271),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_277),
.A2(n_268),
.B1(n_4),
.B2(n_5),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_279),
.B(n_278),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_297),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_10),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_298),
.A2(n_290),
.B1(n_6),
.B2(n_7),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_3),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_4),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_3),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_5),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_307),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_310),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_296),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_309),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_304),
.A2(n_286),
.B1(n_296),
.B2(n_7),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_5),
.C(n_6),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_301),
.B(n_305),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_315),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_300),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_316),
.B1(n_314),
.B2(n_311),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_309),
.B(n_299),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_303),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_311),
.B(n_6),
.Y(n_321)
);


endmodule