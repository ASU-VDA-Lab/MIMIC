module real_jpeg_19122_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_36;
wire n_40;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_10),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_2),
.B(n_27),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g22 ( 
.A(n_3),
.B(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_3),
.B(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_13),
.Y(n_12)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g10 ( 
.A1(n_5),
.A2(n_11),
.B(n_14),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

AO21x1_ASAP7_75t_SL g30 ( 
.A1(n_5),
.A2(n_20),
.B(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_7),
.Y(n_6)
);

OAI221xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_22),
.B1(n_24),
.B2(n_31),
.C(n_34),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_16),
.Y(n_8)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

OA21x2_ASAP7_75t_L g27 ( 
.A1(n_11),
.A2(n_14),
.B(n_19),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_15),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B(n_21),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);


endmodule