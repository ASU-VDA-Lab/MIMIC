module fake_jpeg_17099_n_286 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_286);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_286;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_15),
.B1(n_22),
.B2(n_20),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_46),
.B1(n_21),
.B2(n_27),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_15),
.B1(n_22),
.B2(n_20),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

CKINVDCx12_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_36),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_38),
.B(n_25),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_70),
.B(n_78),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_56),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_47),
.B1(n_42),
.B2(n_49),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_68),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_66),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_46),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_17),
.B(n_25),
.C(n_28),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_37),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_21),
.B1(n_32),
.B2(n_23),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_75),
.B1(n_49),
.B2(n_52),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_77),
.Y(n_102)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_23),
.B1(n_25),
.B2(n_17),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_53),
.B(n_30),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_84),
.B1(n_97),
.B2(n_101),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_81),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_42),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_51),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_41),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_25),
.B1(n_8),
.B2(n_11),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_51),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_28),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_57),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_107),
.B(n_118),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_103),
.Y(n_150)
);

AND2x6_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_57),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_61),
.B1(n_76),
.B2(n_17),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_102),
.B1(n_104),
.B2(n_79),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_121),
.B(n_122),
.Y(n_148)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_116),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_85),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_124),
.Y(n_153)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_87),
.B1(n_104),
.B2(n_85),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_30),
.B(n_16),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_61),
.B1(n_65),
.B2(n_77),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_85),
.B1(n_91),
.B2(n_90),
.Y(n_145)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_12),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_11),
.B(n_12),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_66),
.A3(n_24),
.B1(n_18),
.B2(n_65),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_44),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_44),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_101),
.B1(n_100),
.B2(n_96),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_140),
.A2(n_145),
.B1(n_146),
.B2(n_154),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_99),
.C(n_92),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_150),
.C(n_16),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_103),
.B1(n_80),
.B2(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_121),
.B(n_125),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_92),
.B1(n_94),
.B2(n_72),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_16),
.Y(n_155)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_18),
.Y(n_187)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_64),
.B(n_54),
.C(n_2),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_0),
.B(n_1),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_109),
.A2(n_54),
.B1(n_16),
.B2(n_24),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_113),
.B1(n_120),
.B2(n_124),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_166),
.B(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_174),
.Y(n_204)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_131),
.B(n_140),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_159),
.B(n_1),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_144),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_159),
.B(n_152),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_134),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_119),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_148),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_16),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_118),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_184),
.B(n_187),
.Y(n_201)
);

AO22x1_ASAP7_75t_SL g186 ( 
.A1(n_131),
.A2(n_118),
.B1(n_115),
.B2(n_24),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_188),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_199),
.C(n_178),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_143),
.B1(n_151),
.B2(n_160),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_192),
.A2(n_195),
.B1(n_200),
.B2(n_210),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_185),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_193),
.B(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_154),
.Y(n_194)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_151),
.B1(n_146),
.B2(n_145),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_133),
.Y(n_202)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_159),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_161),
.B1(n_183),
.B2(n_172),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_118),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_209),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_191),
.B(n_175),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_214),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_171),
.B1(n_162),
.B2(n_167),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_221),
.B1(n_222),
.B2(n_165),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_181),
.C(n_183),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_226),
.C(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVxp33_ASAP7_75t_SL g234 ( 
.A(n_219),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_161),
.B(n_179),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_220),
.A2(n_206),
.B1(n_184),
.B2(n_186),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_207),
.B1(n_198),
.B2(n_196),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_198),
.B1(n_194),
.B2(n_202),
.Y(n_222)
);

BUFx4f_ASAP7_75t_SL g225 ( 
.A(n_204),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_201),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_163),
.C(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_186),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_166),
.C(n_200),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_231),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_192),
.C(n_170),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_208),
.C(n_163),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_239),
.C(n_177),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_182),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_237),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_236),
.A2(n_227),
.B1(n_224),
.B2(n_212),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_195),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_164),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_223),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_217),
.B1(n_216),
.B2(n_177),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_235),
.B1(n_24),
.B2(n_18),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_28),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_225),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_176),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_239),
.Y(n_254)
);

NAND3xp33_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_180),
.C(n_220),
.Y(n_251)
);

NOR2xp67_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_235),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_238),
.A2(n_176),
.B1(n_174),
.B2(n_173),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_0),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_262),
.C(n_242),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_249),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_261),
.Y(n_263)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_250),
.B1(n_247),
.B2(n_246),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_259),
.A2(n_256),
.B1(n_248),
.B2(n_252),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_267),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_253),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_266),
.B(n_268),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_243),
.Y(n_268)
);

AOI31xp67_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_8),
.A3(n_12),
.B(n_3),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_272),
.A2(n_273),
.B1(n_270),
.B2(n_275),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_7),
.B1(n_10),
.B2(n_3),
.Y(n_273)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_263),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_277),
.A2(n_278),
.B(n_7),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_267),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_9),
.A3(n_10),
.B1(n_5),
.B2(n_6),
.C1(n_1),
.C2(n_2),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_281),
.A2(n_279),
.B(n_5),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_278),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_6),
.B(n_9),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_2),
.B(n_6),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_18),
.Y(n_286)
);


endmodule