module fake_ariane_1769_n_93 (n_8, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_10, n_93);

input n_8;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_10;

output n_93;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_92;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_66;
wire n_71;
wire n_24;
wire n_49;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_23;
wire n_61;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_88;
wire n_68;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_35;
wire n_54;
wire n_25;

BUFx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_7),
.Y(n_28)
);

OAI21x1_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_14),
.B(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

OA21x2_ASAP7_75t_L g38 ( 
.A1(n_0),
.A2(n_1),
.B(n_12),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

AO221x1_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_3),
.B(n_15),
.C(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

OAI21x1_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_29),
.B(n_35),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_29),
.B(n_28),
.Y(n_50)
);

NAND2x1p5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_38),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_39),
.B1(n_34),
.B2(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx2_ASAP7_75t_SL g61 ( 
.A(n_53),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_51),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_52),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_39),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_54),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_66),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_41),
.B1(n_63),
.B2(n_62),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_60),
.Y(n_73)
);

NAND2x1p5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_50),
.B(n_68),
.C(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

NAND4xp25_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_50),
.C(n_48),
.D(n_26),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_79),
.Y(n_82)
);

AOI211xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_49),
.B(n_24),
.C(n_26),
.Y(n_83)
);

NOR4xp25_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_72),
.C(n_35),
.D(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_38),
.C(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_87),
.Y(n_88)
);

AOI221xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_84),
.B1(n_83),
.B2(n_35),
.C(n_31),
.Y(n_89)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_80),
.B1(n_24),
.B2(n_31),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_25),
.B1(n_27),
.B2(n_88),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_90),
.B(n_25),
.Y(n_92)
);

OR2x6_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_25),
.Y(n_93)
);


endmodule