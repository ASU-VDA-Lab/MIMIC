module fake_jpeg_10958_n_397 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_397);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_397;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_45),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_48),
.B(n_54),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_13),
.C(n_11),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_22),
.C(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_60),
.Y(n_115)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_26),
.Y(n_62)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_67),
.B(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_28),
.B(n_0),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_85),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_79),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_76),
.Y(n_127)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_77),
.B(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx2_ASAP7_75t_R g80 ( 
.A(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_15),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_82),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_28),
.B(n_13),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_83),
.B(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_20),
.B(n_11),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_10),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_30),
.B1(n_43),
.B2(n_37),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_89),
.A2(n_93),
.B1(n_96),
.B2(n_108),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_90),
.B(n_114),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_30),
.B1(n_38),
.B2(n_34),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_123),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_30),
.B1(n_38),
.B2(n_34),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_64),
.A2(n_37),
.B1(n_21),
.B2(n_19),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_97),
.A2(n_130),
.B1(n_66),
.B2(n_63),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_107),
.B(n_59),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_32),
.B1(n_42),
.B2(n_79),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_25),
.B(n_35),
.C(n_39),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_109),
.A2(n_76),
.B(n_7),
.C(n_75),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_58),
.B(n_35),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_114),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_69),
.A2(n_37),
.B1(n_21),
.B2(n_32),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_125),
.B1(n_128),
.B2(n_77),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_70),
.B(n_0),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_65),
.A2(n_42),
.B1(n_33),
.B2(n_4),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_33),
.C(n_8),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_133),
.C(n_95),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_SL g133 ( 
.A1(n_71),
.A2(n_8),
.B(n_9),
.Y(n_133)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_62),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_136),
.B(n_144),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_137),
.B(n_162),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_138),
.A2(n_86),
.B1(n_110),
.B2(n_111),
.Y(n_200)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_141),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

BUFx24_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_143),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_62),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_56),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_172),
.B(n_146),
.Y(n_190)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_150),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_66),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_151),
.B(n_166),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_61),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_153),
.B(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_156),
.A2(n_164),
.B1(n_171),
.B2(n_175),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_87),
.B(n_53),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_157),
.B(n_174),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_100),
.Y(n_158)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_165),
.B(n_168),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_87),
.B(n_59),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_126),
.B(n_121),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_170),
.Y(n_215)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_103),
.B(n_82),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_169),
.B(n_131),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_123),
.B(n_9),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_102),
.A2(n_49),
.B1(n_55),
.B2(n_1),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_120),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_7),
.C(n_89),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_92),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_122),
.A2(n_7),
.B1(n_105),
.B2(n_134),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_179),
.B1(n_113),
.B2(n_129),
.Y(n_197)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_178),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_7),
.B1(n_125),
.B2(n_128),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_103),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_141),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_102),
.A2(n_94),
.B1(n_98),
.B2(n_112),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_182),
.B(n_176),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_109),
.A2(n_113),
.B(n_94),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_183),
.B(n_186),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_165),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_152),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_88),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_187),
.B(n_188),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_174),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_155),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_196),
.B(n_206),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_197),
.A2(n_135),
.B1(n_143),
.B2(n_163),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_159),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_142),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_200),
.A2(n_201),
.B1(n_207),
.B2(n_164),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_138),
.A2(n_86),
.B1(n_110),
.B2(n_129),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_137),
.B(n_131),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_111),
.B1(n_149),
.B2(n_179),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_149),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_212),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_213),
.B(n_218),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_160),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_177),
.A2(n_168),
.B(n_140),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_141),
.B(n_142),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_150),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_224),
.B(n_214),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_225),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_226),
.B(n_227),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_221),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_239),
.C(n_259),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_145),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_230),
.B(n_235),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_231),
.A2(n_234),
.B(n_184),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_183),
.B(n_162),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_236),
.B(n_243),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_175),
.C(n_139),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_249),
.B1(n_253),
.B2(n_203),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_221),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_245),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_242),
.A2(n_247),
.B1(n_248),
.B2(n_252),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_202),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_223),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_246),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_197),
.B1(n_208),
.B2(n_220),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_207),
.B1(n_186),
.B2(n_206),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_188),
.A2(n_210),
.B1(n_187),
.B2(n_201),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_215),
.B(n_217),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_200),
.A2(n_185),
.B1(n_191),
.B2(n_220),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_193),
.B(n_185),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_193),
.A2(n_209),
.B1(n_219),
.B2(n_222),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_256),
.A2(n_209),
.B1(n_199),
.B2(n_195),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_198),
.B(n_202),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_260),
.A2(n_272),
.B1(n_283),
.B2(n_268),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_261),
.A2(n_286),
.B1(n_271),
.B2(n_268),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_204),
.C(n_211),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_273),
.C(n_275),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_247),
.A2(n_222),
.B1(n_195),
.B2(n_204),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_204),
.C(n_184),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_276),
.B(n_278),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_205),
.C(n_192),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_249),
.A2(n_205),
.B1(n_192),
.B2(n_194),
.Y(n_276)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_277),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_255),
.A2(n_194),
.B(n_231),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_229),
.C(n_239),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_262),
.C(n_286),
.Y(n_311)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_257),
.B(n_242),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_245),
.B(n_243),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_234),
.A2(n_254),
.B1(n_237),
.B2(n_238),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_287),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_259),
.Y(n_290)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_227),
.Y(n_291)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_291),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_237),
.B1(n_256),
.B2(n_241),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_295),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_252),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_296),
.B(n_299),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

BUFx12_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_233),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_232),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_309),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_271),
.B(n_228),
.Y(n_303)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_303),
.Y(n_322)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_279),
.B(n_283),
.Y(n_306)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_308),
.A2(n_290),
.B1(n_265),
.B2(n_276),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_279),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_310),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_280),
.C(n_262),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_281),
.B(n_284),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_314),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_288),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_263),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_294),
.B(n_304),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_325),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_332),
.C(n_336),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_275),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_334),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_309),
.C(n_292),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_314),
.A2(n_273),
.B1(n_274),
.B2(n_278),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_333),
.B(n_293),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_260),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_264),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_299),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_338),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_319),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_SL g363 ( 
.A(n_339),
.B(n_345),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_326),
.Y(n_340)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_341),
.Y(n_355)
);

OAI321xp33_ASAP7_75t_L g343 ( 
.A1(n_327),
.A2(n_306),
.A3(n_310),
.B1(n_303),
.B2(n_308),
.C(n_305),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_343),
.B(n_344),
.Y(n_360)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_318),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_326),
.B(n_312),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_325),
.B(n_293),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_348),
.A2(n_329),
.B(n_316),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_312),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_349),
.A2(n_350),
.B1(n_351),
.B2(n_316),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_324),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_322),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_328),
.C(n_334),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_352),
.B(n_353),
.C(n_323),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_301),
.C(n_264),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_348),
.A2(n_333),
.B1(n_329),
.B2(n_323),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_357),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_358),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_317),
.C(n_301),
.Y(n_357)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_361),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_342),
.A2(n_335),
.B1(n_330),
.B2(n_320),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_364),
.B(n_366),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_342),
.A2(n_307),
.B1(n_294),
.B2(n_320),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_365),
.A2(n_338),
.B1(n_282),
.B2(n_263),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_341),
.A2(n_315),
.B1(n_297),
.B2(n_282),
.Y(n_366)
);

NAND2x1_ASAP7_75t_SL g367 ( 
.A(n_357),
.B(n_353),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_369),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_362),
.Y(n_369)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_370),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_355),
.A2(n_359),
.B1(n_360),
.B2(n_356),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_371),
.A2(n_366),
.B1(n_358),
.B2(n_298),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_355),
.A2(n_347),
.B1(n_346),
.B2(n_266),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_374),
.B(n_354),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_363),
.B(n_347),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_375),
.B(n_372),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_364),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_377),
.B(n_379),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_378),
.Y(n_386)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_368),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_346),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_383),
.C(n_376),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_382),
.A2(n_367),
.B(n_298),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_387),
.B(n_384),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_371),
.C(n_373),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_388),
.B(n_389),
.C(n_378),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g393 ( 
.A(n_390),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_391),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_381),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_393),
.B(n_392),
.C(n_386),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_394),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_396),
.B(n_298),
.Y(n_397)
);


endmodule