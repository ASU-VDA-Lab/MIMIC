module fake_jpeg_21929_n_325 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_34),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_44),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_48),
.B(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_27),
.B1(n_19),
.B2(n_17),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_17),
.B1(n_27),
.B2(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_36),
.C(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_28),
.A2(n_19),
.B1(n_17),
.B2(n_27),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_37),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_56),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_43),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_58),
.B(n_62),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_59),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_37),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_19),
.B1(n_27),
.B2(n_35),
.Y(n_82)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_50),
.B1(n_47),
.B2(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx2_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_16),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_48),
.B1(n_51),
.B2(n_42),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_81),
.B1(n_82),
.B2(n_85),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_48),
.B1(n_53),
.B2(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_60),
.A2(n_45),
.B1(n_38),
.B2(n_46),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_92),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_73),
.B(n_66),
.Y(n_114)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_49),
.C(n_40),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_53),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_41),
.Y(n_101)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_45),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_35),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_97),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_75),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_63),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_108),
.Y(n_140)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_117),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_67),
.B1(n_63),
.B2(n_96),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_113),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_114),
.A2(n_115),
.B(n_91),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_76),
.B(n_82),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

OR2x2_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_71),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_81),
.B(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_78),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_129),
.B(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_98),
.B1(n_84),
.B2(n_89),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_133),
.B1(n_138),
.B2(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_128),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_67),
.B1(n_111),
.B2(n_106),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_86),
.B1(n_65),
.B2(n_52),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_136),
.B1(n_31),
.B2(n_59),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_83),
.B1(n_96),
.B2(n_80),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_71),
.B(n_74),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_141),
.B(n_14),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_86),
.B1(n_55),
.B2(n_56),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_109),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_105),
.A2(n_77),
.B1(n_80),
.B2(n_78),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_134),
.C(n_101),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_74),
.B(n_86),
.Y(n_141)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_74),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_69),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_149),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_170),
.C(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_119),
.B1(n_103),
.B2(n_106),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_152),
.A2(n_159),
.B(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_162),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_99),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_155),
.B(n_161),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_156),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_112),
.B1(n_21),
.B2(n_20),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_14),
.B1(n_167),
.B2(n_162),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_100),
.Y(n_160)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_125),
.B(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_112),
.Y(n_164)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_69),
.Y(n_166)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_126),
.B(n_138),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_88),
.C(n_31),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_173),
.B1(n_127),
.B2(n_122),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_172),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_129),
.A2(n_68),
.B1(n_59),
.B2(n_34),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_190),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_135),
.B1(n_136),
.B2(n_124),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_172),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_168),
.Y(n_203)
);

XNOR2x2_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_143),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_184),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_141),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_196),
.C(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_135),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_198),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_68),
.B1(n_25),
.B2(n_23),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_151),
.A2(n_13),
.B1(n_26),
.B2(n_24),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_13),
.B1(n_26),
.B2(n_24),
.Y(n_192)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_18),
.C(n_16),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_163),
.A2(n_25),
.B1(n_21),
.B2(n_23),
.Y(n_197)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_161),
.B(n_18),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_211),
.C(n_214),
.Y(n_241)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_193),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_209),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_164),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_154),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_187),
.B(n_167),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_212),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_166),
.C(n_160),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_155),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_180),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_153),
.C(n_149),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_146),
.B(n_148),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_177),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_148),
.Y(n_221)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_16),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_227),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_204),
.A2(n_178),
.B1(n_177),
.B2(n_175),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_231),
.B1(n_235),
.B2(n_208),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_188),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_189),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_199),
.B1(n_200),
.B2(n_184),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_196),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_242),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_217),
.A2(n_222),
.B1(n_205),
.B2(n_223),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_174),
.C(n_190),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_236),
.B(n_16),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_217),
.A2(n_171),
.B1(n_173),
.B2(n_154),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_197),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_219),
.A2(n_25),
.B1(n_21),
.B2(n_23),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_220),
.B1(n_222),
.B2(n_203),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_211),
.C(n_201),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_241),
.C(n_227),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_255),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_202),
.Y(n_249)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_218),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_256),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_252),
.A2(n_247),
.B1(n_240),
.B2(n_258),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_239),
.B(n_228),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_253),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_214),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_234),
.A2(n_220),
.B1(n_34),
.B2(n_32),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_261),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_226),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_229),
.B(n_10),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_259),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_30),
.B1(n_29),
.B2(n_2),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_233),
.B(n_12),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_262),
.A2(n_26),
.B1(n_24),
.B2(n_12),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_268),
.C(n_272),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_250),
.C(n_263),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_246),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_1),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_271),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_236),
.C(n_244),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_273),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_11),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_275),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_11),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_0),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_272),
.A2(n_256),
.B(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_252),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_285),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_267),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_292),
.B(n_293),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_290),
.B(n_268),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_18),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_286),
.B(n_289),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

XNOR2x2_ASAP7_75t_SL g290 ( 
.A(n_266),
.B(n_270),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_269),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_1),
.B(n_2),
.Y(n_293)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_8),
.C(n_9),
.Y(n_311)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_303),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_278),
.C(n_279),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_4),
.C(n_5),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_281),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_3),
.B(n_4),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_9),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_300),
.A2(n_284),
.B1(n_5),
.B2(n_6),
.Y(n_305)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_310),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_302),
.B1(n_298),
.B2(n_297),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_312),
.B(n_295),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_306),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.C(n_315),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_307),
.C(n_311),
.Y(n_318)
);

NAND3xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_314),
.C(n_9),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

A2O1A1O1Ixp25_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_9),
.B(n_16),
.C(n_22),
.D(n_306),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_22),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_22),
.C(n_156),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_22),
.B(n_298),
.Y(n_325)
);


endmodule