module fake_aes_10593_n_41 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
INVx1_ASAP7_75t_SL g14 ( .A(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_15), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_12), .B(n_0), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_17), .B(n_2), .Y(n_22) );
BUFx3_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_19), .B(n_18), .Y(n_24) );
INVx1_ASAP7_75t_SL g25 ( .A(n_23), .Y(n_25) );
OAI222xp33_ASAP7_75t_L g26 ( .A1(n_22), .A2(n_17), .B1(n_14), .B2(n_13), .C1(n_5), .C2(n_2), .Y(n_26) );
OAI21xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_20), .B(n_19), .Y(n_27) );
NAND3xp33_ASAP7_75t_SL g28 ( .A(n_25), .B(n_20), .C(n_23), .Y(n_28) );
OAI221xp5_ASAP7_75t_L g29 ( .A1(n_24), .A2(n_21), .B1(n_4), .B2(n_5), .C(n_3), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
INVxp67_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
NOR2xp33_ASAP7_75t_L g33 ( .A(n_30), .B(n_26), .Y(n_33) );
AOI321xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_21), .A3(n_30), .B1(n_3), .B2(n_28), .C(n_25), .Y(n_34) );
AND2x2_ASAP7_75t_SL g35 ( .A(n_32), .B(n_21), .Y(n_35) );
AOI21xp33_ASAP7_75t_SL g36 ( .A1(n_33), .A2(n_21), .B(n_8), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_35), .Y(n_37) );
XNOR2xp5_ASAP7_75t_L g38 ( .A(n_35), .B(n_6), .Y(n_38) );
INVx1_ASAP7_75t_L g39 ( .A(n_34), .Y(n_39) );
INVxp33_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
OAI221xp5_ASAP7_75t_R g41 ( .A1(n_40), .A2(n_39), .B1(n_37), .B2(n_36), .C(n_9), .Y(n_41) );
endmodule