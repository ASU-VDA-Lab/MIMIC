module fake_jpeg_13882_n_502 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_50),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_56),
.Y(n_97)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_58),
.Y(n_143)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_27),
.B(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_76),
.Y(n_110)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_85),
.Y(n_121)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g81 ( 
.A(n_38),
.Y(n_81)
);

CKINVDCx9p33_ASAP7_75t_R g119 ( 
.A(n_81),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_84),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_22),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g138 ( 
.A(n_92),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_18),
.B(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_41),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_40),
.B(n_22),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_102),
.B(n_20),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_27),
.B1(n_31),
.B2(n_47),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_114),
.A2(n_32),
.B1(n_27),
.B2(n_31),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_18),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_128),
.B(n_129),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_81),
.A2(n_41),
.B(n_48),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_132),
.B(n_133),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_92),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_60),
.B(n_45),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_69),
.B(n_43),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_135),
.B(n_137),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_63),
.B(n_43),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_86),
.B(n_44),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_86),
.B(n_44),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_34),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_153),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_84),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_34),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_156),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_51),
.B(n_28),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_157),
.Y(n_238)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_158),
.Y(n_244)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_159),
.Y(n_241)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_102),
.A2(n_72),
.B(n_73),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_162),
.A2(n_182),
.B(n_199),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_121),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_163),
.B(n_177),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_165),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_110),
.A2(n_89),
.B1(n_93),
.B2(n_64),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_167),
.A2(n_170),
.B1(n_145),
.B2(n_98),
.Y(n_227)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_115),
.Y(n_174)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_174),
.Y(n_259)
);

CKINVDCx12_ASAP7_75t_R g175 ( 
.A(n_108),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_175),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_116),
.A2(n_40),
.B1(n_21),
.B2(n_87),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_176),
.A2(n_185),
.B1(n_198),
.B2(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_125),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_201),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_97),
.B(n_95),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_181),
.B(n_205),
.Y(n_235)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_116),
.A2(n_40),
.B1(n_21),
.B2(n_28),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_25),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_213),
.Y(n_215)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_193),
.Y(n_232)
);

CKINVDCx12_ASAP7_75t_R g191 ( 
.A(n_113),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_191),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_113),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_192),
.B(n_196),
.Y(n_231)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_118),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_194),
.B(n_195),
.Y(n_258)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_131),
.B(n_42),
.Y(n_196)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_99),
.A2(n_57),
.B1(n_70),
.B2(n_31),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_125),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_204),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_107),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_203),
.B(n_208),
.Y(n_254)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_143),
.B(n_25),
.Y(n_205)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_125),
.A2(n_88),
.B1(n_83),
.B2(n_82),
.Y(n_206)
);

OA22x2_ASAP7_75t_SL g261 ( 
.A1(n_206),
.A2(n_209),
.B1(n_4),
.B2(n_5),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_99),
.A2(n_80),
.B1(n_49),
.B2(n_42),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_207),
.A2(n_103),
.B(n_6),
.Y(n_262)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_140),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_210),
.B(n_212),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_143),
.B(n_16),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_107),
.B(n_16),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_147),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_214),
.A2(n_208),
.B1(n_195),
.B2(n_127),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_182),
.A2(n_140),
.B1(n_151),
.B2(n_150),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_216),
.A2(n_236),
.B1(n_241),
.B2(n_233),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_154),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_233),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_152),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_221),
.B(n_226),
.C(n_228),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_162),
.A2(n_147),
.B(n_136),
.C(n_139),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_225),
.A2(n_201),
.B(n_7),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_152),
.C(n_122),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_262),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_180),
.B(n_127),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_154),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_200),
.A2(n_145),
.B1(n_120),
.B2(n_109),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_234),
.A2(n_243),
.B1(n_246),
.B2(n_260),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_170),
.B1(n_209),
.B2(n_174),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_207),
.A2(n_199),
.B1(n_179),
.B2(n_196),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_173),
.B(n_130),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_249),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_120),
.B1(n_130),
.B2(n_98),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_193),
.B(n_122),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_206),
.A2(n_136),
.B1(n_139),
.B2(n_14),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_209),
.B1(n_198),
.B2(n_168),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_194),
.B(n_4),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_4),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_158),
.B(n_165),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_264),
.A2(n_271),
.B(n_282),
.Y(n_333)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_265),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_187),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_266),
.B(n_275),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_209),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_291),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_231),
.A2(n_184),
.B(n_189),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_272),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_257),
.Y(n_273)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_254),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_274),
.B(n_296),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_210),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_276),
.B(n_299),
.C(n_259),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_172),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_277),
.B(n_295),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_278),
.A2(n_285),
.B1(n_290),
.B2(n_244),
.Y(n_309)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_280),
.A2(n_292),
.B1(n_304),
.B2(n_229),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_216),
.A2(n_159),
.B(n_157),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_218),
.A2(n_157),
.B(n_186),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_300),
.B(n_305),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_236),
.A2(n_164),
.B1(n_183),
.B2(n_190),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_286),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_225),
.A2(n_204),
.B(n_211),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_287),
.A2(n_298),
.B(n_302),
.Y(n_312)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_219),
.Y(n_289)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_171),
.B1(n_103),
.B2(n_201),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_215),
.B(n_14),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_261),
.A2(n_103),
.B1(n_7),
.B2(n_8),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

AND2x6_ASAP7_75t_L g294 ( 
.A(n_228),
.B(n_6),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_297),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_215),
.B(n_6),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_258),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_245),
.B(n_6),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_242),
.A2(n_11),
.B(n_8),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_226),
.B(n_7),
.C(n_9),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_239),
.B(n_11),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_222),
.B(n_11),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_307),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_232),
.B(n_9),
.Y(n_302)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_308),
.B1(n_248),
.B2(n_217),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_263),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_230),
.A2(n_10),
.B(n_244),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_258),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_302),
.B1(n_269),
.B2(n_281),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_223),
.B(n_10),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_248),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_313),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_278),
.A2(n_285),
.B1(n_269),
.B2(n_290),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_L g350 ( 
.A1(n_314),
.A2(n_302),
.B(n_283),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_276),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_315),
.B(n_323),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_270),
.A2(n_247),
.B1(n_239),
.B2(n_224),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_316),
.A2(n_322),
.B1(n_331),
.B2(n_332),
.Y(n_360)
);

AOI32xp33_ASAP7_75t_L g317 ( 
.A1(n_288),
.A2(n_253),
.A3(n_247),
.B1(n_232),
.B2(n_258),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_337),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_318),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_232),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_330),
.Y(n_365)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_321),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_280),
.A2(n_240),
.B1(n_217),
.B2(n_251),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_267),
.B(n_252),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_251),
.B(n_252),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_329),
.A2(n_338),
.B(n_300),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_267),
.B(n_220),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_270),
.A2(n_273),
.B1(n_293),
.B2(n_272),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_293),
.A2(n_220),
.B1(n_259),
.B2(n_237),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_334),
.A2(n_347),
.B1(n_268),
.B2(n_294),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_287),
.B(n_288),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_340),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_271),
.B(n_237),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_344),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_229),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_265),
.Y(n_346)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_346),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_268),
.A2(n_294),
.B1(n_269),
.B2(n_277),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_348),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_350),
.A2(n_336),
.B1(n_314),
.B2(n_311),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_325),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_371),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_335),
.B(n_275),
.Y(n_358)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_266),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_359),
.B(n_362),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_301),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_363),
.A2(n_327),
.B(n_312),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_330),
.B(n_297),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_364),
.B(n_378),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_326),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_307),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_367),
.B(n_375),
.Y(n_401)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_326),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_368),
.Y(n_383)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_369),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_328),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_316),
.B(n_323),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_376),
.Y(n_402)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_311),
.Y(n_373)
);

A2O1A1Ixp33_ASAP7_75t_SL g384 ( 
.A1(n_373),
.A2(n_333),
.B(n_303),
.C(n_329),
.Y(n_384)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_346),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_374),
.B(n_377),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_320),
.B(n_291),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_340),
.B(n_295),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_341),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_300),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_380),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_338),
.B(n_304),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_324),
.B(n_308),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_381),
.B(n_345),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_319),
.C(n_315),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_386),
.C(n_404),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_384),
.B(n_406),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_337),
.C(n_342),
.Y(n_386)
);

NOR3xp33_ASAP7_75t_SL g387 ( 
.A(n_380),
.B(n_324),
.C(n_310),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_387),
.B(n_378),
.Y(n_420)
);

AO22x1_ASAP7_75t_L g388 ( 
.A1(n_363),
.A2(n_336),
.B1(n_327),
.B2(n_333),
.Y(n_388)
);

OAI31xp33_ASAP7_75t_SL g426 ( 
.A1(n_388),
.A2(n_373),
.A3(n_354),
.B(n_353),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_365),
.B(n_347),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_389),
.B(n_409),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_310),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_396),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_397),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_313),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_403),
.B(n_407),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_357),
.B(n_309),
.C(n_312),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_349),
.A2(n_298),
.B1(n_282),
.B2(n_279),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_405),
.A2(n_396),
.B1(n_406),
.B2(n_360),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_361),
.A2(n_279),
.B(n_349),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_358),
.B(n_376),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_364),
.B(n_352),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_408),
.B(n_377),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_357),
.B(n_351),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_395),
.Y(n_411)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_411),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_398),
.A2(n_372),
.B1(n_361),
.B2(n_379),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_414),
.A2(n_427),
.B1(n_428),
.B2(n_405),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_356),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_423),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_383),
.Y(n_416)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_416),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_401),
.A2(n_360),
.B1(n_398),
.B2(n_392),
.Y(n_418)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_418),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_422),
.B1(n_384),
.B2(n_388),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_420),
.A2(n_383),
.B1(n_373),
.B2(n_366),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_421),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_404),
.A2(n_353),
.B1(n_354),
.B2(n_369),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_395),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_426),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_385),
.B(n_356),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_385),
.B(n_366),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_394),
.B(n_374),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_429),
.B(n_430),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_355),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_386),
.B(n_382),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_433),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_390),
.Y(n_433)
);

INVx11_ASAP7_75t_L g434 ( 
.A(n_426),
.Y(n_434)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_431),
.B(n_391),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_445),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_412),
.B(n_389),
.C(n_409),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_442),
.B(n_443),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_384),
.C(n_397),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_384),
.C(n_402),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_447),
.C(n_449),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_432),
.B(n_388),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_446),
.A2(n_414),
.B1(n_413),
.B2(n_416),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_432),
.C(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_448),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_355),
.C(n_387),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_450),
.B(n_419),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_441),
.B1(n_451),
.B2(n_437),
.Y(n_453)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_440),
.B(n_430),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_435),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_455),
.A2(n_459),
.B1(n_425),
.B2(n_399),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_447),
.B(n_424),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_SL g471 ( 
.A(n_456),
.B(n_463),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_434),
.Y(n_459)
);

FAx1_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_443),
.CI(n_449),
.CON(n_460),
.SN(n_460)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_445),
.Y(n_468)
);

BUFx12_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_410),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_464),
.A2(n_425),
.B(n_442),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_465),
.A2(n_435),
.B1(n_399),
.B2(n_368),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_438),
.B(n_413),
.C(n_429),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_467),
.C(n_457),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_470),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_458),
.A2(n_439),
.B1(n_413),
.B2(n_433),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_472),
.B(n_473),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_474),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_477),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_458),
.A2(n_368),
.B1(n_436),
.B2(n_462),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_476),
.B(n_478),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_466),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_478),
.B(n_461),
.Y(n_479)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_479),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_461),
.C(n_465),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_481),
.B(n_471),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_460),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_482),
.A2(n_469),
.B(n_472),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_487),
.B(n_490),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_489),
.A2(n_483),
.B(n_484),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_470),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_476),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_491),
.B(n_481),
.Y(n_493)
);

OAI21x1_ASAP7_75t_SL g495 ( 
.A1(n_493),
.A2(n_494),
.B(n_488),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_495),
.B(n_496),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_492),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_497),
.Y(n_498)
);

AOI321xp33_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_454),
.A3(n_486),
.B1(n_460),
.B2(n_483),
.C(n_475),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_499),
.B(n_463),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_500),
.Y(n_501)
);

AO21x1_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_463),
.B(n_456),
.Y(n_502)
);


endmodule