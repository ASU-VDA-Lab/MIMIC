module fake_netlist_5_2561_n_131 (n_16, n_0, n_12, n_9, n_18, n_22, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_131);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_131;

wire n_91;
wire n_82;
wire n_122;
wire n_24;
wire n_124;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_114;
wire n_96;
wire n_57;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_128;
wire n_73;
wire n_92;
wire n_120;
wire n_30;
wire n_33;
wire n_126;
wire n_84;
wire n_23;
wire n_130;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_118;
wire n_28;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_21),
.Y(n_23)
);

INVxp67_ASAP7_75t_SL g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NAND2x1p5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

AO21x2_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_35),
.B(n_23),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_52),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_49),
.B(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_52),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_48),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_60),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_55),
.Y(n_77)
);

O2A1O1Ixp5_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_49),
.B(n_42),
.C(n_41),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_58),
.B1(n_25),
.B2(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_48),
.Y(n_80)
);

AOI221x1_ASAP7_75t_SL g81 ( 
.A1(n_66),
.A2(n_43),
.B1(n_36),
.B2(n_27),
.C(n_45),
.Y(n_81)
);

AOI21x1_ASAP7_75t_SL g82 ( 
.A1(n_64),
.A2(n_46),
.B(n_49),
.Y(n_82)
);

AO21x2_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_73),
.B(n_74),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_64),
.B1(n_65),
.B2(n_41),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_90),
.A2(n_78),
.B(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_66),
.B(n_43),
.Y(n_96)
);

OA21x2_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_66),
.B(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_81),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_102),
.A2(n_93),
.B(n_83),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_64),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_46),
.B1(n_97),
.B2(n_71),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_71),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_83),
.B(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_91),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_91),
.Y(n_114)
);

OAI221xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_41),
.B1(n_42),
.B2(n_49),
.C(n_46),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_96),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_42),
.B(n_91),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_97),
.B(n_57),
.C(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_106),
.B(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_105),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_SL g123 ( 
.A(n_121),
.B(n_107),
.C(n_118),
.Y(n_123)
);

OR3x1_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_0),
.C(n_1),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

OAI221xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_122),
.B1(n_57),
.B2(n_4),
.C(n_5),
.Y(n_126)
);

OAI322xp33_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_1),
.A3(n_3),
.B1(n_5),
.B2(n_91),
.C1(n_63),
.C2(n_8),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_123),
.B1(n_127),
.B2(n_97),
.Y(n_129)
);

NAND4xp25_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_63),
.C(n_7),
.D(n_10),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_63),
.B1(n_16),
.B2(n_17),
.Y(n_131)
);


endmodule