module fake_jpeg_5070_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_1),
.B(n_0),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx24_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_10),
.B1(n_7),
.B2(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_14),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_8),
.B(n_5),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_10),
.B1(n_6),
.B2(n_5),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_16),
.B(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_16),
.B(n_17),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_18),
.B1(n_7),
.B2(n_9),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_16),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_11),
.B1(n_13),
.B2(n_2),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_11),
.C(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_11),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_33),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_30),
.C(n_31),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_35),
.Y(n_36)
);

AOI322xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_0),
.A3(n_1),
.B1(n_3),
.B2(n_4),
.C1(n_34),
.C2(n_32),
.Y(n_37)
);

AOI221xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.C(n_20),
.Y(n_38)
);


endmodule