module fake_jpeg_17572_n_208 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_1),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_15),
.B(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_58),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_35),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_31),
.B1(n_30),
.B2(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_19),
.B1(n_15),
.B2(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_30),
.B1(n_31),
.B2(n_24),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_62),
.B(n_22),
.Y(n_75)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_28),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_63),
.A2(n_43),
.B(n_51),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_71),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_36),
.Y(n_69)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_75),
.A2(n_82),
.B1(n_68),
.B2(n_45),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_56),
.B1(n_59),
.B2(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_55),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_20),
.B(n_16),
.C(n_26),
.Y(n_82)
);

AO22x1_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_20),
.B1(n_50),
.B2(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_101),
.B(n_20),
.Y(n_122)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_80),
.B1(n_77),
.B2(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_97),
.Y(n_112)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_63),
.B(n_22),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_21),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_70),
.B1(n_16),
.B2(n_26),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_44),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_110),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_63),
.B1(n_75),
.B2(n_82),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_109),
.B1(n_117),
.B2(n_119),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_65),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_123),
.C(n_22),
.Y(n_135)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_115),
.B(n_120),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_99),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_79),
.B1(n_44),
.B2(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_53),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_86),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_26),
.B1(n_21),
.B2(n_28),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_92),
.B(n_5),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_20),
.B(n_28),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_88),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_88),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_135),
.C(n_139),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_90),
.B(n_53),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_128),
.B(n_140),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_143),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_132),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_115),
.B(n_116),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

AOI221xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_20),
.B1(n_21),
.B2(n_28),
.C(n_25),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_138),
.C(n_38),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

NOR4xp25_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_53),
.C(n_87),
.D(n_38),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_113),
.C(n_118),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_92),
.B(n_38),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_131),
.Y(n_146)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_117),
.C(n_124),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_159),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_153),
.B(n_156),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_154),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_130),
.B(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_128),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_37),
.C(n_38),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_138),
.B(n_133),
.C(n_139),
.D(n_142),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_160),
.A2(n_158),
.B(n_155),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_140),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_171),
.C(n_172),
.Y(n_173)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_97),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_142),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_25),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_159),
.C(n_144),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_178),
.C(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_148),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_165),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_144),
.B(n_154),
.C(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_161),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_78),
.C(n_28),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_183),
.A2(n_187),
.B(n_4),
.C(n_7),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_180),
.B(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_171),
.B1(n_172),
.B2(n_162),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_174),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_96),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_25),
.C(n_18),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_181),
.A3(n_173),
.B1(n_182),
.B2(n_12),
.C1(n_14),
.C2(n_13),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_8),
.B(n_9),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_186),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_194),
.A2(n_8),
.B(n_9),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_14),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_200),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_201),
.C(n_18),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_194),
.B1(n_196),
.B2(n_10),
.Y(n_202)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_204),
.B(n_203),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_203),
.A2(n_10),
.B(n_11),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_18),
.Y(n_208)
);


endmodule