module fake_ariane_306_n_1496 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_323, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_39, n_155, n_127, n_1496);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_323;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1496;

wire n_913;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_1495;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_272),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_8),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_38),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_256),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_156),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_137),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_192),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_244),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_318),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_67),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_35),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_148),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_215),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_285),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_93),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_2),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_149),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_310),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_154),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_186),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_304),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_125),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_266),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_200),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_66),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_15),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_115),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_100),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_312),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_229),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_55),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_5),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_214),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_164),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_194),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_224),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_150),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_21),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_64),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_21),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_123),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_240),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_237),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_120),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_283),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_29),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_136),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_257),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_27),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_174),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_295),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_265),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_6),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_168),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_27),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_177),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_104),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_254),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_264),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_30),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_238),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_92),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_179),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_23),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_54),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_213),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_276),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_16),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_199),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_321),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_25),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

BUFx10_ASAP7_75t_L g400 ( 
.A(n_222),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_323),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_53),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_259),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_89),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_217),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_113),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_53),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_223),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_165),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_294),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_195),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_24),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_277),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_231),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_267),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_178),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_144),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_227),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_212),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_274),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_261),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_26),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_119),
.Y(n_424)
);

BUFx8_ASAP7_75t_SL g425 ( 
.A(n_64),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_3),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_25),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_151),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_41),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_303),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_26),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_2),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_55),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_139),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_203),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_302),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_44),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_34),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_306),
.Y(n_439)
);

BUFx10_ASAP7_75t_L g440 ( 
.A(n_43),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_142),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_0),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_278),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_286),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_114),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_91),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_196),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_1),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_191),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_298),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_249),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_107),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_201),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_57),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_218),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_133),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_116),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_92),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_117),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_170),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_202),
.Y(n_461)
);

BUFx10_ASAP7_75t_L g462 ( 
.A(n_24),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_88),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_287),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_84),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_77),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_155),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_34),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_22),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_145),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_305),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_138),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_275),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_9),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_316),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_66),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_247),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_172),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_233),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_234),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_311),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_44),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_72),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_103),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_181),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_43),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_3),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_288),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_171),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_293),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_61),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_307),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_128),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_219),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_205),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_86),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_166),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_129),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_93),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_159),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_268),
.Y(n_501)
);

BUFx8_ASAP7_75t_SL g502 ( 
.A(n_169),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_248),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_270),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_309),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_314),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_35),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_134),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_141),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_96),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_300),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_60),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_180),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_230),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_198),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_226),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_252),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_255),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_78),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_130),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_91),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_161),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_5),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_109),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_106),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_9),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_22),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_86),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_251),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_152),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_188),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_99),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_153),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_162),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_246),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_206),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_62),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_301),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_140),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_111),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_70),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_51),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_60),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_29),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_253),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_241),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_0),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_121),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_320),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_110),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_87),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_208),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_282),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_426),
.B(n_1),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_327),
.B(n_402),
.Y(n_555)
);

AND2x6_ASAP7_75t_L g556 ( 
.A(n_329),
.B(n_97),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_400),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_468),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_327),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_329),
.B(n_98),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_336),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_337),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_400),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_343),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_4),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_388),
.B(n_4),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_400),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_494),
.B(n_6),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_326),
.B(n_7),
.Y(n_570)
);

BUFx12f_ASAP7_75t_L g571 ( 
.A(n_509),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_425),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_509),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_331),
.B(n_7),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_440),
.B(n_8),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_402),
.B(n_10),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_509),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_342),
.Y(n_578)
);

BUFx12f_ASAP7_75t_L g579 ( 
.A(n_440),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_339),
.B(n_10),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_342),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_340),
.B(n_11),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_547),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_344),
.B(n_11),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_521),
.B(n_12),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_345),
.B(n_12),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_440),
.B(n_13),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_502),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_521),
.B(n_13),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_347),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_342),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_352),
.B(n_14),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_333),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_462),
.B(n_14),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_363),
.B(n_15),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_462),
.B(n_16),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_347),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_353),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_539),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_371),
.B(n_17),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_352),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_342),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_365),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_374),
.B(n_17),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_458),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_458),
.B(n_18),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_381),
.B(n_18),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_539),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_373),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_333),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_376),
.B(n_19),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_380),
.Y(n_612)
);

CKINVDCx11_ASAP7_75t_R g613 ( 
.A(n_499),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_386),
.B(n_19),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_462),
.B(n_20),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_539),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_334),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_396),
.B(n_20),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_399),
.B(n_23),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_405),
.B(n_28),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_547),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_551),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_409),
.B(n_28),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_403),
.B(n_30),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_334),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_412),
.B(n_31),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_551),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_476),
.B(n_31),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_382),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_476),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_539),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_502),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_328),
.Y(n_634)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_358),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_356),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_356),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_360),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_349),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_389),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_360),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_479),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_417),
.B(n_32),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_420),
.B(n_32),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_479),
.B(n_33),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_346),
.Y(n_646)
);

BUFx12f_ASAP7_75t_L g647 ( 
.A(n_366),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_346),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_422),
.B(n_33),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_434),
.B(n_36),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_490),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_490),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_484),
.Y(n_653)
);

BUFx8_ASAP7_75t_L g654 ( 
.A(n_484),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_498),
.B(n_515),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_436),
.B(n_36),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_349),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_325),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_498),
.Y(n_659)
);

CKINVDCx11_ASAP7_75t_R g660 ( 
.A(n_499),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_515),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_439),
.B(n_443),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_456),
.B(n_37),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_330),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_481),
.B(n_37),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_532),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_495),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_532),
.Y(n_668)
);

INVx5_ASAP7_75t_L g669 ( 
.A(n_531),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_357),
.B(n_38),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_398),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_348),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_357),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_404),
.B(n_39),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_367),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_408),
.B(n_39),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_332),
.B(n_40),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_335),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_431),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_432),
.B(n_40),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_332),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_433),
.B(n_41),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_485),
.B(n_42),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_438),
.B(n_42),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_379),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_454),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_379),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_488),
.B(n_45),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_383),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_387),
.Y(n_690)
);

INVx5_ASAP7_75t_L g691 ( 
.A(n_383),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_393),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_492),
.B(n_45),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_493),
.B(n_46),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_473),
.B(n_46),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_469),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_508),
.B(n_47),
.Y(n_697)
);

NOR2x1_ASAP7_75t_L g698 ( 
.A(n_513),
.B(n_101),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_393),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_407),
.Y(n_700)
);

BUFx8_ASAP7_75t_SL g701 ( 
.A(n_372),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_407),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_474),
.B(n_482),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_496),
.B(n_47),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_483),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_523),
.Y(n_706)
);

BUFx8_ASAP7_75t_L g707 ( 
.A(n_470),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_518),
.B(n_48),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_522),
.B(n_48),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_561),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_590),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_670),
.A2(n_372),
.B1(n_428),
.B2(n_378),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_591),
.Y(n_713)
);

INVxp33_ASAP7_75t_L g714 ( 
.A(n_701),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_695),
.B(n_378),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_565),
.B(n_359),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_667),
.B(n_527),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_670),
.A2(n_444),
.B1(n_457),
.B2(n_428),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_L g719 ( 
.A1(n_657),
.A2(n_457),
.B1(n_472),
.B2(n_444),
.Y(n_719)
);

OA22x2_ASAP7_75t_L g720 ( 
.A1(n_558),
.A2(n_542),
.B1(n_491),
.B2(n_392),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_562),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_566),
.A2(n_478),
.B1(n_497),
.B2(n_472),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_704),
.A2(n_497),
.B1(n_506),
.B2(n_478),
.Y(n_723)
);

AND2x2_ASAP7_75t_SL g724 ( 
.A(n_575),
.B(n_480),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_587),
.A2(n_525),
.B1(n_506),
.B2(n_395),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_SL g726 ( 
.A1(n_569),
.A2(n_413),
.B1(n_423),
.B2(n_391),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_667),
.B(n_348),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_657),
.A2(n_525),
.B1(n_429),
.B2(n_437),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_SL g729 ( 
.A1(n_639),
.A2(n_442),
.B1(n_446),
.B2(n_427),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_591),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_667),
.B(n_448),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_564),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_SL g733 ( 
.A1(n_569),
.A2(n_465),
.B1(n_466),
.B2(n_463),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_SL g734 ( 
.A1(n_625),
.A2(n_487),
.B1(n_507),
.B2(n_486),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_669),
.B(n_510),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_588),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_673),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_636),
.Y(n_738)
);

OAI22xp33_ASAP7_75t_L g739 ( 
.A1(n_558),
.A2(n_519),
.B1(n_526),
.B2(n_512),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_658),
.B(n_529),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_578),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_557),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_SL g743 ( 
.A(n_594),
.B(n_528),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_581),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_622),
.B(n_537),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_596),
.A2(n_543),
.B1(n_541),
.B2(n_390),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_615),
.A2(n_629),
.B1(n_554),
.B2(n_589),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_669),
.B(n_350),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_602),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_669),
.B(n_350),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_585),
.A2(n_362),
.B1(n_354),
.B2(n_355),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_L g752 ( 
.A1(n_633),
.A2(n_516),
.B1(n_441),
.B2(n_451),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_590),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_590),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_633),
.B(n_351),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_608),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_658),
.B(n_533),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_SL g758 ( 
.A1(n_567),
.A2(n_538),
.B1(n_552),
.B2(n_534),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_573),
.B(n_351),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_675),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_622),
.B(n_49),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_557),
.B(n_451),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_557),
.B(n_548),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_608),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_633),
.A2(n_548),
.B1(n_550),
.B2(n_549),
.Y(n_765)
);

AND2x2_ASAP7_75t_SL g766 ( 
.A(n_645),
.B(n_416),
.Y(n_766)
);

AO22x2_ASAP7_75t_L g767 ( 
.A1(n_585),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_SL g768 ( 
.A1(n_611),
.A2(n_550),
.B1(n_549),
.B2(n_341),
.Y(n_768)
);

AND2x6_ASAP7_75t_L g769 ( 
.A(n_645),
.B(n_102),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_563),
.B(n_338),
.Y(n_770)
);

OAI22xp33_ASAP7_75t_L g771 ( 
.A1(n_623),
.A2(n_364),
.B1(n_368),
.B2(n_361),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_563),
.B(n_568),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_563),
.B(n_568),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_589),
.A2(n_623),
.B1(n_628),
.B2(n_583),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_608),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_628),
.A2(n_370),
.B1(n_375),
.B2(n_369),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_568),
.B(n_377),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_592),
.A2(n_385),
.B1(n_394),
.B2(n_384),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_620),
.A2(n_579),
.B1(n_631),
.B2(n_577),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_620),
.A2(n_401),
.B1(n_406),
.B2(n_397),
.Y(n_780)
);

OAI22xp33_ASAP7_75t_SL g781 ( 
.A1(n_662),
.A2(n_411),
.B1(n_414),
.B2(n_410),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_598),
.Y(n_782)
);

OAI22xp33_ASAP7_75t_SL g783 ( 
.A1(n_662),
.A2(n_418),
.B1(n_419),
.B2(n_415),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_577),
.B(n_421),
.Y(n_784)
);

NAND3x1_ASAP7_75t_L g785 ( 
.A(n_570),
.B(n_50),
.C(n_52),
.Y(n_785)
);

AND2x2_ASAP7_75t_SL g786 ( 
.A(n_592),
.B(n_606),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_606),
.A2(n_430),
.B1(n_435),
.B2(n_424),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_593),
.Y(n_788)
);

INVx5_ASAP7_75t_L g789 ( 
.A(n_577),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_603),
.Y(n_790)
);

INVx8_ASAP7_75t_L g791 ( 
.A(n_571),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_609),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_612),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_SL g794 ( 
.A1(n_570),
.A2(n_447),
.B1(n_449),
.B2(n_445),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_SL g795 ( 
.A1(n_572),
.A2(n_553),
.B1(n_546),
.B2(n_545),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_SL g796 ( 
.A1(n_555),
.A2(n_540),
.B1(n_536),
.B2(n_535),
.Y(n_796)
);

NOR2x1p5_ASAP7_75t_L g797 ( 
.A(n_635),
.B(n_450),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_632),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_632),
.Y(n_799)
);

OAI22xp33_ASAP7_75t_L g800 ( 
.A1(n_574),
.A2(n_530),
.B1(n_524),
.B2(n_520),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_655),
.B(n_452),
.Y(n_801)
);

AO22x2_ASAP7_75t_L g802 ( 
.A1(n_555),
.A2(n_703),
.B1(n_676),
.B2(n_680),
.Y(n_802)
);

AND2x2_ASAP7_75t_SL g803 ( 
.A(n_674),
.B(n_453),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_632),
.Y(n_804)
);

CKINVDCx6p67_ASAP7_75t_R g805 ( 
.A(n_613),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_626),
.B(n_455),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_630),
.Y(n_807)
);

OA22x2_ASAP7_75t_L g808 ( 
.A1(n_703),
.A2(n_517),
.B1(n_514),
.B2(n_511),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_559),
.B(n_52),
.Y(n_809)
);

OAI22xp33_ASAP7_75t_L g810 ( 
.A1(n_574),
.A2(n_505),
.B1(n_504),
.B2(n_503),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_661),
.B(n_459),
.Y(n_811)
);

AO22x2_ASAP7_75t_L g812 ( 
.A1(n_674),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_668),
.B(n_460),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_636),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_672),
.B(n_461),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_801),
.B(n_664),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_814),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_710),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_721),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_732),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_791),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_788),
.B(n_676),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_786),
.B(n_690),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_737),
.Y(n_824)
);

OR2x6_ASAP7_75t_L g825 ( 
.A(n_791),
.B(n_647),
.Y(n_825)
);

INVxp33_ASAP7_75t_SL g826 ( 
.A(n_795),
.Y(n_826)
);

INVxp33_ASAP7_75t_L g827 ( 
.A(n_760),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_SL g828 ( 
.A(n_766),
.B(n_654),
.Y(n_828)
);

XOR2xp5_ASAP7_75t_L g829 ( 
.A(n_712),
.B(n_634),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_759),
.B(n_601),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_782),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_740),
.B(n_664),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_757),
.B(n_678),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_790),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_712),
.Y(n_835)
);

XNOR2x2_ASAP7_75t_L g836 ( 
.A(n_718),
.B(n_660),
.Y(n_836)
);

XOR2xp5_ASAP7_75t_L g837 ( 
.A(n_718),
.B(n_698),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_792),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_805),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_793),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_778),
.B(n_678),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_713),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_807),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_730),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_741),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_778),
.B(n_654),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_744),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_749),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_729),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_753),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_738),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_787),
.B(n_610),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_787),
.B(n_617),
.Y(n_853)
);

XOR2x2_ASAP7_75t_L g854 ( 
.A(n_722),
.B(n_576),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_809),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_791),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_736),
.Y(n_857)
);

INVxp33_ASAP7_75t_L g858 ( 
.A(n_796),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_717),
.Y(n_859)
);

XOR2xp5_ASAP7_75t_L g860 ( 
.A(n_714),
.B(n_698),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_748),
.B(n_651),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_711),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_754),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_756),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_764),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_775),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_803),
.B(n_580),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_736),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_798),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_795),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_799),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_804),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_802),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_802),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_806),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_711),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_811),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_813),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_724),
.B(n_646),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_761),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_750),
.B(n_652),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_722),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_711),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_731),
.Y(n_884)
);

CKINVDCx14_ASAP7_75t_R g885 ( 
.A(n_715),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_735),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_815),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_762),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_763),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_773),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_770),
.B(n_784),
.Y(n_891)
);

XOR2xp5_ASAP7_75t_L g892 ( 
.A(n_723),
.B(n_601),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_794),
.B(n_580),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_780),
.B(n_666),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_747),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_742),
.B(n_646),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_747),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_751),
.B(n_646),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_796),
.B(n_680),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_745),
.B(n_605),
.Y(n_900)
);

CKINVDCx16_ASAP7_75t_R g901 ( 
.A(n_723),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_808),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_751),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_720),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_772),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_729),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_758),
.Y(n_907)
);

INVxp33_ASAP7_75t_L g908 ( 
.A(n_725),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_769),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_769),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_769),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_SL g912 ( 
.A(n_719),
.B(n_707),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_727),
.A2(n_586),
.B(n_582),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_725),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_824),
.Y(n_915)
);

AND2x6_ASAP7_75t_L g916 ( 
.A(n_909),
.B(n_769),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_830),
.B(n_746),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_832),
.B(n_746),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_827),
.B(n_716),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_818),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_900),
.B(n_767),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_821),
.B(n_789),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_819),
.Y(n_923)
);

BUFx8_ASAP7_75t_L g924 ( 
.A(n_899),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_827),
.B(n_716),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_823),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_895),
.B(n_897),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_840),
.B(n_767),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_840),
.B(n_812),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_820),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_845),
.Y(n_931)
);

NAND2x1p5_ASAP7_75t_L g932 ( 
.A(n_873),
.B(n_789),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_852),
.B(n_812),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_856),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_910),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_911),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_847),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_831),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_848),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_834),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_832),
.B(n_776),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_841),
.B(n_794),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_833),
.B(n_776),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_876),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_899),
.B(n_781),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_874),
.B(n_797),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_833),
.B(n_800),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_852),
.B(n_682),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_817),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_816),
.B(n_810),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_825),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_838),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_822),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_816),
.B(n_774),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_843),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_822),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_844),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_850),
.Y(n_958)
);

INVxp67_ASAP7_75t_SL g959 ( 
.A(n_891),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_880),
.B(n_605),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_908),
.B(n_682),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_907),
.B(n_684),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_828),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_861),
.B(n_707),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_901),
.B(n_728),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_887),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_841),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_861),
.B(n_771),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_846),
.B(n_684),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_846),
.B(n_640),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_853),
.B(n_679),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_853),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_851),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_825),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_913),
.A2(n_777),
.B(n_586),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_842),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_864),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_881),
.B(n_582),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_857),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_888),
.B(n_755),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_889),
.B(n_595),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_867),
.B(n_768),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_894),
.Y(n_983)
);

AND2x2_ASAP7_75t_SL g984 ( 
.A(n_912),
.B(n_595),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_855),
.B(n_679),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_825),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_867),
.B(n_894),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_868),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_884),
.B(n_686),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_892),
.B(n_739),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_859),
.B(n_886),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_903),
.B(n_696),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_879),
.B(n_614),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_893),
.A2(n_743),
.B1(n_600),
.B2(n_607),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_858),
.B(n_696),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_875),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_829),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_839),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_865),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_858),
.B(n_671),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_866),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_905),
.B(n_619),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_877),
.B(n_783),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_902),
.B(n_705),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_878),
.B(n_734),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_898),
.B(n_624),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_869),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_890),
.B(n_765),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_904),
.B(n_706),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_885),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_885),
.B(n_584),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_883),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_862),
.A2(n_627),
.B(n_624),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_849),
.B(n_584),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_854),
.B(n_649),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_871),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_872),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_862),
.A2(n_643),
.B(n_627),
.Y(n_1018)
);

BUFx2_ASAP7_75t_L g1019 ( 
.A(n_915),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_927),
.B(n_870),
.Y(n_1020)
);

BUFx12f_ASAP7_75t_L g1021 ( 
.A(n_915),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_919),
.Y(n_1022)
);

CKINVDCx14_ASAP7_75t_R g1023 ( 
.A(n_998),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_934),
.Y(n_1024)
);

AND2x6_ASAP7_75t_L g1025 ( 
.A(n_936),
.B(n_863),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_917),
.B(n_837),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_920),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_961),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_SL g1029 ( 
.A(n_942),
.B(n_826),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_936),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_936),
.Y(n_1031)
);

INVx5_ASAP7_75t_L g1032 ( 
.A(n_951),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_967),
.B(n_726),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_927),
.B(n_835),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_983),
.B(n_726),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_951),
.B(n_914),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_923),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_951),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_974),
.B(n_882),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_974),
.B(n_906),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_953),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_936),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_974),
.B(n_896),
.Y(n_1043)
);

INVx6_ASAP7_75t_L g1044 ( 
.A(n_986),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_972),
.B(n_860),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1015),
.B(n_970),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_930),
.Y(n_1047)
);

NAND2x1p5_ASAP7_75t_L g1048 ( 
.A(n_987),
.B(n_677),
.Y(n_1048)
);

OR2x6_ASAP7_75t_SL g1049 ( 
.A(n_990),
.B(n_836),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_SL g1050 ( 
.A(n_942),
.B(n_556),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_935),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_1000),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_986),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_941),
.B(n_779),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_986),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_971),
.Y(n_1056)
);

NOR2x1_ASAP7_75t_L g1057 ( 
.A(n_943),
.B(n_922),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_938),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_940),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_987),
.B(n_681),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_956),
.B(n_681),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_979),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_976),
.Y(n_1063)
);

BUFx8_ASAP7_75t_L g1064 ( 
.A(n_925),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_1012),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_954),
.B(n_733),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_918),
.B(n_752),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1015),
.B(n_636),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_971),
.B(n_681),
.Y(n_1069)
);

NOR2x1_ASAP7_75t_L g1070 ( 
.A(n_948),
.B(n_643),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_926),
.B(n_637),
.Y(n_1071)
);

NOR2x1_ASAP7_75t_L g1072 ( 
.A(n_948),
.B(n_969),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_976),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_924),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_1012),
.Y(n_1075)
);

CKINVDCx8_ASAP7_75t_R g1076 ( 
.A(n_946),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_959),
.B(n_685),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_952),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_947),
.B(n_685),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_935),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_1014),
.B(n_637),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_931),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_955),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_973),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1014),
.B(n_637),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_978),
.B(n_685),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_931),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_956),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_950),
.B(n_648),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_988),
.Y(n_1090)
);

BUFx12f_ASAP7_75t_L g1091 ( 
.A(n_924),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_926),
.B(n_638),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_995),
.B(n_638),
.Y(n_1093)
);

INVxp67_ASAP7_75t_SL g1094 ( 
.A(n_928),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_937),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_935),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1006),
.B(n_687),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_939),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_995),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_973),
.Y(n_1100)
);

OR2x6_ASAP7_75t_L g1101 ( 
.A(n_1010),
.B(n_785),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_993),
.B(n_687),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_965),
.B(n_650),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_939),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1027),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1031),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1037),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1031),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_1041),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_1091),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1047),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_1031),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_1032),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_1021),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1063),
.Y(n_1115)
);

CKINVDCx16_ASAP7_75t_R g1116 ( 
.A(n_1062),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1090),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_1032),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_1094),
.Y(n_1119)
);

INVx5_ASAP7_75t_L g1120 ( 
.A(n_1025),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1084),
.Y(n_1121)
);

INVx5_ASAP7_75t_L g1122 ( 
.A(n_1025),
.Y(n_1122)
);

INVxp67_ASAP7_75t_SL g1123 ( 
.A(n_1094),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1073),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1020),
.B(n_929),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_1038),
.B(n_973),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1044),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1024),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1058),
.Y(n_1129)
);

BUFx5_ASAP7_75t_L g1130 ( 
.A(n_1025),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1084),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_1044),
.Y(n_1132)
);

INVx6_ASAP7_75t_L g1133 ( 
.A(n_1038),
.Y(n_1133)
);

CKINVDCx6p67_ASAP7_75t_R g1134 ( 
.A(n_1019),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1067),
.B(n_933),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_1020),
.Y(n_1136)
);

INVx3_ASAP7_75t_SL g1137 ( 
.A(n_1101),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_1053),
.Y(n_1138)
);

INVx8_ASAP7_75t_L g1139 ( 
.A(n_1025),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_1042),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1042),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1059),
.Y(n_1142)
);

INVx6_ASAP7_75t_L g1143 ( 
.A(n_1065),
.Y(n_1143)
);

BUFx4_ASAP7_75t_SL g1144 ( 
.A(n_1074),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1078),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1029),
.B(n_1054),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1083),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1087),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1082),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1046),
.B(n_933),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_1055),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1100),
.B(n_1042),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1100),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1030),
.Y(n_1154)
);

CKINVDCx8_ASAP7_75t_R g1155 ( 
.A(n_1040),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1104),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_1068),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1095),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1099),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1098),
.Y(n_1160)
);

INVx5_ASAP7_75t_SL g1161 ( 
.A(n_1065),
.Y(n_1161)
);

BUFx2_ASAP7_75t_SL g1162 ( 
.A(n_1076),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1081),
.B(n_928),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_1065),
.Y(n_1164)
);

INVx5_ASAP7_75t_L g1165 ( 
.A(n_1075),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_1075),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1075),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1030),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1051),
.Y(n_1169)
);

OR2x2_ASAP7_75t_L g1170 ( 
.A(n_1103),
.B(n_997),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1051),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1080),
.Y(n_1172)
);

NAND2x1p5_ASAP7_75t_L g1173 ( 
.A(n_1080),
.B(n_1017),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1105),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1146),
.B(n_1034),
.Y(n_1175)
);

BUFx4f_ASAP7_75t_SL g1176 ( 
.A(n_1134),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1144),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1146),
.B(n_1034),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1135),
.B(n_1026),
.Y(n_1179)
);

BUFx12f_ASAP7_75t_L g1180 ( 
.A(n_1114),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1136),
.A2(n_1029),
.B1(n_1045),
.B2(n_984),
.Y(n_1181)
);

CKINVDCx6p67_ASAP7_75t_R g1182 ( 
.A(n_1116),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1107),
.Y(n_1183)
);

CKINVDCx11_ASAP7_75t_R g1184 ( 
.A(n_1134),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_SL g1185 ( 
.A1(n_1125),
.A2(n_984),
.B1(n_1066),
.B2(n_929),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1170),
.A2(n_1072),
.B1(n_1011),
.B2(n_1040),
.Y(n_1186)
);

OAI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1150),
.A2(n_1033),
.B1(n_1028),
.B2(n_968),
.Y(n_1187)
);

BUFx8_ASAP7_75t_L g1188 ( 
.A(n_1128),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1125),
.A2(n_1011),
.B1(n_1039),
.B2(n_1036),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1123),
.A2(n_1056),
.B1(n_1028),
.B2(n_994),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1125),
.A2(n_1039),
.B1(n_1036),
.B2(n_1052),
.Y(n_1191)
);

INVx6_ASAP7_75t_L g1192 ( 
.A(n_1110),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1149),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1119),
.A2(n_1052),
.B1(n_946),
.B2(n_924),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1111),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1149),
.Y(n_1196)
);

CKINVDCx11_ASAP7_75t_R g1197 ( 
.A(n_1110),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_SL g1198 ( 
.A1(n_1119),
.A2(n_982),
.B1(n_1033),
.B2(n_1050),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1158),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1157),
.A2(n_982),
.B1(n_1056),
.B2(n_1035),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1117),
.Y(n_1201)
);

INVx1_ASAP7_75t_SL g1202 ( 
.A(n_1109),
.Y(n_1202)
);

INVx4_ASAP7_75t_SL g1203 ( 
.A(n_1137),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1158),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1160),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1163),
.A2(n_946),
.B1(n_945),
.B2(n_966),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_L g1207 ( 
.A(n_1137),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1129),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1109),
.A2(n_1070),
.B1(n_1035),
.B2(n_996),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1139),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1171),
.A2(n_1057),
.B(n_1002),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1142),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_1143),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1138),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_1161),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1159),
.B(n_1085),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1162),
.A2(n_1050),
.B1(n_921),
.B2(n_1049),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1145),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1138),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1127),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1147),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1169),
.A2(n_996),
.B1(n_966),
.B2(n_1048),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1148),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1127),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1132),
.Y(n_1225)
);

INVx8_ASAP7_75t_L g1226 ( 
.A(n_1139),
.Y(n_1226)
);

INVx6_ASAP7_75t_L g1227 ( 
.A(n_1165),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1160),
.A2(n_945),
.B1(n_1093),
.B2(n_1005),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1155),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1143),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1132),
.Y(n_1231)
);

INVx8_ASAP7_75t_L g1232 ( 
.A(n_1139),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1171),
.A2(n_1008),
.B(n_1013),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1169),
.A2(n_981),
.B1(n_1096),
.B2(n_1018),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1156),
.A2(n_1093),
.B1(n_921),
.B2(n_1008),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1115),
.A2(n_1005),
.B1(n_1022),
.B2(n_1003),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_1139),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_SL g1238 ( 
.A1(n_1120),
.A2(n_964),
.B1(n_963),
.B2(n_1023),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1120),
.A2(n_1064),
.B1(n_1092),
.B2(n_1071),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1216),
.B(n_1071),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1226),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1175),
.B(n_1092),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1179),
.A2(n_1003),
.B1(n_618),
.B2(n_621),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1200),
.A2(n_1120),
.B1(n_1122),
.B2(n_1130),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1185),
.A2(n_644),
.B1(n_604),
.B2(n_649),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1187),
.A2(n_1217),
.B1(n_1178),
.B2(n_1181),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1198),
.A2(n_1173),
.B1(n_1169),
.B2(n_1096),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1202),
.A2(n_1173),
.B1(n_1172),
.B2(n_991),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1186),
.A2(n_989),
.B1(n_1089),
.B2(n_1124),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1174),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1226),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1202),
.A2(n_1172),
.B1(n_1133),
.B2(n_1120),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1189),
.A2(n_989),
.B1(n_1089),
.B2(n_1124),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1183),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1193),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1235),
.A2(n_1060),
.B1(n_650),
.B2(n_663),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1190),
.A2(n_1200),
.B1(n_1209),
.B2(n_1235),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1201),
.A2(n_1176),
.B1(n_1222),
.B2(n_1206),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1215),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1191),
.A2(n_1194),
.B1(n_1228),
.B2(n_1236),
.Y(n_1260)
);

NAND2x1_ASAP7_75t_L g1261 ( 
.A(n_1210),
.B(n_1237),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1195),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1238),
.A2(n_989),
.B1(n_1017),
.B2(n_1064),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1239),
.A2(n_992),
.B1(n_980),
.B2(n_977),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1229),
.A2(n_992),
.B1(n_980),
.B2(n_999),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1197),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1196),
.A2(n_980),
.B1(n_1007),
.B2(n_1001),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1201),
.A2(n_1088),
.B1(n_962),
.B2(n_709),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_SL g1269 ( 
.A1(n_1177),
.A2(n_665),
.B(n_656),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1199),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1220),
.B(n_1161),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1204),
.A2(n_1016),
.B1(n_957),
.B2(n_958),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1182),
.B(n_1167),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1208),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1212),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1234),
.A2(n_1133),
.B1(n_1122),
.B2(n_1154),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1218),
.B(n_1221),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1223),
.A2(n_1069),
.B1(n_962),
.B2(n_688),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1233),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1220),
.B(n_960),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1211),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1205),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1210),
.A2(n_688),
.B(n_683),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1207),
.A2(n_1133),
.B1(n_1122),
.B2(n_1154),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1192),
.A2(n_1154),
.B1(n_693),
.B2(n_694),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1214),
.A2(n_693),
.B1(n_694),
.B2(n_683),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1224),
.B(n_985),
.Y(n_1287)
);

NOR2x1_ASAP7_75t_SL g1288 ( 
.A(n_1237),
.B(n_1113),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1230),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1219),
.A2(n_708),
.B1(n_697),
.B2(n_1077),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1230),
.Y(n_1291)
);

INVx8_ASAP7_75t_L g1292 ( 
.A(n_1226),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1192),
.A2(n_1086),
.B1(n_1126),
.B2(n_1102),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1232),
.Y(n_1294)
);

INVx1_ASAP7_75t_SL g1295 ( 
.A(n_1224),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1225),
.A2(n_1086),
.B1(n_1126),
.B2(n_1102),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1232),
.A2(n_1130),
.B1(n_1151),
.B2(n_1079),
.Y(n_1297)
);

BUFx4f_ASAP7_75t_SL g1298 ( 
.A(n_1180),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1257),
.A2(n_641),
.B1(n_642),
.B2(n_638),
.Y(n_1299)
);

AOI222xp33_ASAP7_75t_L g1300 ( 
.A1(n_1246),
.A2(n_1203),
.B1(n_985),
.B2(n_1004),
.C1(n_1009),
.C2(n_1188),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1255),
.Y(n_1301)
);

OAI222xp33_ASAP7_75t_L g1302 ( 
.A1(n_1260),
.A2(n_1079),
.B1(n_1097),
.B2(n_1061),
.C1(n_1164),
.C2(n_1166),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1260),
.A2(n_659),
.B1(n_958),
.B2(n_949),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1249),
.A2(n_958),
.B1(n_949),
.B2(n_1097),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1245),
.A2(n_1253),
.B1(n_1242),
.B2(n_1265),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1264),
.A2(n_949),
.B1(n_699),
.B2(n_700),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1277),
.B(n_1250),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1240),
.A2(n_1243),
.B1(n_1256),
.B2(n_1280),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1254),
.B(n_1225),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1243),
.A2(n_699),
.B1(n_700),
.B2(n_689),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1286),
.B(n_975),
.C(n_1188),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1279),
.B(n_56),
.Y(n_1312)
);

OAI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1286),
.A2(n_1278),
.B1(n_1290),
.B2(n_1268),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1259),
.B(n_1225),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1278),
.A2(n_1165),
.B1(n_1166),
.B2(n_1164),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1279),
.B(n_58),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1290),
.A2(n_1164),
.B1(n_1108),
.B2(n_1112),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1287),
.A2(n_699),
.B1(n_700),
.B2(n_689),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1244),
.A2(n_702),
.B1(n_689),
.B2(n_1043),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1262),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1282),
.A2(n_702),
.B1(n_1043),
.B2(n_1231),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1263),
.A2(n_702),
.B1(n_1231),
.B2(n_944),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1267),
.A2(n_1231),
.B1(n_944),
.B2(n_1004),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1270),
.A2(n_1248),
.B1(n_1258),
.B2(n_1281),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1269),
.B(n_653),
.C(n_648),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1283),
.A2(n_1285),
.B1(n_1247),
.B2(n_1273),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1281),
.A2(n_944),
.B1(n_1004),
.B2(n_1009),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1274),
.A2(n_1203),
.B1(n_1184),
.B2(n_1232),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1272),
.A2(n_1009),
.B1(n_1130),
.B2(n_560),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1275),
.A2(n_1130),
.B1(n_560),
.B2(n_556),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1289),
.A2(n_1168),
.B1(n_916),
.B2(n_691),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_SL g1332 ( 
.A(n_1266),
.B(n_467),
.C(n_464),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1276),
.A2(n_1140),
.B1(n_1108),
.B2(n_1112),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1241),
.A2(n_1140),
.B1(n_1106),
.B2(n_1141),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1291),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1295),
.B(n_1106),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1252),
.A2(n_1293),
.B1(n_1296),
.B2(n_1297),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1241),
.A2(n_1141),
.B1(n_1168),
.B2(n_1227),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1284),
.A2(n_1168),
.B1(n_916),
.B2(n_691),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1271),
.A2(n_1168),
.B1(n_916),
.B2(n_692),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1292),
.Y(n_1341)
);

OAI222xp33_ASAP7_75t_L g1342 ( 
.A1(n_1298),
.A2(n_1118),
.B1(n_1113),
.B2(n_1152),
.C1(n_932),
.C2(n_475),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1251),
.A2(n_1121),
.B1(n_1153),
.B2(n_1131),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1294),
.B(n_1121),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1292),
.A2(n_1153),
.B1(n_1131),
.B2(n_1118),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1261),
.A2(n_1153),
.B1(n_1131),
.B2(n_1118),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1288),
.A2(n_1153),
.B1(n_1131),
.B2(n_1113),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1245),
.A2(n_477),
.B1(n_501),
.B2(n_500),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1277),
.B(n_1213),
.Y(n_1349)
);

OAI21xp33_ASAP7_75t_L g1350 ( 
.A1(n_1245),
.A2(n_489),
.B(n_471),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1307),
.B(n_59),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1313),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_1352)
);

OAI221xp5_ASAP7_75t_L g1353 ( 
.A1(n_1350),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.C(n_68),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1326),
.B(n_616),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1320),
.B(n_1335),
.Y(n_1355)
);

NAND4xp25_ASAP7_75t_L g1356 ( 
.A(n_1325),
.B(n_69),
.C(n_70),
.D(n_71),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1311),
.A2(n_71),
.B(n_72),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1350),
.A2(n_616),
.B1(n_599),
.B2(n_597),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1311),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1337),
.A2(n_73),
.B(n_74),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1312),
.B(n_75),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1333),
.A2(n_76),
.B(n_77),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1314),
.B(n_76),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1316),
.B(n_79),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1308),
.B(n_80),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1309),
.B(n_81),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1324),
.B(n_82),
.Y(n_1367)
);

OAI221xp5_ASAP7_75t_L g1368 ( 
.A1(n_1305),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.C(n_87),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1349),
.B(n_83),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1328),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1336),
.B(n_105),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1328),
.B(n_324),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1344),
.B(n_108),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1341),
.B(n_315),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1301),
.B(n_313),
.Y(n_1375)
);

OAI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1300),
.A2(n_112),
.B1(n_118),
.B2(n_122),
.C(n_124),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1301),
.Y(n_1377)
);

NAND2x1p5_ASAP7_75t_L g1378 ( 
.A(n_1341),
.B(n_126),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1317),
.B(n_308),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1299),
.B(n_127),
.Y(n_1380)
);

NAND3xp33_ASAP7_75t_L g1381 ( 
.A(n_1348),
.B(n_131),
.C(n_132),
.Y(n_1381)
);

AOI211xp5_ASAP7_75t_L g1382 ( 
.A1(n_1332),
.A2(n_135),
.B(n_143),
.C(n_146),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1347),
.B(n_1343),
.Y(n_1383)
);

AOI221xp5_ASAP7_75t_L g1384 ( 
.A1(n_1310),
.A2(n_1302),
.B1(n_1342),
.B2(n_1327),
.C(n_1303),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1315),
.A2(n_147),
.B1(n_157),
.B2(n_158),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1355),
.B(n_1345),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1354),
.B(n_1334),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1357),
.B(n_1346),
.C(n_1318),
.Y(n_1388)
);

OA211x2_ASAP7_75t_L g1389 ( 
.A1(n_1354),
.A2(n_1319),
.B(n_1339),
.C(n_1331),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1355),
.B(n_1338),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1366),
.Y(n_1391)
);

NAND3xp33_ASAP7_75t_L g1392 ( 
.A(n_1360),
.B(n_1304),
.C(n_1321),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1360),
.B(n_1329),
.C(n_1340),
.Y(n_1393)
);

NAND4xp25_ASAP7_75t_L g1394 ( 
.A(n_1352),
.B(n_1356),
.C(n_1359),
.D(n_1370),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1363),
.B(n_1322),
.Y(n_1395)
);

NOR3xp33_ASAP7_75t_L g1396 ( 
.A(n_1353),
.B(n_1306),
.C(n_1323),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1351),
.B(n_160),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1352),
.B(n_1330),
.C(n_163),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1364),
.B(n_167),
.Y(n_1399)
);

OAI211xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1361),
.A2(n_173),
.B(n_175),
.C(n_176),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1383),
.B(n_182),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1377),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1365),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1369),
.B(n_187),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1362),
.A2(n_189),
.B(n_190),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1365),
.A2(n_193),
.B1(n_197),
.B2(n_204),
.Y(n_1406)
);

AO21x2_ASAP7_75t_L g1407 ( 
.A1(n_1375),
.A2(n_207),
.B(n_209),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1367),
.B(n_210),
.Y(n_1408)
);

NAND4xp75_ASAP7_75t_L g1409 ( 
.A(n_1405),
.B(n_1372),
.C(n_1384),
.D(n_1383),
.Y(n_1409)
);

NAND4xp75_ASAP7_75t_L g1410 ( 
.A(n_1389),
.B(n_1379),
.C(n_1358),
.D(n_1374),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1402),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1390),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1386),
.Y(n_1413)
);

NAND4xp75_ASAP7_75t_L g1414 ( 
.A(n_1401),
.B(n_1380),
.C(n_1373),
.D(n_1371),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1391),
.B(n_1378),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1408),
.Y(n_1416)
);

XNOR2xp5_ASAP7_75t_L g1417 ( 
.A(n_1404),
.B(n_1399),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1395),
.Y(n_1418)
);

XNOR2xp5_ASAP7_75t_L g1419 ( 
.A(n_1394),
.B(n_1368),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1387),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1407),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1403),
.A2(n_1376),
.B1(n_1382),
.B2(n_1381),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1407),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1397),
.B(n_1388),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1411),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_1417),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1411),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1418),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1413),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1420),
.B(n_1385),
.Y(n_1430)
);

XNOR2x2_ASAP7_75t_L g1431 ( 
.A(n_1409),
.B(n_1393),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1412),
.B(n_1406),
.Y(n_1432)
);

XOR2x2_ASAP7_75t_L g1433 ( 
.A(n_1419),
.B(n_1396),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1416),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1424),
.B(n_1400),
.Y(n_1435)
);

CKINVDCx16_ASAP7_75t_R g1436 ( 
.A(n_1415),
.Y(n_1436)
);

XOR2x2_ASAP7_75t_L g1437 ( 
.A(n_1410),
.B(n_1414),
.Y(n_1437)
);

INVxp67_ASAP7_75t_SL g1438 ( 
.A(n_1435),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1425),
.Y(n_1439)
);

OA22x2_ASAP7_75t_L g1440 ( 
.A1(n_1426),
.A2(n_1430),
.B1(n_1431),
.B2(n_1432),
.Y(n_1440)
);

XOR2x2_ASAP7_75t_SL g1441 ( 
.A(n_1437),
.B(n_1422),
.Y(n_1441)
);

XNOR2xp5_ASAP7_75t_L g1442 ( 
.A(n_1433),
.B(n_1414),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1427),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1434),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_SL g1445 ( 
.A1(n_1436),
.A2(n_1423),
.B1(n_1421),
.B2(n_1398),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1428),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1429),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1439),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1443),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1443),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1446),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1440),
.Y(n_1452)
);

XOR2xp5_ASAP7_75t_L g1453 ( 
.A(n_1442),
.B(n_1392),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1444),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1438),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_L g1456 ( 
.A1(n_1452),
.A2(n_1445),
.B1(n_1441),
.B2(n_1444),
.C(n_1447),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1455),
.Y(n_1457)
);

AND4x1_ASAP7_75t_L g1458 ( 
.A(n_1451),
.B(n_1454),
.C(n_1450),
.D(n_1448),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1449),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_SL g1460 ( 
.A1(n_1456),
.A2(n_1449),
.B(n_1453),
.C(n_1400),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1457),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1459),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1458),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1461),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1460),
.A2(n_211),
.B(n_216),
.C(n_220),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1463),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1462),
.B(n_221),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1461),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1464),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1467),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1468),
.Y(n_1471)
);

NOR3xp33_ASAP7_75t_L g1472 ( 
.A(n_1465),
.B(n_225),
.C(n_228),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1466),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1473),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1469),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1471),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1470),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1472),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1474),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1475),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1476),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1478),
.Y(n_1482)
);

AO22x2_ASAP7_75t_L g1483 ( 
.A1(n_1479),
.A2(n_1477),
.B1(n_242),
.B2(n_243),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1482),
.A2(n_239),
.B1(n_245),
.B2(n_250),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1480),
.Y(n_1485)
);

INVxp67_ASAP7_75t_SL g1486 ( 
.A(n_1485),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1483),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1487),
.A2(n_1481),
.B1(n_1484),
.B2(n_258),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1486),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1489),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1488),
.Y(n_1491)
);

AO22x2_ASAP7_75t_L g1492 ( 
.A1(n_1490),
.A2(n_271),
.B1(n_279),
.B2(n_280),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1491),
.A2(n_281),
.B1(n_284),
.B2(n_289),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1492),
.Y(n_1494)
);

AOI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1494),
.A2(n_1493),
.B1(n_290),
.B2(n_291),
.C(n_292),
.Y(n_1495)
);

AOI211xp5_ASAP7_75t_L g1496 ( 
.A1(n_1495),
.A2(n_296),
.B(n_297),
.C(n_299),
.Y(n_1496)
);


endmodule