module fake_ariane_1110_n_29 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_29);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_29;

wire n_24;
wire n_22;
wire n_13;
wire n_20;
wire n_27;
wire n_17;
wire n_18;
wire n_28;
wire n_11;
wire n_26;
wire n_14;
wire n_19;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_10;
wire n_25;

INVx4_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_9),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

AND2x6_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_3),
.Y(n_13)
);

AND2x6_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_7),
.Y(n_15)
);

OAI22xp33_ASAP7_75t_L g16 ( 
.A1(n_10),
.A2(n_0),
.B1(n_2),
.B2(n_6),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_8),
.B(n_0),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NAND2x1p5_ASAP7_75t_SL g20 ( 
.A(n_18),
.B(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_23),
.A2(n_17),
.B(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_20),
.B(n_26),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_20),
.B1(n_26),
.B2(n_28),
.Y(n_29)
);


endmodule