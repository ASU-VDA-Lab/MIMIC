module fake_jpeg_596_n_111 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_38),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_36),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_31),
.B1(n_30),
.B2(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_51),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_32),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_29),
.B1(n_39),
.B2(n_32),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_41),
.C(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_60),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_1),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_51),
.B1(n_47),
.B2(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_5),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_47),
.B1(n_48),
.B2(n_44),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_44),
.B1(n_39),
.B2(n_14),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_15),
.B(n_26),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_77),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_1),
.B(n_2),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_80),
.B(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_2),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_17),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_3),
.B(n_4),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_3),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_16),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_71),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_92),
.B(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_6),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_21),
.C(n_24),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_81),
.B(n_22),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_23),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_93),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_96),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_94),
.B(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_97),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_SL g107 ( 
.A(n_106),
.B(n_87),
.C(n_9),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_81),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_28),
.Y(n_111)
);


endmodule