module real_aes_16280_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_1983, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_1983;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1694;
wire n_1224;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_1940;
wire n_715;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_1648;
wire n_724;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_1951;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_1689;
wire n_998;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1908;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1899;
wire n_816;
wire n_1470;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1638;
wire n_1072;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1939;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1671;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1855;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_1969;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
AOI221xp5_ASAP7_75t_L g1652 ( .A1(n_0), .A2(n_102), .B1(n_577), .B2(n_695), .C(n_1019), .Y(n_1652) );
AOI22xp33_ASAP7_75t_SL g1665 ( .A1(n_0), .A2(n_243), .B1(n_1122), .B2(n_1666), .Y(n_1665) );
OAI22xp5_ASAP7_75t_L g1423 ( .A1(n_1), .A2(n_105), .B1(n_531), .B2(n_540), .Y(n_1423) );
OAI22xp33_ASAP7_75t_L g1454 ( .A1(n_1), .A2(n_187), .B1(n_488), .B2(n_491), .Y(n_1454) );
INVx1_ASAP7_75t_L g389 ( .A(n_2), .Y(n_389) );
AND2x2_ASAP7_75t_L g418 ( .A(n_2), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g534 ( .A(n_2), .B(n_260), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_2), .B(n_399), .Y(n_560) );
INVx1_ASAP7_75t_L g1011 ( .A(n_3), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_3), .A2(n_72), .B1(n_440), .B2(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1564 ( .A(n_4), .Y(n_1564) );
AOI22xp5_ASAP7_75t_L g1585 ( .A1(n_4), .A2(n_11), .B1(n_694), .B2(n_1141), .Y(n_1585) );
AOI22xp33_ASAP7_75t_SL g1901 ( .A1(n_5), .A2(n_39), .B1(n_480), .B2(n_722), .Y(n_1901) );
INVxp67_ASAP7_75t_SL g1922 ( .A(n_5), .Y(n_1922) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_6), .A2(n_282), .B1(n_1205), .B2(n_1208), .Y(n_1204) );
OAI22xp33_ASAP7_75t_L g1236 ( .A1(n_6), .A2(n_282), .B1(n_1237), .B2(n_1240), .Y(n_1236) );
INVx1_ASAP7_75t_L g1601 ( .A(n_7), .Y(n_1601) );
OAI221xp5_ASAP7_75t_L g1625 ( .A1(n_7), .A2(n_144), .B1(n_677), .B2(n_1626), .C(n_1627), .Y(n_1625) );
INVx1_ASAP7_75t_L g1646 ( .A(n_8), .Y(n_1646) );
OAI22xp33_ASAP7_75t_L g1670 ( .A1(n_8), .A2(n_85), .B1(n_1613), .B2(n_1671), .Y(n_1670) );
INVx1_ASAP7_75t_L g999 ( .A(n_9), .Y(n_999) );
INVx1_ASAP7_75t_L g728 ( .A(n_10), .Y(n_728) );
OA222x2_ASAP7_75t_L g750 ( .A1(n_10), .A2(n_146), .B1(n_174), .B2(n_751), .C1(n_753), .C2(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g1573 ( .A(n_11), .Y(n_1573) );
OAI221xp5_ASAP7_75t_L g1050 ( .A1(n_12), .A2(n_363), .B1(n_440), .B2(n_445), .C(n_451), .Y(n_1050) );
OAI21xp33_ASAP7_75t_SL g1078 ( .A1(n_12), .A2(n_596), .B(n_754), .Y(n_1078) );
INVx1_ASAP7_75t_L g1197 ( .A(n_13), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1522 ( .A1(n_14), .A2(n_60), .B1(n_713), .B2(n_935), .Y(n_1522) );
AOI221xp5_ASAP7_75t_L g1537 ( .A1(n_14), .A2(n_332), .B1(n_1018), .B2(n_1141), .C(n_1142), .Y(n_1537) );
AOI221xp5_ASAP7_75t_L g1638 ( .A1(n_15), .A2(n_84), .B1(n_577), .B2(n_1639), .C(n_1641), .Y(n_1638) );
AOI22xp33_ASAP7_75t_SL g1669 ( .A1(n_15), .A2(n_204), .B1(n_480), .B2(n_639), .Y(n_1669) );
INVx2_ASAP7_75t_L g435 ( .A(n_16), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g1720 ( .A1(n_17), .A2(n_20), .B1(n_1684), .B2(n_1692), .Y(n_1720) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_18), .A2(n_176), .B1(n_710), .B2(n_719), .Y(n_718) );
INVxp67_ASAP7_75t_SL g777 ( .A(n_18), .Y(n_777) );
INVx1_ASAP7_75t_L g1158 ( .A(n_19), .Y(n_1158) );
OAI22xp33_ASAP7_75t_L g1061 ( .A1(n_21), .A2(n_306), .B1(n_488), .B2(n_491), .Y(n_1061) );
INVx1_ASAP7_75t_L g1077 ( .A(n_21), .Y(n_1077) );
INVx1_ASAP7_75t_L g1467 ( .A(n_22), .Y(n_1467) );
OAI211xp5_ASAP7_75t_L g1191 ( .A1(n_23), .A2(n_1192), .B(n_1193), .C(n_1196), .Y(n_1191) );
INVx1_ASAP7_75t_L g1235 ( .A(n_23), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_24), .A2(n_362), .B1(n_620), .B2(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_24), .A2(n_160), .B1(n_580), .B2(n_581), .Y(n_668) );
CKINVDCx5p33_ASAP7_75t_R g1510 ( .A(n_25), .Y(n_1510) );
XOR2x1_ASAP7_75t_L g409 ( .A(n_26), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g969 ( .A(n_27), .Y(n_969) );
AOI221x1_ASAP7_75t_SL g974 ( .A1(n_27), .A2(n_202), .B1(n_526), .B2(n_886), .C(n_975), .Y(n_974) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_28), .Y(n_384) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_28), .B(n_382), .Y(n_1685) );
INVx1_ASAP7_75t_L g1168 ( .A(n_29), .Y(n_1168) );
OA22x2_ASAP7_75t_L g1300 ( .A1(n_30), .A2(n_1301), .B1(n_1367), .B2(n_1368), .Y(n_1300) );
INVxp67_ASAP7_75t_L g1368 ( .A(n_30), .Y(n_1368) );
AOI22xp33_ASAP7_75t_L g1765 ( .A1(n_31), .A2(n_192), .B1(n_1692), .B2(n_1716), .Y(n_1765) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_32), .A2(n_234), .B1(n_629), .B2(n_723), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_32), .A2(n_314), .B1(n_780), .B2(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g963 ( .A(n_33), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_33), .A2(n_178), .B1(n_548), .B2(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g1323 ( .A(n_34), .Y(n_1323) );
OAI211xp5_ASAP7_75t_SL g1463 ( .A1(n_35), .A2(n_1464), .B(n_1466), .C(n_1469), .Y(n_1463) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_35), .A2(n_291), .B1(n_650), .B2(n_1502), .Y(n_1501) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_36), .A2(n_269), .B1(n_457), .B2(n_464), .Y(n_456) );
INVxp33_ASAP7_75t_L g594 ( .A(n_36), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_37), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_37), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_38), .Y(n_959) );
AOI221xp5_ASAP7_75t_L g1915 ( .A1(n_39), .A2(n_88), .B1(n_563), .B2(n_1088), .C(n_1641), .Y(n_1915) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_40), .A2(n_288), .B1(n_707), .B2(n_710), .Y(n_706) );
INVxp67_ASAP7_75t_SL g764 ( .A(n_40), .Y(n_764) );
INVx1_ASAP7_75t_L g1386 ( .A(n_41), .Y(n_1386) );
INVx1_ASAP7_75t_L g1383 ( .A(n_42), .Y(n_1383) );
AOI221xp5_ASAP7_75t_L g1405 ( .A1(n_42), .A2(n_279), .B1(n_576), .B2(n_578), .C(n_1406), .Y(n_1405) );
OAI221xp5_ASAP7_75t_L g1472 ( .A1(n_43), .A2(n_111), .B1(n_681), .B2(n_1473), .C(n_1474), .Y(n_1472) );
OAI22xp33_ASAP7_75t_L g1494 ( .A1(n_43), .A2(n_111), .B1(n_1495), .B2(n_1497), .Y(n_1494) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_44), .A2(n_195), .B1(n_526), .B2(n_779), .Y(n_890) );
INVx1_ASAP7_75t_L g925 ( .A(n_44), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g1428 ( .A1(n_45), .A2(n_57), .B1(n_583), .B2(n_1429), .C(n_1430), .Y(n_1428) );
AOI221xp5_ASAP7_75t_L g1451 ( .A1(n_45), .A2(n_134), .B1(n_480), .B2(n_710), .C(n_1452), .Y(n_1451) );
AOI22xp33_ASAP7_75t_SL g1478 ( .A1(n_46), .A2(n_264), .B1(n_1479), .B2(n_1480), .Y(n_1478) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_46), .A2(n_366), .B1(n_480), .B2(n_640), .Y(n_1489) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_47), .A2(n_123), .B1(n_615), .B2(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_SL g691 ( .A(n_47), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g1714 ( .A1(n_48), .A2(n_211), .B1(n_1684), .B2(n_1689), .Y(n_1714) );
AOI22xp5_ASAP7_75t_L g1700 ( .A1(n_49), .A2(n_351), .B1(n_1692), .B2(n_1701), .Y(n_1700) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_50), .Y(n_396) );
INVx1_ASAP7_75t_L g1563 ( .A(n_51), .Y(n_1563) );
AOI22xp33_ASAP7_75t_L g1587 ( .A1(n_51), .A2(n_188), .B1(n_576), .B2(n_694), .Y(n_1587) );
AOI22xp5_ASAP7_75t_L g1715 ( .A1(n_52), .A2(n_330), .B1(n_1692), .B2(n_1716), .Y(n_1715) );
AOI22xp5_ASAP7_75t_L g1724 ( .A1(n_53), .A2(n_127), .B1(n_1684), .B2(n_1689), .Y(n_1724) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_54), .A2(n_225), .B1(n_840), .B2(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g919 ( .A(n_54), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1902 ( .A1(n_55), .A2(n_274), .B1(n_935), .B2(n_1903), .Y(n_1902) );
AOI22xp33_ASAP7_75t_L g1916 ( .A1(n_55), .A2(n_141), .B1(n_581), .B2(n_1135), .Y(n_1916) );
OAI222xp33_ASAP7_75t_L g1251 ( .A1(n_56), .A2(n_73), .B1(n_1252), .B2(n_1253), .C1(n_1261), .C2(n_1269), .Y(n_1251) );
INVx1_ASAP7_75t_L g1284 ( .A(n_56), .Y(n_1284) );
INVx1_ASAP7_75t_L g1448 ( .A(n_57), .Y(n_1448) );
AOI22xp33_ASAP7_75t_SL g1121 ( .A1(n_58), .A2(n_169), .B1(n_1112), .B2(n_1122), .Y(n_1121) );
AOI221xp5_ASAP7_75t_L g1140 ( .A1(n_58), .A2(n_121), .B1(n_665), .B2(n_1141), .C(n_1142), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1387 ( .A1(n_59), .A2(n_303), .B1(n_457), .B2(n_464), .Y(n_1387) );
INVxp67_ASAP7_75t_SL g1390 ( .A(n_59), .Y(n_1390) );
AOI22xp33_ASAP7_75t_SL g1535 ( .A1(n_60), .A2(n_145), .B1(n_580), .B2(n_581), .Y(n_1535) );
INVx1_ASAP7_75t_L g1126 ( .A(n_61), .Y(n_1126) );
AOI21xp33_ASAP7_75t_L g1062 ( .A1(n_62), .A2(n_1063), .B(n_1066), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1087 ( .A1(n_62), .A2(n_101), .B1(n_577), .B2(n_1088), .C(n_1090), .Y(n_1087) );
INVx1_ASAP7_75t_L g790 ( .A(n_63), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g800 ( .A(n_64), .Y(n_800) );
INVxp67_ASAP7_75t_SL g1440 ( .A(n_65), .Y(n_1440) );
OAI22xp5_ASAP7_75t_L g1444 ( .A1(n_65), .A2(n_103), .B1(n_457), .B2(n_464), .Y(n_1444) );
AOI22xp33_ASAP7_75t_L g1906 ( .A1(n_66), .A2(n_88), .B1(n_722), .B2(n_1520), .Y(n_1906) );
INVxp67_ASAP7_75t_SL g1923 ( .A(n_66), .Y(n_1923) );
INVx1_ASAP7_75t_L g1129 ( .A(n_67), .Y(n_1129) );
INVx1_ASAP7_75t_L g613 ( .A(n_68), .Y(n_613) );
AOI21xp33_ASAP7_75t_L g1477 ( .A1(n_69), .A2(n_694), .B(n_695), .Y(n_1477) );
INVx1_ASAP7_75t_L g1484 ( .A(n_69), .Y(n_1484) );
XOR2x2_ASAP7_75t_L g1045 ( .A(n_70), .B(n_1046), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1955 ( .A1(n_71), .A2(n_336), .B1(n_625), .B2(n_1956), .Y(n_1955) );
AOI221xp5_ASAP7_75t_L g1963 ( .A1(n_71), .A2(n_353), .B1(n_667), .B2(n_694), .C(n_1964), .Y(n_1963) );
INVx1_ASAP7_75t_L g1004 ( .A(n_72), .Y(n_1004) );
INVx1_ASAP7_75t_L g1285 ( .A(n_73), .Y(n_1285) );
OAI22xp33_ASAP7_75t_L g1316 ( .A1(n_74), .A2(n_190), .B1(n_1317), .B2(n_1318), .Y(n_1316) );
OAI22xp5_ASAP7_75t_L g1360 ( .A1(n_74), .A2(n_190), .B1(n_1361), .B2(n_1363), .Y(n_1360) );
XNOR2xp5_ASAP7_75t_L g600 ( .A(n_75), .B(n_601), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g1705 ( .A1(n_76), .A2(n_365), .B1(n_1684), .B2(n_1689), .Y(n_1705) );
NAND2xp33_ASAP7_75t_SL g1427 ( .A(n_77), .B(n_771), .Y(n_1427) );
INVx1_ASAP7_75t_L g1453 ( .A(n_77), .Y(n_1453) );
OAI221xp5_ASAP7_75t_L g868 ( .A1(n_78), .A2(n_122), .B1(n_765), .B2(n_869), .C(n_870), .Y(n_868) );
INVx1_ASAP7_75t_L g899 ( .A(n_78), .Y(n_899) );
AOI22xp33_ASAP7_75t_SL g1609 ( .A1(n_79), .A2(n_370), .B1(n_480), .B2(n_743), .Y(n_1609) );
AOI221xp5_ASAP7_75t_L g1618 ( .A1(n_79), .A2(n_208), .B1(n_762), .B2(n_886), .C(n_1619), .Y(n_1618) );
OAI22xp33_ASAP7_75t_L g487 ( .A1(n_80), .A2(n_205), .B1(n_488), .B2(n_491), .Y(n_487) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_80), .Y(n_544) );
INVx1_ASAP7_75t_L g1337 ( .A(n_81), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1656 ( .A1(n_82), .A2(n_209), .B1(n_648), .B2(n_650), .Y(n_1656) );
INVx1_ASAP7_75t_L g872 ( .A(n_83), .Y(n_872) );
OAI221xp5_ASAP7_75t_SL g907 ( .A1(n_83), .A2(n_117), .B1(n_443), .B2(n_611), .C(n_815), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g1663 ( .A1(n_84), .A2(n_290), .B1(n_639), .B2(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1645 ( .A(n_85), .Y(n_1645) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_86), .A2(n_218), .B1(n_457), .B2(n_464), .Y(n_1051) );
INVxp67_ASAP7_75t_SL g1086 ( .A(n_86), .Y(n_1086) );
INVx1_ASAP7_75t_L g1102 ( .A(n_87), .Y(n_1102) );
AOI22xp5_ASAP7_75t_SL g1706 ( .A1(n_89), .A2(n_223), .B1(n_1692), .B2(n_1701), .Y(n_1706) );
AND2x2_ASAP7_75t_L g485 ( .A(n_90), .B(n_486), .Y(n_485) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_90), .A2(n_230), .B1(n_580), .B2(n_581), .C(n_583), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_91), .A2(n_108), .B1(n_722), .B2(n_723), .C(n_725), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_91), .A2(n_288), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_92), .A2(n_333), .B1(n_486), .B2(n_709), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_92), .A2(n_137), .B1(n_1135), .B2(n_1139), .Y(n_1138) );
AOI222xp33_ASAP7_75t_L g1067 ( .A1(n_93), .A2(n_151), .B1(n_352), .B2(n_466), .C1(n_620), .C2(n_962), .Y(n_1067) );
INVx1_ASAP7_75t_L g1092 ( .A(n_93), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_94), .B(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_94), .A2(n_173), .B1(n_576), .B2(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g1378 ( .A(n_95), .Y(n_1378) );
AOI221xp5_ASAP7_75t_L g1397 ( .A1(n_95), .A2(n_199), .B1(n_1398), .B2(n_1400), .C(n_1402), .Y(n_1397) );
INVx1_ASAP7_75t_L g1108 ( .A(n_96), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_97), .A2(n_200), .B1(n_625), .B2(n_626), .Y(n_624) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_97), .Y(n_689) );
INVxp67_ASAP7_75t_SL g1262 ( .A(n_98), .Y(n_1262) );
AOI22xp33_ASAP7_75t_SL g1290 ( .A1(n_98), .A2(n_297), .B1(n_480), .B2(n_639), .Y(n_1290) );
INVx1_ASAP7_75t_L g1340 ( .A(n_99), .Y(n_1340) );
OAI221xp5_ASAP7_75t_L g1938 ( .A1(n_100), .A2(n_239), .B1(n_1296), .B2(n_1939), .C(n_1940), .Y(n_1938) );
OAI211xp5_ASAP7_75t_L g1961 ( .A1(n_100), .A2(n_677), .B(n_1962), .C(n_1965), .Y(n_1961) );
AOI221xp5_ASAP7_75t_L g1053 ( .A1(n_101), .A2(n_233), .B1(n_1054), .B2(n_1056), .C(n_1058), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1668 ( .A1(n_102), .A2(n_293), .B1(n_629), .B2(n_632), .Y(n_1668) );
INVxp67_ASAP7_75t_SL g1456 ( .A(n_103), .Y(n_1456) );
INVx1_ASAP7_75t_L g382 ( .A(n_104), .Y(n_382) );
OAI221xp5_ASAP7_75t_L g1443 ( .A1(n_105), .A2(n_132), .B1(n_440), .B2(n_445), .C(n_451), .Y(n_1443) );
AOI221xp5_ASAP7_75t_L g891 ( .A1(n_106), .A2(n_152), .B1(n_762), .B2(n_886), .C(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g913 ( .A(n_106), .Y(n_913) );
INVx1_ASAP7_75t_L g1049 ( .A(n_107), .Y(n_1049) );
OAI21xp33_ASAP7_75t_L g1074 ( .A1(n_107), .A2(n_521), .B(n_1075), .Y(n_1074) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_108), .A2(n_158), .B1(n_760), .B2(n_762), .C(n_763), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g1959 ( .A1(n_109), .A2(n_276), .B1(n_648), .B2(n_650), .Y(n_1959) );
INVx1_ASAP7_75t_L g1161 ( .A(n_110), .Y(n_1161) );
INVx1_ASAP7_75t_L g1571 ( .A(n_112), .Y(n_1571) );
AOI22xp33_ASAP7_75t_L g1586 ( .A1(n_112), .A2(n_162), .B1(n_526), .B2(n_779), .Y(n_1586) );
AOI22xp5_ASAP7_75t_L g1708 ( .A1(n_113), .A2(n_340), .B1(n_1689), .B2(n_1701), .Y(n_1708) );
AOI22xp33_ASAP7_75t_SL g1111 ( .A1(n_114), .A2(n_121), .B1(n_1112), .B2(n_1114), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1132 ( .A1(n_114), .A2(n_324), .B1(n_547), .B2(n_577), .C(n_667), .Y(n_1132) );
INVx1_ASAP7_75t_L g1434 ( .A(n_115), .Y(n_1434) );
INVx1_ASAP7_75t_L g1899 ( .A(n_116), .Y(n_1899) );
OAI221xp5_ASAP7_75t_L g1920 ( .A1(n_116), .A2(n_124), .B1(n_1252), .B2(n_1269), .C(n_1921), .Y(n_1920) );
INVx1_ASAP7_75t_L g881 ( .A(n_117), .Y(n_881) );
CKINVDCx5p33_ASAP7_75t_R g1560 ( .A(n_118), .Y(n_1560) );
INVx1_ASAP7_75t_L g938 ( .A(n_119), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g985 ( .A1(n_119), .A2(n_257), .B1(n_986), .B2(n_988), .Y(n_985) );
INVx1_ASAP7_75t_L g1277 ( .A(n_120), .Y(n_1277) );
INVx1_ASAP7_75t_L g897 ( .A(n_122), .Y(n_897) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_123), .A2(n_200), .B1(n_660), .B2(n_665), .C(n_667), .Y(n_659) );
INVx1_ASAP7_75t_L g1898 ( .A(n_124), .Y(n_1898) );
OAI21xp5_ASAP7_75t_SL g1146 ( .A1(n_125), .A2(n_648), .B(n_1147), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1471 ( .A1(n_126), .A2(n_247), .B1(n_581), .B2(n_780), .Y(n_1471) );
INVx1_ASAP7_75t_L g1488 ( .A(n_126), .Y(n_1488) );
XOR2x2_ASAP7_75t_L g1591 ( .A(n_127), .B(n_1592), .Y(n_1591) );
OAI221xp5_ASAP7_75t_L g1553 ( .A1(n_128), .A2(n_302), .B1(n_457), .B2(n_464), .C(n_1554), .Y(n_1553) );
INVx1_ASAP7_75t_L g1589 ( .A(n_128), .Y(n_1589) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_129), .A2(n_787), .B1(n_788), .B2(n_856), .Y(n_786) );
INVx1_ASAP7_75t_L g856 ( .A(n_129), .Y(n_856) );
INVx1_ASAP7_75t_L g876 ( .A(n_130), .Y(n_876) );
OAI21xp33_ASAP7_75t_L g905 ( .A1(n_130), .A2(n_643), .B(n_906), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g1511 ( .A(n_131), .Y(n_1511) );
INVxp67_ASAP7_75t_SL g1439 ( .A(n_132), .Y(n_1439) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_133), .A2(n_331), .B1(n_440), .B2(n_445), .C(n_451), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_133), .B(n_552), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g1435 ( .A1(n_134), .A2(n_140), .B1(n_557), .B2(n_1430), .C(n_1436), .Y(n_1435) );
AOI22xp33_ASAP7_75t_SL g1009 ( .A1(n_135), .A2(n_266), .B1(n_780), .B2(n_894), .Y(n_1009) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_135), .A2(n_350), .B1(n_480), .B2(n_722), .C(n_725), .Y(n_1030) );
OAI22xp33_ASAP7_75t_L g1211 ( .A1(n_136), .A2(n_338), .B1(n_1212), .B2(n_1213), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_136), .A2(n_338), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1119 ( .A1(n_137), .A2(n_324), .B1(n_625), .B2(n_1114), .C(n_1120), .Y(n_1119) );
CKINVDCx5p33_ASAP7_75t_R g1594 ( .A(n_138), .Y(n_1594) );
AOI22xp33_ASAP7_75t_SL g1519 ( .A1(n_139), .A2(n_320), .B1(n_1295), .B2(n_1520), .Y(n_1519) );
AOI22xp33_ASAP7_75t_L g1538 ( .A1(n_139), .A2(n_308), .B1(n_580), .B2(n_581), .Y(n_1538) );
INVx1_ASAP7_75t_L g1450 ( .A(n_140), .Y(n_1450) );
AOI22xp33_ASAP7_75t_L g1904 ( .A1(n_141), .A2(n_170), .B1(n_935), .B2(n_1903), .Y(n_1904) );
INVx1_ASAP7_75t_L g1948 ( .A(n_142), .Y(n_1948) );
INVx1_ASAP7_75t_L g1258 ( .A(n_143), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_143), .A2(n_214), .B1(n_486), .B2(n_1029), .Y(n_1291) );
INVx1_ASAP7_75t_L g1599 ( .A(n_144), .Y(n_1599) );
AOI22xp33_ASAP7_75t_L g1523 ( .A1(n_145), .A2(n_332), .B1(n_486), .B2(n_620), .Y(n_1523) );
INVx1_ASAP7_75t_L g744 ( .A(n_146), .Y(n_744) );
AOI221xp5_ASAP7_75t_SL g885 ( .A1(n_147), .A2(n_329), .B1(n_762), .B2(n_886), .C(n_889), .Y(n_885) );
INVx1_ASAP7_75t_L g922 ( .A(n_147), .Y(n_922) );
OAI222xp33_ASAP7_75t_L g641 ( .A1(n_148), .A2(n_254), .B1(n_261), .B2(n_642), .C1(n_648), .C2(n_650), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g654 ( .A1(n_148), .A2(n_655), .B(n_658), .C(n_670), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_149), .Y(n_883) );
OAI22xp33_ASAP7_75t_L g1907 ( .A1(n_150), .A2(n_299), .B1(n_1671), .B2(n_1908), .Y(n_1907) );
INVx1_ASAP7_75t_L g1919 ( .A(n_150), .Y(n_1919) );
INVx1_ASAP7_75t_L g1083 ( .A(n_151), .Y(n_1083) );
INVx1_ASAP7_75t_L g926 ( .A(n_152), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1604 ( .A1(n_153), .A2(n_323), .B1(n_634), .B2(n_1029), .Y(n_1604) );
AOI22xp33_ASAP7_75t_L g1620 ( .A1(n_153), .A2(n_277), .B1(n_839), .B2(n_1621), .Y(n_1620) );
AOI221xp5_ASAP7_75t_L g1470 ( .A1(n_154), .A2(n_366), .B1(n_564), .B2(n_892), .C(n_1141), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g1492 ( .A1(n_154), .A2(n_264), .B1(n_480), .B2(n_626), .Y(n_1492) );
INVxp67_ASAP7_75t_SL g1943 ( .A(n_155), .Y(n_1943) );
AOI221xp5_ASAP7_75t_L g1973 ( .A1(n_155), .A2(n_263), .B1(n_578), .B2(n_889), .C(n_1964), .Y(n_1973) );
INVx1_ASAP7_75t_L g1556 ( .A(n_156), .Y(n_1556) );
OAI22xp5_ASAP7_75t_L g1583 ( .A1(n_156), .A2(n_346), .B1(n_531), .B2(n_540), .Y(n_1583) );
CKINVDCx5p33_ASAP7_75t_R g950 ( .A(n_157), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_158), .A2(n_189), .B1(n_712), .B2(n_713), .C(n_716), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g1379 ( .A1(n_159), .A2(n_199), .B1(n_935), .B2(n_1380), .C(n_1382), .Y(n_1379) );
INVx1_ASAP7_75t_L g1408 ( .A(n_159), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_160), .A2(n_359), .B1(n_632), .B2(n_634), .Y(n_631) );
INVxp67_ASAP7_75t_SL g795 ( .A(n_161), .Y(n_795) );
OAI221xp5_ASAP7_75t_L g811 ( .A1(n_161), .A2(n_451), .B1(n_457), .B2(n_812), .C(n_821), .Y(n_811) );
INVx1_ASAP7_75t_L g1566 ( .A(n_162), .Y(n_1566) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_163), .A2(n_632), .B(n_716), .Y(n_809) );
INVx1_ASAP7_75t_L g836 ( .A(n_163), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g1911 ( .A1(n_164), .A2(n_185), .B1(n_648), .B2(n_792), .Y(n_1911) );
OAI211xp5_ASAP7_75t_L g1913 ( .A1(n_164), .A2(n_1616), .B(n_1914), .C(n_1917), .Y(n_1913) );
INVx1_ASAP7_75t_L g820 ( .A(n_165), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_165), .A2(n_234), .B1(n_839), .B2(n_840), .Y(n_838) );
INVx1_ASAP7_75t_L g1958 ( .A(n_166), .Y(n_1958) );
INVx1_ASAP7_75t_L g1762 ( .A(n_167), .Y(n_1762) );
AOI22xp5_ASAP7_75t_SL g1723 ( .A1(n_168), .A2(n_179), .B1(n_1692), .B2(n_1701), .Y(n_1723) );
AOI22xp33_ASAP7_75t_SL g1133 ( .A1(n_169), .A2(n_333), .B1(n_1134), .B2(n_1135), .Y(n_1133) );
AOI221xp5_ASAP7_75t_L g1924 ( .A1(n_170), .A2(n_274), .B1(n_762), .B2(n_886), .C(n_1260), .Y(n_1924) );
INVx1_ASAP7_75t_L g605 ( .A(n_171), .Y(n_605) );
OAI221xp5_ASAP7_75t_SL g676 ( .A1(n_171), .A2(n_180), .B1(n_677), .B2(n_681), .C(n_685), .Y(n_676) );
INVx1_ASAP7_75t_L g1200 ( .A(n_172), .Y(n_1200) );
OAI211xp5_ASAP7_75t_L g1224 ( .A1(n_172), .A2(n_1173), .B(n_1225), .C(n_1227), .Y(n_1224) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_173), .A2(n_213), .B1(n_495), .B2(n_500), .C(n_501), .Y(n_494) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_174), .A2(n_175), .B1(n_735), .B2(n_736), .C(n_740), .Y(n_734) );
INVxp67_ASAP7_75t_SL g756 ( .A(n_175), .Y(n_756) );
INVxp33_ASAP7_75t_SL g766 ( .A(n_176), .Y(n_766) );
INVx1_ASAP7_75t_L g438 ( .A(n_177), .Y(n_438) );
INVx1_ASAP7_75t_L g953 ( .A(n_178), .Y(n_953) );
INVx1_ASAP7_75t_L g608 ( .A(n_180), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g1932 ( .A1(n_181), .A2(n_1933), .B1(n_1934), .B2(n_1976), .Y(n_1932) );
CKINVDCx5p33_ASAP7_75t_R g1976 ( .A(n_181), .Y(n_1976) );
INVx2_ASAP7_75t_L g1687 ( .A(n_182), .Y(n_1687) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_182), .B(n_1688), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1695 ( .A(n_182), .B(n_316), .Y(n_1695) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_183), .A2(n_480), .B(n_482), .Y(n_479) );
INVx1_ASAP7_75t_L g567 ( .A(n_183), .Y(n_567) );
INVxp67_ASAP7_75t_SL g1268 ( .A(n_184), .Y(n_1268) );
AOI22xp33_ASAP7_75t_SL g1294 ( .A1(n_184), .A2(n_334), .B1(n_942), .B2(n_1295), .Y(n_1294) );
XNOR2xp5_ASAP7_75t_L g1460 ( .A(n_186), .B(n_1461), .Y(n_1460) );
AOI22xp5_ASAP7_75t_SL g1719 ( .A1(n_186), .A2(n_265), .B1(n_1689), .B2(n_1694), .Y(n_1719) );
OAI211xp5_ASAP7_75t_L g1421 ( .A1(n_187), .A2(n_748), .B(n_1422), .C(n_1437), .Y(n_1421) );
INVx1_ASAP7_75t_L g1570 ( .A(n_188), .Y(n_1570) );
INVx1_ASAP7_75t_L g774 ( .A(n_189), .Y(n_774) );
INVx1_ASAP7_75t_L g1590 ( .A(n_191), .Y(n_1590) );
OAI21xp33_ASAP7_75t_L g1001 ( .A1(n_193), .A2(n_751), .B(n_1002), .Y(n_1001) );
OAI221xp5_ASAP7_75t_L g1035 ( .A1(n_193), .A2(n_301), .B1(n_824), .B2(n_1036), .C(n_1037), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1691 ( .A1(n_194), .A2(n_335), .B1(n_1692), .B2(n_1694), .Y(n_1691) );
XOR2x2_ASAP7_75t_L g1893 ( .A(n_194), .B(n_1894), .Y(n_1893) );
AOI22xp33_ASAP7_75t_L g1928 ( .A1(n_194), .A2(n_1929), .B1(n_1932), .B2(n_1977), .Y(n_1928) );
INVx1_ASAP7_75t_L g912 ( .A(n_195), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g1699 ( .A1(n_196), .A2(n_271), .B1(n_1684), .B2(n_1689), .Y(n_1699) );
OAI221xp5_ASAP7_75t_L g1388 ( .A1(n_197), .A2(n_294), .B1(n_440), .B2(n_445), .C(n_451), .Y(n_1388) );
INVx1_ASAP7_75t_L g1413 ( .A(n_197), .Y(n_1413) );
INVx1_ASAP7_75t_L g1159 ( .A(n_198), .Y(n_1159) );
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_201), .Y(n_947) );
INVx1_ASAP7_75t_L g957 ( .A(n_202), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g1709 ( .A1(n_203), .A2(n_295), .B1(n_1684), .B2(n_1692), .Y(n_1709) );
INVxp67_ASAP7_75t_SL g1651 ( .A(n_204), .Y(n_1651) );
INVx1_ASAP7_75t_L g411 ( .A(n_205), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g1517 ( .A(n_206), .Y(n_1517) );
INVx1_ASAP7_75t_L g742 ( .A(n_207), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_207), .A2(n_245), .B1(n_531), .B2(n_540), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g1603 ( .A1(n_208), .A2(n_219), .B1(n_480), .B2(n_743), .Y(n_1603) );
OAI211xp5_ASAP7_75t_L g1636 ( .A1(n_209), .A2(n_655), .B(n_1637), .C(n_1644), .Y(n_1636) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_210), .Y(n_823) );
INVx1_ASAP7_75t_L g1457 ( .A(n_211), .Y(n_1457) );
AOI22xp33_ASAP7_75t_SL g1008 ( .A1(n_212), .A2(n_339), .B1(n_576), .B2(n_888), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1028 ( .A1(n_212), .A2(n_240), .B1(n_716), .B2(n_722), .C(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g569 ( .A(n_213), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_214), .A2(n_371), .B1(n_984), .B2(n_1274), .Y(n_1273) );
AOI22xp33_ASAP7_75t_SL g1524 ( .A1(n_215), .A2(n_308), .B1(n_615), .B2(n_1295), .Y(n_1524) );
AOI221xp5_ASAP7_75t_L g1531 ( .A1(n_215), .A2(n_320), .B1(n_577), .B2(n_667), .C(n_1532), .Y(n_1531) );
INVx2_ASAP7_75t_L g437 ( .A(n_216), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_216), .B(n_435), .Y(n_460) );
INVx1_ASAP7_75t_L g506 ( .A(n_216), .Y(n_506) );
INVx1_ASAP7_75t_L g1500 ( .A(n_217), .Y(n_1500) );
INVxp67_ASAP7_75t_SL g1070 ( .A(n_218), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1630 ( .A1(n_219), .A2(n_370), .B1(n_894), .B2(n_1621), .Y(n_1630) );
XOR2xp5_ASAP7_75t_L g928 ( .A(n_220), .B(n_929), .Y(n_928) );
OAI221xp5_ASAP7_75t_SL g1647 ( .A1(n_221), .A2(n_317), .B1(n_1252), .B2(n_1626), .C(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1660 ( .A(n_221), .Y(n_1660) );
INVx1_ASAP7_75t_L g1574 ( .A(n_222), .Y(n_1574) );
AOI22xp33_ASAP7_75t_L g1588 ( .A1(n_222), .A2(n_342), .B1(n_580), .B2(n_581), .Y(n_1588) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_224), .A2(n_328), .B1(n_498), .B2(n_714), .Y(n_939) );
INVx1_ASAP7_75t_L g992 ( .A(n_224), .Y(n_992) );
INVx1_ASAP7_75t_L g923 ( .A(n_225), .Y(n_923) );
INVx1_ASAP7_75t_L g1331 ( .A(n_226), .Y(n_1331) );
CKINVDCx5p33_ASAP7_75t_R g1528 ( .A(n_227), .Y(n_1528) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_228), .A2(n_349), .B1(n_894), .B2(n_1015), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_228), .A2(n_266), .B1(n_480), .B2(n_503), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1595 ( .A1(n_229), .A2(n_322), .B1(n_792), .B2(n_1502), .Y(n_1595) );
OAI211xp5_ASAP7_75t_L g1615 ( .A1(n_229), .A2(n_1616), .B(n_1617), .C(n_1622), .Y(n_1615) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_230), .A2(n_284), .B1(n_473), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g1256 ( .A(n_231), .Y(n_1256) );
AOI22xp33_ASAP7_75t_SL g1292 ( .A1(n_231), .A2(n_371), .B1(n_486), .B2(n_1293), .Y(n_1292) );
BUFx3_ASAP7_75t_L g429 ( .A(n_232), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_233), .B(n_693), .Y(n_1080) );
INVx1_ASAP7_75t_L g1059 ( .A(n_235), .Y(n_1059) );
OAI21xp5_ASAP7_75t_SL g1540 ( .A1(n_236), .A2(n_648), .B(n_1541), .Y(n_1540) );
INVx1_ASAP7_75t_L g1003 ( .A(n_237), .Y(n_1003) );
OAI21xp5_ASAP7_75t_SL g1278 ( .A1(n_238), .A2(n_648), .B(n_1279), .Y(n_1278) );
OAI221xp5_ASAP7_75t_SL g1966 ( .A1(n_239), .A2(n_345), .B1(n_1269), .B2(n_1967), .C(n_1969), .Y(n_1966) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_240), .A2(n_350), .B1(n_1018), .B2(n_1019), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g1683 ( .A1(n_241), .A2(n_292), .B1(n_1684), .B2(n_1689), .Y(n_1683) );
XOR2xp5_ASAP7_75t_L g1633 ( .A(n_242), .B(n_1634), .Y(n_1633) );
AOI22xp33_ASAP7_75t_L g1642 ( .A1(n_243), .A2(n_293), .B1(n_1015), .B2(n_1643), .Y(n_1642) );
OAI22xp33_ASAP7_75t_L g1610 ( .A1(n_244), .A2(n_364), .B1(n_1611), .B2(n_1613), .Y(n_1610) );
INVx1_ASAP7_75t_L g1623 ( .A(n_244), .Y(n_1623) );
INVx1_ASAP7_75t_L g727 ( .A(n_245), .Y(n_727) );
OAI211xp5_ASAP7_75t_SL g1309 ( .A1(n_246), .A2(n_1225), .B(n_1310), .C(n_1312), .Y(n_1309) );
INVx1_ASAP7_75t_L g1357 ( .A(n_246), .Y(n_1357) );
INVx1_ASAP7_75t_L g1491 ( .A(n_247), .Y(n_1491) );
CKINVDCx5p33_ASAP7_75t_R g1655 ( .A(n_248), .Y(n_1655) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_249), .Y(n_794) );
INVx1_ASAP7_75t_L g1315 ( .A(n_250), .Y(n_1315) );
OAI211xp5_ASAP7_75t_SL g1353 ( .A1(n_250), .A2(n_1193), .B(n_1354), .C(n_1355), .Y(n_1353) );
INVx1_ASAP7_75t_L g1438 ( .A(n_251), .Y(n_1438) );
INVx1_ASAP7_75t_L g470 ( .A(n_252), .Y(n_470) );
INVx1_ASAP7_75t_L g1276 ( .A(n_253), .Y(n_1276) );
AOI22xp33_ASAP7_75t_L g1605 ( .A1(n_255), .A2(n_277), .B1(n_1029), .B2(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1628 ( .A(n_255), .Y(n_1628) );
OAI211xp5_ASAP7_75t_L g1557 ( .A1(n_256), .A2(n_426), .B(n_451), .C(n_1558), .Y(n_1557) );
INVxp33_ASAP7_75t_SL g1582 ( .A(n_256), .Y(n_1582) );
OAI221xp5_ASAP7_75t_L g943 ( .A1(n_257), .A2(n_281), .B1(n_443), .B2(n_611), .C(n_914), .Y(n_943) );
INVx1_ASAP7_75t_L g1468 ( .A(n_258), .Y(n_1468) );
INVx1_ASAP7_75t_L g1107 ( .A(n_259), .Y(n_1107) );
BUFx3_ASAP7_75t_L g399 ( .A(n_260), .Y(n_399) );
INVx1_ASAP7_75t_L g419 ( .A(n_260), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g1270 ( .A1(n_262), .A2(n_655), .B(n_1271), .C(n_1275), .Y(n_1270) );
INVx1_ASAP7_75t_L g1287 ( .A(n_262), .Y(n_1287) );
INVx1_ASAP7_75t_L g1951 ( .A(n_263), .Y(n_1951) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_267), .B(n_853), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_268), .Y(n_965) );
INVxp67_ASAP7_75t_SL g512 ( .A(n_269), .Y(n_512) );
OAI322xp33_ASAP7_75t_SL g1941 ( .A1(n_270), .A2(n_1169), .A3(n_1342), .B1(n_1611), .B2(n_1942), .C1(n_1947), .C2(n_1950), .Y(n_1941) );
OAI22xp33_ASAP7_75t_SL g1974 ( .A1(n_270), .A2(n_276), .B1(n_655), .B2(n_1975), .Y(n_1974) );
INVxp67_ASAP7_75t_SL g995 ( .A(n_271), .Y(n_995) );
CKINVDCx5p33_ASAP7_75t_R g871 ( .A(n_272), .Y(n_871) );
INVx1_ASAP7_75t_L g802 ( .A(n_273), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g1104 ( .A(n_275), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1375 ( .A1(n_278), .A2(n_348), .B1(n_625), .B2(n_935), .C(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1403 ( .A(n_278), .Y(n_1403) );
INVx1_ASAP7_75t_L g1377 ( .A(n_279), .Y(n_1377) );
INVx1_ASAP7_75t_L g1954 ( .A(n_280), .Y(n_1954) );
OA222x2_ASAP7_75t_L g989 ( .A1(n_281), .A2(n_298), .B1(n_354), .B2(n_521), .C1(n_751), .C2(n_754), .Y(n_989) );
INVx1_ASAP7_75t_L g1172 ( .A(n_283), .Y(n_1172) );
AOI32xp33_ASAP7_75t_L g546 ( .A1(n_284), .A2(n_547), .A3(n_550), .B1(n_555), .B2(n_1983), .Y(n_546) );
XNOR2x2_ASAP7_75t_L g1370 ( .A(n_285), .B(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1060 ( .A(n_286), .Y(n_1060) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_287), .Y(n_816) );
XOR2x2_ASAP7_75t_L g1248 ( .A(n_289), .B(n_1249), .Y(n_1248) );
INVxp67_ASAP7_75t_SL g1649 ( .A(n_290), .Y(n_1649) );
INVxp67_ASAP7_75t_SL g1393 ( .A(n_294), .Y(n_1393) );
INVx1_ASAP7_75t_L g432 ( .A(n_296), .Y(n_432) );
INVx1_ASAP7_75t_L g450 ( .A(n_296), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g1272 ( .A1(n_297), .A2(n_334), .B1(n_547), .B2(n_886), .C(n_892), .Y(n_1272) );
INVx1_ASAP7_75t_L g941 ( .A(n_298), .Y(n_941) );
INVx1_ASAP7_75t_L g1918 ( .A(n_299), .Y(n_1918) );
INVx1_ASAP7_75t_L g1012 ( .A(n_300), .Y(n_1012) );
INVxp67_ASAP7_75t_SL g1042 ( .A(n_301), .Y(n_1042) );
INVxp67_ASAP7_75t_SL g1580 ( .A(n_302), .Y(n_1580) );
INVx1_ASAP7_75t_L g1396 ( .A(n_303), .Y(n_1396) );
OAI22xp5_ASAP7_75t_L g1374 ( .A1(n_304), .A2(n_341), .B1(n_488), .B2(n_491), .Y(n_1374) );
INVx1_ASAP7_75t_L g1394 ( .A(n_304), .Y(n_1394) );
INVx1_ASAP7_75t_L g1333 ( .A(n_305), .Y(n_1333) );
INVxp67_ASAP7_75t_SL g1073 ( .A(n_306), .Y(n_1073) );
INVx1_ASAP7_75t_L g1166 ( .A(n_307), .Y(n_1166) );
INVx1_ASAP7_75t_L g1334 ( .A(n_309), .Y(n_1334) );
INVx1_ASAP7_75t_L g741 ( .A(n_310), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_310), .B(n_748), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g1529 ( .A(n_311), .Y(n_1529) );
INVx1_ASAP7_75t_L g1328 ( .A(n_312), .Y(n_1328) );
CKINVDCx5p33_ASAP7_75t_R g1475 ( .A(n_313), .Y(n_1475) );
INVx1_ASAP7_75t_L g826 ( .A(n_314), .Y(n_826) );
INVx1_ASAP7_75t_L g618 ( .A(n_315), .Y(n_618) );
INVx1_ASAP7_75t_L g1688 ( .A(n_316), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_316), .B(n_1687), .Y(n_1693) );
INVx1_ASAP7_75t_L g1661 ( .A(n_317), .Y(n_1661) );
CKINVDCx5p33_ASAP7_75t_R g1281 ( .A(n_318), .Y(n_1281) );
XNOR2xp5_ASAP7_75t_L g1098 ( .A(n_319), .B(n_1099), .Y(n_1098) );
OAI22xp33_ASAP7_75t_L g1305 ( .A1(n_321), .A2(n_374), .B1(n_1306), .B2(n_1308), .Y(n_1305) );
OAI22xp33_ASAP7_75t_L g1365 ( .A1(n_321), .A2(n_374), .B1(n_391), .B2(n_1366), .Y(n_1365) );
AOI21xp33_ASAP7_75t_L g1629 ( .A1(n_323), .A2(n_886), .B(n_889), .Y(n_1629) );
INVx1_ASAP7_75t_L g1433 ( .A(n_325), .Y(n_1433) );
AOI221xp5_ASAP7_75t_L g1446 ( .A1(n_325), .A2(n_375), .B1(n_472), .B2(n_710), .C(n_1447), .Y(n_1446) );
INVx1_ASAP7_75t_L g1163 ( .A(n_326), .Y(n_1163) );
INVx1_ASAP7_75t_L g1764 ( .A(n_327), .Y(n_1764) );
INVx1_ASAP7_75t_L g991 ( .A(n_328), .Y(n_991) );
INVx1_ASAP7_75t_L g916 ( .A(n_329), .Y(n_916) );
INVxp67_ASAP7_75t_SL g538 ( .A(n_331), .Y(n_538) );
INVxp67_ASAP7_75t_SL g1972 ( .A(n_336), .Y(n_1972) );
INVx1_ASAP7_75t_L g803 ( .A(n_337), .Y(n_803) );
OAI221xp5_ASAP7_75t_L g841 ( .A1(n_337), .A2(n_754), .B1(n_842), .B2(n_850), .C(n_851), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_339), .A2(n_349), .B1(n_503), .B2(n_1032), .Y(n_1031) );
INVxp67_ASAP7_75t_SL g1411 ( .A(n_341), .Y(n_1411) );
INVx1_ASAP7_75t_L g1567 ( .A(n_342), .Y(n_1567) );
INVx1_ASAP7_75t_L g1314 ( .A(n_343), .Y(n_1314) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_344), .Y(n_395) );
INVxp67_ASAP7_75t_SL g1936 ( .A(n_345), .Y(n_1936) );
INVx1_ASAP7_75t_L g1559 ( .A(n_346), .Y(n_1559) );
CKINVDCx5p33_ASAP7_75t_R g1514 ( .A(n_347), .Y(n_1514) );
INVx1_ASAP7_75t_L g1407 ( .A(n_348), .Y(n_1407) );
AOI21xp33_ASAP7_75t_L g1084 ( .A1(n_352), .A2(n_547), .B(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1949 ( .A(n_353), .Y(n_1949) );
INVx1_ASAP7_75t_L g936 ( .A(n_354), .Y(n_936) );
INVx1_ASAP7_75t_L g784 ( .A(n_355), .Y(n_784) );
XOR2xp5_ASAP7_75t_L g1507 ( .A(n_356), .B(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g416 ( .A(n_357), .Y(n_416) );
INVx2_ASAP7_75t_L g510 ( .A(n_357), .Y(n_510) );
INVx1_ASAP7_75t_L g525 ( .A(n_357), .Y(n_525) );
XOR2x2_ASAP7_75t_L g1152 ( .A(n_358), .B(n_1153), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_359), .A2(n_362), .B1(n_547), .B2(n_693), .C(n_695), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g1910 ( .A(n_360), .Y(n_1910) );
INVx1_ASAP7_75t_L g1384 ( .A(n_361), .Y(n_1384) );
INVx1_ASAP7_75t_L g1076 ( .A(n_363), .Y(n_1076) );
INVx1_ASAP7_75t_L g1624 ( .A(n_364), .Y(n_1624) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_367), .Y(n_805) );
OAI21xp33_ASAP7_75t_SL g1551 ( .A1(n_368), .A2(n_748), .B(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_L g1555 ( .A(n_368), .Y(n_1555) );
INVx1_ASAP7_75t_L g1174 ( .A(n_369), .Y(n_1174) );
INVx1_ASAP7_75t_L g1946 ( .A(n_372), .Y(n_1946) );
INVx1_ASAP7_75t_L g1330 ( .A(n_373), .Y(n_1330) );
INVx1_ASAP7_75t_L g1426 ( .A(n_375), .Y(n_1426) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_400), .B(n_1675), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_385), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g1927 ( .A(n_379), .B(n_388), .Y(n_1927) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1931 ( .A(n_381), .B(n_384), .Y(n_1931) );
INVx1_ASAP7_75t_L g1979 ( .A(n_381), .Y(n_1979) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g1981 ( .A(n_384), .B(n_1979), .Y(n_1981) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g1216 ( .A(n_388), .B(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g587 ( .A(n_389), .B(n_399), .Y(n_587) );
AND2x4_ASAP7_75t_L g696 ( .A(n_389), .B(n_398), .Y(n_696) );
INVx1_ASAP7_75t_L g1212 ( .A(n_390), .Y(n_1212) );
AND2x4_ASAP7_75t_SL g1926 ( .A(n_390), .B(n_1927), .Y(n_1926) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_397), .Y(n_391) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_392), .Y(n_568) );
OR2x6_ASAP7_75t_L g1206 ( .A(n_392), .B(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g1327 ( .A(n_392), .Y(n_1327) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx4f_ASAP7_75t_L g688 ( .A(n_393), .Y(n_688) );
INVx3_ASAP7_75t_L g977 ( .A(n_393), .Y(n_977) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx2_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
AND2x2_ASAP7_75t_L g516 ( .A(n_395), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g529 ( .A(n_395), .Y(n_529) );
INVx1_ASAP7_75t_L g543 ( .A(n_395), .Y(n_543) );
AND2x2_ASAP7_75t_L g549 ( .A(n_395), .B(n_396), .Y(n_549) );
NAND2x1_ASAP7_75t_L g554 ( .A(n_395), .B(n_396), .Y(n_554) );
INVx1_ASAP7_75t_L g422 ( .A(n_396), .Y(n_422) );
INVx2_ASAP7_75t_L g517 ( .A(n_396), .Y(n_517) );
AND2x2_ASAP7_75t_L g528 ( .A(n_396), .B(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g537 ( .A(n_396), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_396), .B(n_529), .Y(n_574) );
OR2x2_ASAP7_75t_L g773 ( .A(n_396), .B(n_421), .Y(n_773) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g1195 ( .A(n_398), .Y(n_1195) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx2_ASAP7_75t_L g1199 ( .A(n_399), .Y(n_1199) );
AND2x4_ASAP7_75t_L g1203 ( .A(n_399), .B(n_542), .Y(n_1203) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_1148), .B2(n_1149), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_1095), .B2(n_1096), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
XNOR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_858), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_407), .B1(n_700), .B2(n_857), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OA22x2_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_599), .B2(n_600), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AO211x2_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_423), .C(n_518), .Y(n_410) );
INVx3_ASAP7_75t_L g748 ( .A(n_412), .Y(n_748) );
AOI222xp33_ASAP7_75t_L g789 ( .A1(n_412), .A2(n_513), .B1(n_790), .B2(n_791), .C1(n_794), .C2(n_795), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g990 ( .A1(n_412), .A2(n_513), .B1(n_991), .B2(n_992), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_412), .B(n_999), .Y(n_998) );
AOI211xp5_ASAP7_75t_L g1072 ( .A1(n_412), .A2(n_1073), .B(n_1074), .C(n_1078), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_412), .B(n_1411), .Y(n_1410) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_417), .Y(n_412) );
AND2x4_ASAP7_75t_L g513 ( .A(n_413), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g540 ( .A(n_414), .B(n_541), .Y(n_540) );
INVxp67_ASAP7_75t_L g651 ( .A(n_414), .Y(n_651) );
OR2x2_ASAP7_75t_L g988 ( .A(n_414), .B(n_541), .Y(n_988) );
INVx1_ASAP7_75t_L g1217 ( .A(n_414), .Y(n_1217) );
BUFx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g586 ( .A(n_415), .Y(n_586) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g672 ( .A(n_417), .Y(n_672) );
BUFx6f_ASAP7_75t_L g1128 ( .A(n_417), .Y(n_1128) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
AND2x2_ASAP7_75t_L g514 ( .A(n_418), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_418), .B(n_525), .Y(n_524) );
AND2x4_ASAP7_75t_L g656 ( .A(n_418), .B(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g675 ( .A(n_418), .B(n_515), .Y(n_675) );
AND2x4_ASAP7_75t_SL g680 ( .A(n_418), .B(n_548), .Y(n_680) );
BUFx2_ASAP7_75t_L g873 ( .A(n_418), .Y(n_873) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_418), .B(n_526), .Y(n_1465) );
HB1xp67_ASAP7_75t_L g1207 ( .A(n_419), .Y(n_1207) );
INVx3_ASAP7_75t_L g582 ( .A(n_420), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_420), .B(n_534), .Y(n_593) );
BUFx6f_ASAP7_75t_L g779 ( .A(n_420), .Y(n_779) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
A2O1A1Ixp33_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_467), .B(n_507), .C(n_511), .Y(n_423) );
AOI211xp5_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_438), .B(n_439), .C(n_456), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_425), .A2(n_731), .B1(n_734), .B2(n_744), .Y(n_730) );
INVx2_ASAP7_75t_L g1039 ( .A(n_425), .Y(n_1039) );
AOI211xp5_ASAP7_75t_SL g1048 ( .A1(n_425), .A2(n_1049), .B(n_1050), .C(n_1051), .Y(n_1048) );
AOI211xp5_ASAP7_75t_SL g1385 ( .A1(n_425), .A2(n_1386), .B(n_1387), .C(n_1388), .Y(n_1385) );
AOI211xp5_ASAP7_75t_SL g1442 ( .A1(n_425), .A2(n_1438), .B(n_1443), .C(n_1444), .Y(n_1442) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OR2x6_ASAP7_75t_L g650 ( .A(n_426), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g792 ( .A(n_426), .B(n_651), .Y(n_792) );
NAND2x1p5_ASAP7_75t_L g426 ( .A(n_427), .B(n_433), .Y(n_426) );
INVx8_ASAP7_75t_L g481 ( .A(n_427), .Y(n_481) );
AND2x2_ASAP7_75t_L g489 ( .A(n_427), .B(n_490), .Y(n_489) );
BUFx3_ASAP7_75t_L g709 ( .A(n_427), .Y(n_709) );
BUFx3_ASAP7_75t_L g724 ( .A(n_427), .Y(n_724) );
AND2x4_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
AND2x4_ASAP7_75t_L g462 ( .A(n_428), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_429), .Y(n_444) );
AND2x4_ASAP7_75t_L g493 ( .A(n_429), .B(n_449), .Y(n_493) );
OR2x2_ASAP7_75t_L g499 ( .A(n_429), .B(n_431), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_429), .B(n_450), .Y(n_646) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g463 ( .A(n_432), .Y(n_463) );
AND2x6_ASAP7_75t_L g441 ( .A(n_433), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g446 ( .A(n_433), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g455 ( .A(n_433), .Y(n_455) );
AND2x4_ASAP7_75t_L g607 ( .A(n_433), .B(n_591), .Y(n_607) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g505 ( .A(n_434), .B(n_506), .Y(n_505) );
NAND3x1_ASAP7_75t_L g636 ( .A(n_434), .B(n_506), .C(n_637), .Y(n_636) );
OR2x4_ASAP7_75t_L g1220 ( .A(n_434), .B(n_499), .Y(n_1220) );
INVx1_ASAP7_75t_L g1223 ( .A(n_434), .Y(n_1223) );
AND2x4_ASAP7_75t_L g1226 ( .A(n_434), .B(n_493), .Y(n_1226) );
OR2x6_ASAP7_75t_L g1241 ( .A(n_434), .B(n_739), .Y(n_1241) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx3_ASAP7_75t_L g484 ( .A(n_435), .Y(n_484) );
NAND2xp33_ASAP7_75t_SL g717 ( .A(n_435), .B(n_437), .Y(n_717) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g483 ( .A(n_437), .B(n_484), .Y(n_483) );
AND3x4_ASAP7_75t_L g623 ( .A(n_437), .B(n_484), .C(n_509), .Y(n_623) );
HB1xp67_ASAP7_75t_L g1245 ( .A(n_437), .Y(n_1245) );
AOI222xp33_ASAP7_75t_L g519 ( .A1(n_438), .A2(n_520), .B1(n_530), .B2(n_538), .C1(n_539), .C2(n_544), .Y(n_519) );
INVx4_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_441), .A2(n_446), .B1(n_727), .B2(n_728), .C(n_729), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_441), .A2(n_446), .B1(n_802), .B2(n_803), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g1558 ( .A1(n_441), .A2(n_446), .B1(n_1559), .B2(n_1560), .Y(n_1558) );
AND2x2_ASAP7_75t_L g606 ( .A(n_442), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_SL g1496 ( .A(n_442), .B(n_607), .Y(n_1496) );
NAND2x1_ASAP7_75t_L g1516 ( .A(n_442), .B(n_607), .Y(n_1516) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_442), .B(n_607), .Y(n_1600) );
INVx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_444), .B(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g466 ( .A(n_444), .B(n_448), .Y(n_466) );
BUFx2_ASAP7_75t_L g1231 ( .A(n_444), .Y(n_1231) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_446), .Y(n_1025) );
INVx1_ASAP7_75t_L g611 ( .A(n_447), .Y(n_611) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g454 ( .A(n_450), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g729 ( .A(n_451), .Y(n_729) );
OR2x6_ASAP7_75t_L g451 ( .A(n_452), .B(n_455), .Y(n_451) );
INVx1_ASAP7_75t_L g500 ( .A(n_452), .Y(n_500) );
INVx1_ASAP7_75t_L g1065 ( .A(n_452), .Y(n_1065) );
INVx1_ASAP7_75t_L g1311 ( .A(n_452), .Y(n_1311) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_453), .Y(n_478) );
BUFx3_ASAP7_75t_L g815 ( .A(n_453), .Y(n_815) );
BUFx2_ASAP7_75t_L g1234 ( .A(n_454), .Y(n_1234) );
INVx1_ASAP7_75t_L g944 ( .A(n_455), .Y(n_944) );
OR2x6_ASAP7_75t_SL g457 ( .A(n_458), .B(n_461), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g465 ( .A(n_459), .B(n_466), .Y(n_465) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_459), .Y(n_733) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g490 ( .A(n_460), .Y(n_490) );
OR2x2_ASAP7_75t_L g617 ( .A(n_460), .B(n_586), .Y(n_617) );
INVx3_ASAP7_75t_L g901 ( .A(n_461), .Y(n_901) );
BUFx2_ASAP7_75t_L g1113 ( .A(n_461), .Y(n_1113) );
BUFx2_ASAP7_75t_L g1667 ( .A(n_461), .Y(n_1667) );
INVx1_ASAP7_75t_L g1945 ( .A(n_461), .Y(n_1945) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_462), .Y(n_473) );
BUFx8_ASAP7_75t_L g620 ( .A(n_462), .Y(n_620) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_462), .Y(n_715) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_465), .B(n_746), .Y(n_855) );
BUFx3_ASAP7_75t_L g486 ( .A(n_466), .Y(n_486) );
BUFx12f_ASAP7_75t_L g503 ( .A(n_466), .Y(n_503) );
INVx5_ASAP7_75t_L g630 ( .A(n_466), .Y(n_630) );
BUFx2_ASAP7_75t_L g710 ( .A(n_466), .Y(n_710) );
BUFx3_ASAP7_75t_L g935 ( .A(n_466), .Y(n_935) );
NOR3xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_487), .C(n_494), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_474), .C(n_485), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_470), .B(n_551), .Y(n_562) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g968 ( .A(n_473), .Y(n_968) );
INVx2_ASAP7_75t_L g1036 ( .A(n_473), .Y(n_1036) );
INVx1_ASAP7_75t_L g1055 ( .A(n_473), .Y(n_1055) );
INVx2_ASAP7_75t_L g1162 ( .A(n_473), .Y(n_1162) );
AND2x4_ASAP7_75t_L g1222 ( .A(n_473), .B(n_1223), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g649 ( .A(n_478), .B(n_617), .Y(n_649) );
INVx3_ASAP7_75t_L g808 ( .A(n_478), .Y(n_808) );
BUFx6f_ASAP7_75t_L g914 ( .A(n_478), .Y(n_914) );
INVx4_ASAP7_75t_L g955 ( .A(n_478), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_480), .A2(n_712), .B1(n_794), .B2(n_800), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g906 ( .A1(n_480), .A2(n_607), .B(n_871), .C(n_907), .Y(n_906) );
INVx8_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g615 ( .A(n_481), .Y(n_615) );
INVx2_ASAP7_75t_L g625 ( .A(n_481), .Y(n_625) );
INVx3_ASAP7_75t_L g942 ( .A(n_481), .Y(n_942) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI221xp5_ASAP7_75t_L g964 ( .A1(n_483), .A2(n_965), .B1(n_966), .B2(n_967), .C(n_969), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g1058 ( .A1(n_483), .A2(n_630), .B1(n_708), .B2(n_1059), .C(n_1060), .Y(n_1058) );
OAI221xp5_ASAP7_75t_L g1376 ( .A1(n_483), .A2(n_714), .B1(n_815), .B2(n_1377), .C(n_1378), .Y(n_1376) );
OAI221xp5_ASAP7_75t_L g1452 ( .A1(n_483), .A2(n_1381), .B1(n_1434), .B2(n_1449), .C(n_1453), .Y(n_1452) );
OAI221xp5_ASAP7_75t_L g1562 ( .A1(n_483), .A2(n_914), .B1(n_1033), .B2(n_1563), .C(n_1564), .Y(n_1562) );
INVx3_ASAP7_75t_L g1230 ( .A(n_484), .Y(n_1230) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g1554 ( .A1(n_489), .A2(n_492), .B1(n_1555), .B2(n_1556), .Y(n_1554) );
AND2x2_ASAP7_75t_L g492 ( .A(n_490), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g627 ( .A(n_493), .Y(n_627) );
BUFx2_ASAP7_75t_L g640 ( .A(n_493), .Y(n_640) );
BUFx2_ASAP7_75t_L g712 ( .A(n_493), .Y(n_712) );
BUFx3_ASAP7_75t_L g722 ( .A(n_493), .Y(n_722) );
BUFx2_ASAP7_75t_L g743 ( .A(n_493), .Y(n_743) );
BUFx2_ASAP7_75t_L g1295 ( .A(n_493), .Y(n_1295) );
BUFx2_ASAP7_75t_L g1956 ( .A(n_493), .Y(n_1956) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI22xp33_ASAP7_75t_L g1343 ( .A1(n_496), .A2(n_1323), .B1(n_1333), .B2(n_1344), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1947 ( .A1(n_496), .A2(n_1173), .B1(n_1948), .B2(n_1949), .Y(n_1947) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g1569 ( .A1(n_498), .A2(n_504), .B1(n_966), .B2(n_1570), .C(n_1571), .Y(n_1569) );
BUFx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx4f_ASAP7_75t_L g819 ( .A(n_499), .Y(n_819) );
BUFx3_ASAP7_75t_L g956 ( .A(n_499), .Y(n_956) );
INVx2_ASAP7_75t_L g962 ( .A(n_499), .Y(n_962) );
OR2x4_ASAP7_75t_L g1239 ( .A(n_499), .B(n_1223), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
BUFx2_ASAP7_75t_L g1122 ( .A(n_503), .Y(n_1122) );
INVx3_ASAP7_75t_L g725 ( .A(n_504), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g812 ( .A1(n_504), .A2(n_813), .B1(n_816), .B2(n_817), .C(n_820), .Y(n_812) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_504), .A2(n_953), .B1(n_954), .B2(n_956), .C(n_957), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_504), .B(n_1067), .Y(n_1066) );
OAI221xp5_ASAP7_75t_L g1382 ( .A1(n_504), .A2(n_815), .B1(n_819), .B2(n_1383), .C(n_1384), .Y(n_1382) );
OAI221xp5_ASAP7_75t_L g1447 ( .A1(n_504), .A2(n_817), .B1(n_1448), .B2(n_1449), .C(n_1450), .Y(n_1447) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g927 ( .A(n_505), .B(n_559), .Y(n_927) );
OR2x6_ASAP7_75t_L g1608 ( .A(n_505), .B(n_559), .Y(n_1608) );
OAI21xp33_ASAP7_75t_L g1462 ( .A1(n_507), .A2(n_1463), .B(n_1472), .Y(n_1462) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g699 ( .A(n_508), .Y(n_699) );
BUFx2_ASAP7_75t_L g1653 ( .A(n_508), .Y(n_1653) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_509), .A2(n_1021), .B1(n_1040), .B2(n_1042), .Y(n_1020) );
INVx2_ASAP7_75t_SL g1068 ( .A(n_509), .Y(n_1068) );
OAI31xp33_ASAP7_75t_SL g1552 ( .A1(n_509), .A2(n_1553), .A3(n_1557), .B(n_1561), .Y(n_1552) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_510), .B(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g559 ( .A(n_510), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_513), .Y(n_757) );
INVx1_ASAP7_75t_L g1041 ( .A(n_513), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_513), .B(n_1070), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1579 ( .A(n_513), .B(n_1580), .Y(n_1579) );
INVx2_ASAP7_75t_L g565 ( .A(n_515), .Y(n_565) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_515), .Y(n_694) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx3_ASAP7_75t_L g578 ( .A(n_516), .Y(n_578) );
INVx2_ASAP7_75t_L g761 ( .A(n_516), .Y(n_761) );
AND2x4_ASAP7_75t_L g1214 ( .A(n_516), .B(n_1207), .Y(n_1214) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_545), .C(n_588), .Y(n_518) );
INVxp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVxp67_ASAP7_75t_L g753 ( .A(n_522), .Y(n_753) );
INVx1_ASAP7_75t_L g793 ( .A(n_522), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_522), .A2(n_1003), .B1(n_1004), .B2(n_1005), .Y(n_1002) );
AOI222xp33_ASAP7_75t_L g1392 ( .A1(n_522), .A2(n_530), .B1(n_539), .B2(n_1386), .C1(n_1393), .C2(n_1394), .Y(n_1392) );
AOI222xp33_ASAP7_75t_L g1437 ( .A1(n_522), .A2(n_589), .B1(n_1005), .B2(n_1438), .C1(n_1439), .C2(n_1440), .Y(n_1437) );
AOI21xp33_ASAP7_75t_L g1581 ( .A1(n_522), .A2(n_1582), .B(n_1583), .Y(n_1581) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_526), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OR2x2_ASAP7_75t_L g552 ( .A(n_524), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g754 ( .A(n_524), .B(n_553), .Y(n_754) );
INVx1_ASAP7_75t_L g591 ( .A(n_525), .Y(n_591) );
INVx1_ASAP7_75t_L g637 ( .A(n_525), .Y(n_637) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g1480 ( .A(n_527), .Y(n_1480) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx3_ASAP7_75t_L g580 ( .A(n_528), .Y(n_580) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_528), .Y(n_657) );
BUFx3_ASAP7_75t_L g780 ( .A(n_528), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g851 ( .A1(n_530), .A2(n_539), .B1(n_800), .B2(n_802), .Y(n_851) );
AOI22xp33_ASAP7_75t_SL g1010 ( .A1(n_530), .A2(n_539), .B1(n_1011), .B2(n_1012), .Y(n_1010) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_530), .A2(n_539), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_SL g987 ( .A(n_531), .Y(n_987) );
NAND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_535), .Y(n_531) );
INVx1_ASAP7_75t_L g598 ( .A(n_532), .Y(n_598) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_534), .B(n_542), .Y(n_541) );
AND2x6_ASAP7_75t_L g669 ( .A(n_534), .B(n_548), .Y(n_669) );
INVx1_ASAP7_75t_L g684 ( .A(n_534), .Y(n_684) );
AND2x2_ASAP7_75t_L g879 ( .A(n_534), .B(n_880), .Y(n_879) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g683 ( .A(n_537), .Y(n_683) );
BUFx2_ASAP7_75t_L g880 ( .A(n_537), .Y(n_880) );
AND2x4_ASAP7_75t_L g1198 ( .A(n_537), .B(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g648 ( .A(n_540), .B(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_L g1502 ( .A(n_540), .B(n_649), .Y(n_1502) );
INVx1_ASAP7_75t_L g882 ( .A(n_541), .Y(n_882) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_561), .B1(n_575), .B2(n_579), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_547), .A2(n_580), .B1(n_871), .B2(n_872), .Y(n_870) );
A2O1A1Ixp33_ASAP7_75t_L g875 ( .A1(n_547), .A2(n_848), .B(n_876), .C(n_877), .Y(n_875) );
BUFx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx3_ASAP7_75t_L g576 ( .A(n_548), .Y(n_576) );
BUFx3_ASAP7_75t_L g762 ( .A(n_548), .Y(n_762) );
BUFx6f_ASAP7_75t_L g1089 ( .A(n_548), .Y(n_1089) );
BUFx3_ASAP7_75t_L g1141 ( .A(n_548), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_548), .B(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1399 ( .A(n_548), .Y(n_1399) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g664 ( .A(n_549), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_550), .A2(n_562), .B1(n_563), .B2(n_566), .Y(n_561) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g1005 ( .A(n_552), .Y(n_1005) );
BUFx3_ASAP7_75t_L g978 ( .A(n_553), .Y(n_978) );
INVx2_ASAP7_75t_SL g1255 ( .A(n_553), .Y(n_1255) );
BUFx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_554), .Y(n_597) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g832 ( .A(n_557), .Y(n_832) );
INVx4_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g782 ( .A(n_558), .Y(n_782) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_558), .Y(n_973) );
AOI31xp33_ASAP7_75t_L g1007 ( .A1(n_558), .A2(n_595), .A3(n_1008), .B(n_1009), .Y(n_1007) );
INVx2_ASAP7_75t_L g1085 ( .A(n_558), .Y(n_1085) );
AOI222xp33_ASAP7_75t_L g1395 ( .A1(n_558), .A2(n_589), .B1(n_767), .B2(n_1396), .C1(n_1397), .C2(n_1405), .Y(n_1395) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g746 ( .A(n_559), .Y(n_746) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g666 ( .A(n_564), .Y(n_666) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_569), .B2(n_570), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_568), .A2(n_570), .B1(n_1060), .B2(n_1083), .Y(n_1082) );
OAI22xp33_ASAP7_75t_L g1322 ( .A1(n_570), .A2(n_1323), .B1(n_1324), .B2(n_1328), .Y(n_1322) );
INVx5_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx6_ASAP7_75t_L g690 ( .A(n_571), .Y(n_690) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g1093 ( .A(n_572), .Y(n_1093) );
INVx4_ASAP7_75t_L g1180 ( .A(n_572), .Y(n_1180) );
INVx2_ASAP7_75t_L g1267 ( .A(n_572), .Y(n_1267) );
INVx1_ASAP7_75t_L g1339 ( .A(n_572), .Y(n_1339) );
INVx2_ASAP7_75t_SL g1409 ( .A(n_572), .Y(n_1409) );
INVx1_ASAP7_75t_L g1650 ( .A(n_572), .Y(n_1650) );
INVx8_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_573), .B(n_1199), .Y(n_1210) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g1401 ( .A(n_578), .Y(n_1401) );
BUFx3_ASAP7_75t_L g1135 ( .A(n_580), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1274 ( .A(n_580), .Y(n_1274) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g839 ( .A(n_582), .Y(n_839) );
INVx2_ASAP7_75t_L g984 ( .A(n_582), .Y(n_984) );
INVx2_ASAP7_75t_L g1134 ( .A(n_582), .Y(n_1134) );
INVx1_ASAP7_75t_L g1139 ( .A(n_582), .Y(n_1139) );
INVx1_ASAP7_75t_L g1479 ( .A(n_582), .Y(n_1479) );
INVx1_ASAP7_75t_L g1186 ( .A(n_583), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_587), .Y(n_583) );
AND2x4_ASAP7_75t_L g767 ( .A(n_584), .B(n_587), .Y(n_767) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g910 ( .A(n_586), .B(n_717), .Y(n_910) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_586), .Y(n_1247) );
INVx4_ASAP7_75t_L g667 ( .A(n_587), .Y(n_667) );
INVx4_ASAP7_75t_L g892 ( .A(n_587), .Y(n_892) );
INVx1_ASAP7_75t_SL g1619 ( .A(n_587), .Y(n_1619) );
AOI21xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_594), .B(n_595), .Y(n_588) );
AOI322xp5_ASAP7_75t_L g1079 ( .A1(n_589), .A2(n_767), .A3(n_1080), .B1(n_1081), .B2(n_1084), .C1(n_1086), .C2(n_1087), .Y(n_1079) );
AOI332xp33_ASAP7_75t_L g1584 ( .A1(n_589), .A2(n_767), .A3(n_832), .B1(n_1585), .B2(n_1586), .B3(n_1587), .C1(n_1588), .C2(n_1589), .Y(n_1584) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g647 ( .A(n_591), .B(n_593), .Y(n_647) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g1412 ( .A1(n_595), .A2(n_1005), .B(n_1413), .Y(n_1412) );
NOR3xp33_ASAP7_75t_L g1422 ( .A(n_595), .B(n_1423), .C(n_1424), .Y(n_1422) );
AOI21xp5_ASAP7_75t_L g1578 ( .A1(n_595), .A2(n_1005), .B(n_1560), .Y(n_1578) );
CKINVDCx5p33_ASAP7_75t_R g595 ( .A(n_596), .Y(n_595) );
OAI21xp5_ASAP7_75t_L g768 ( .A1(n_596), .A2(n_769), .B(n_781), .Y(n_768) );
OAI21xp5_ASAP7_75t_SL g829 ( .A1(n_596), .A2(n_830), .B(n_833), .Y(n_829) );
OAI21xp5_ASAP7_75t_L g979 ( .A1(n_596), .A2(n_850), .B(n_980), .Y(n_979) );
OR2x6_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx4_ASAP7_75t_L g776 ( .A(n_597), .Y(n_776) );
BUFx4f_ASAP7_75t_L g837 ( .A(n_597), .Y(n_837) );
BUFx4f_ASAP7_75t_L g846 ( .A(n_597), .Y(n_846) );
BUFx6f_ASAP7_75t_L g1192 ( .A(n_597), .Y(n_1192) );
BUFx4f_ASAP7_75t_L g1476 ( .A(n_597), .Y(n_1476) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_653), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_641), .C(n_652), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_612), .C(n_621), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_608), .B2(n_609), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_606), .A2(n_609), .B1(n_1107), .B2(n_1108), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_606), .A2(n_609), .B1(n_1284), .B2(n_1285), .Y(n_1283) );
AOI22xp33_ASAP7_75t_L g1659 ( .A1(n_606), .A2(n_609), .B1(n_1660), .B2(n_1661), .Y(n_1659) );
AND2x4_ASAP7_75t_L g609 ( .A(n_607), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g652 ( .A(n_607), .B(n_640), .Y(n_652) );
AND2x4_ASAP7_75t_SL g1498 ( .A(n_607), .B(n_610), .Y(n_1498) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_609), .A2(n_1514), .B1(n_1515), .B2(n_1517), .Y(n_1513) );
AOI22xp33_ASAP7_75t_L g1598 ( .A1(n_609), .A2(n_1599), .B1(n_1600), .B2(n_1601), .Y(n_1598) );
AOI22xp33_ASAP7_75t_L g1897 ( .A1(n_609), .A2(n_1515), .B1(n_1898), .B2(n_1899), .Y(n_1897) );
INVx1_ASAP7_75t_L g1940 ( .A(n_609), .Y(n_1940) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B1(n_618), .B2(n_619), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_613), .A2(n_618), .B1(n_671), .B2(n_673), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_614), .B(n_897), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_614), .A2(n_619), .B1(n_1126), .B2(n_1129), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_614), .A2(n_619), .B1(n_1276), .B2(n_1277), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1541 ( .A1(n_614), .A2(n_619), .B1(n_1528), .B2(n_1529), .Y(n_1541) );
AND2x4_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x4_ASAP7_75t_L g1504 ( .A(n_615), .B(n_616), .Y(n_1504) );
AND2x4_ASAP7_75t_L g619 ( .A(n_616), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g643 ( .A(n_617), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g902 ( .A(n_617), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_619), .A2(n_1467), .B1(n_1468), .B2(n_1504), .Y(n_1503) );
INVx2_ASAP7_75t_L g1613 ( .A(n_619), .Y(n_1613) );
INVx2_ASAP7_75t_L g1908 ( .A(n_619), .Y(n_1908) );
INVx3_ASAP7_75t_L g633 ( .A(n_620), .Y(n_633) );
INVx2_ASAP7_75t_SL g822 ( .A(n_620), .Y(n_822) );
INVx3_ASAP7_75t_L g1033 ( .A(n_620), .Y(n_1033) );
HB1xp67_ASAP7_75t_L g1293 ( .A(n_620), .Y(n_1293) );
INVx2_ASAP7_75t_SL g1381 ( .A(n_620), .Y(n_1381) );
AOI33xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .A3(n_628), .B1(n_631), .B2(n_635), .B3(n_638), .Y(n_621) );
INVx1_ASAP7_75t_L g1120 ( .A(n_622), .Y(n_1120) );
AOI33xp33_ASAP7_75t_L g1289 ( .A1(n_622), .A2(n_1170), .A3(n_1290), .B1(n_1291), .B2(n_1292), .B3(n_1294), .Y(n_1289) );
AOI33xp33_ASAP7_75t_L g1518 ( .A1(n_622), .A2(n_1170), .A3(n_1519), .B1(n_1522), .B2(n_1523), .B3(n_1524), .Y(n_1518) );
AOI33xp33_ASAP7_75t_L g1662 ( .A1(n_622), .A2(n_635), .A3(n_1663), .B1(n_1665), .B2(n_1668), .B3(n_1669), .Y(n_1662) );
BUFx3_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI33xp33_ASAP7_75t_L g1602 ( .A1(n_623), .A2(n_1603), .A3(n_1604), .B1(n_1605), .B2(n_1607), .B3(n_1609), .Y(n_1602) );
AOI33xp33_ASAP7_75t_L g1900 ( .A1(n_623), .A2(n_1901), .A3(n_1902), .B1(n_1904), .B2(n_1905), .B3(n_1906), .Y(n_1900) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_625), .A2(n_741), .B1(n_742), .B2(n_743), .Y(n_740) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g937 ( .A(n_627), .Y(n_937) );
INVx2_ASAP7_75t_L g1114 ( .A(n_627), .Y(n_1114) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g634 ( .A(n_630), .Y(n_634) );
INVx2_ASAP7_75t_R g1606 ( .A(n_630), .Y(n_1606) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g1348 ( .A(n_635), .Y(n_1348) );
CKINVDCx5p33_ASAP7_75t_R g1493 ( .A(n_635), .Y(n_1493) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx3_ASAP7_75t_L g1117 ( .A(n_636), .Y(n_1117) );
BUFx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_640), .A2(n_942), .B1(n_999), .B2(n_1012), .Y(n_1037) );
INVx8_ASAP7_75t_L g1103 ( .A(n_642), .Y(n_1103) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_647), .Y(n_642) );
BUFx3_ASAP7_75t_L g1167 ( .A(n_644), .Y(n_1167) );
INVx1_ASAP7_75t_L g1576 ( .A(n_644), .Y(n_1576) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_645), .Y(n_825) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx2_ASAP7_75t_L g739 ( .A(n_646), .Y(n_739) );
INVx1_ASAP7_75t_L g752 ( .A(n_647), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_647), .B(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g903 ( .A(n_649), .Y(n_903) );
INVx3_ASAP7_75t_L g1101 ( .A(n_650), .Y(n_1101) );
INVx5_ASAP7_75t_L g1288 ( .A(n_650), .Y(n_1288) );
INVx3_ASAP7_75t_L g1109 ( .A(n_652), .Y(n_1109) );
INVx3_ASAP7_75t_L g1296 ( .A(n_652), .Y(n_1296) );
NOR3xp33_ASAP7_75t_L g1481 ( .A(n_652), .B(n_1482), .C(n_1494), .Y(n_1481) );
NOR3xp33_ASAP7_75t_L g1596 ( .A(n_652), .B(n_1597), .C(n_1610), .Y(n_1596) );
OAI21xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_676), .B(n_697), .Y(n_653) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_656), .A2(n_669), .B1(n_1102), .B2(n_1132), .C(n_1133), .Y(n_1131) );
AOI221xp5_ASAP7_75t_L g1530 ( .A1(n_656), .A2(n_669), .B1(n_1510), .B2(n_1531), .C(n_1535), .Y(n_1530) );
INVx2_ASAP7_75t_SL g1616 ( .A(n_656), .Y(n_1616) );
BUFx2_ASAP7_75t_L g840 ( .A(n_657), .Y(n_840) );
INVx1_ASAP7_75t_L g1016 ( .A(n_657), .Y(n_1016) );
HB1xp67_ASAP7_75t_L g1621 ( .A(n_657), .Y(n_1621) );
AOI21xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_668), .B(n_669), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g1019 ( .A(n_663), .Y(n_1019) );
BUFx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g1534 ( .A(n_664), .Y(n_1534) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
HB1xp67_ASAP7_75t_SL g1641 ( .A(n_667), .Y(n_1641) );
AOI21xp5_ASAP7_75t_L g1271 ( .A1(n_669), .A2(n_1272), .B(n_1273), .Y(n_1271) );
AOI21xp5_ASAP7_75t_L g1469 ( .A1(n_669), .A2(n_1470), .B(n_1471), .Y(n_1469) );
AOI21xp5_ASAP7_75t_L g1617 ( .A1(n_669), .A2(n_1618), .B(n_1620), .Y(n_1617) );
AOI21xp5_ASAP7_75t_L g1637 ( .A1(n_669), .A2(n_1638), .B(n_1642), .Y(n_1637) );
AOI21xp5_ASAP7_75t_SL g1914 ( .A1(n_669), .A2(n_1915), .B(n_1916), .Y(n_1914) );
INVx1_ASAP7_75t_L g1965 ( .A(n_669), .Y(n_1965) );
AOI22xp33_ASAP7_75t_L g1917 ( .A1(n_671), .A2(n_1130), .B1(n_1918), .B2(n_1919), .Y(n_1917) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g1644 ( .A1(n_673), .A2(n_1127), .B1(n_1645), .B2(n_1646), .Y(n_1644) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx6f_ASAP7_75t_L g1130 ( .A(n_675), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_675), .A2(n_1128), .B1(n_1467), .B2(n_1468), .Y(n_1466) );
AOI22xp33_ASAP7_75t_L g1622 ( .A1(n_675), .A2(n_1128), .B1(n_1623), .B2(n_1624), .Y(n_1622) );
HB1xp67_ASAP7_75t_L g1968 ( .A(n_675), .Y(n_1968) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g1252 ( .A(n_678), .Y(n_1252) );
INVx2_ASAP7_75t_L g1473 ( .A(n_678), .Y(n_1473) );
INVx4_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
BUFx3_ASAP7_75t_L g1137 ( .A(n_680), .Y(n_1137) );
BUFx2_ASAP7_75t_L g1626 ( .A(n_681), .Y(n_1626) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g1269 ( .A(n_682), .Y(n_1269) );
NOR2x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g877 ( .A(n_684), .Y(n_877) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_689), .B1(n_690), .B2(n_691), .C(n_692), .Y(n_685) );
OAI221xp5_ASAP7_75t_L g1648 ( .A1(n_686), .A2(n_1649), .B1(n_1650), .B2(n_1651), .C(n_1652), .Y(n_1648) );
OAI221xp5_ASAP7_75t_L g1921 ( .A1(n_686), .A2(n_1266), .B1(n_1922), .B2(n_1923), .C(n_1924), .Y(n_1921) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_SL g1336 ( .A(n_687), .Y(n_1336) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx3_ASAP7_75t_L g765 ( .A(n_688), .Y(n_765) );
INVx4_ASAP7_75t_L g1404 ( .A(n_688), .Y(n_1404) );
OAI22xp33_ASAP7_75t_L g763 ( .A1(n_690), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_763) );
OAI221xp5_ASAP7_75t_L g980 ( .A1(n_690), .A2(n_950), .B1(n_965), .B2(n_981), .C(n_983), .Y(n_980) );
BUFx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx3_ASAP7_75t_L g889 ( .A(n_696), .Y(n_889) );
INVx1_ASAP7_75t_L g1142 ( .A(n_696), .Y(n_1142) );
INVx2_ASAP7_75t_L g1260 ( .A(n_696), .Y(n_1260) );
A2O1A1Ixp33_ASAP7_75t_SL g1441 ( .A1(n_697), .A2(n_1442), .B(n_1445), .C(n_1455), .Y(n_1441) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g827 ( .A(n_699), .Y(n_827) );
INVx2_ASAP7_75t_SL g857 ( .A(n_700), .Y(n_857) );
XNOR2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_786), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_784), .B(n_785), .Y(n_701) );
AND3x1_ASAP7_75t_L g702 ( .A(n_703), .B(n_749), .C(n_758), .Y(n_702) );
AOI31xp33_ASAP7_75t_L g785 ( .A1(n_703), .A2(n_749), .A3(n_758), .B(n_784), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_745), .B(n_747), .Y(n_703) );
NAND3xp33_ASAP7_75t_SL g704 ( .A(n_705), .B(n_726), .C(n_730), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_711), .B1(n_718), .B2(n_721), .Y(n_705) );
BUFx2_ASAP7_75t_SL g1664 ( .A(n_707), .Y(n_1664) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g1521 ( .A(n_709), .Y(n_1521) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_714), .A2(n_1330), .B1(n_1337), .B2(n_1346), .Y(n_1345) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_SL g720 ( .A(n_715), .Y(n_720) );
INVx3_ASAP7_75t_L g735 ( .A(n_715), .Y(n_735) );
INVx5_ASAP7_75t_L g917 ( .A(n_715), .Y(n_917) );
HB1xp67_ASAP7_75t_L g949 ( .A(n_715), .Y(n_949) );
BUFx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
BUFx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g1022 ( .A(n_729), .B(n_1023), .Y(n_1022) );
INVxp67_ASAP7_75t_L g798 ( .A(n_731), .Y(n_798) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g933 ( .A(n_733), .Y(n_933) );
INVx2_ASAP7_75t_L g1953 ( .A(n_735), .Y(n_1953) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_736), .A2(n_959), .B1(n_960), .B2(n_963), .Y(n_958) );
OAI21xp33_ASAP7_75t_L g1487 ( .A1(n_736), .A2(n_1488), .B(n_1489), .Y(n_1487) );
INVx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g918 ( .A(n_738), .Y(n_918) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
BUFx3_ASAP7_75t_L g951 ( .A(n_739), .Y(n_951) );
INVx2_ASAP7_75t_L g1145 ( .A(n_745), .Y(n_1145) );
INVx1_ASAP7_75t_L g1539 ( .A(n_745), .Y(n_1539) );
BUFx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI21xp5_ASAP7_75t_SL g866 ( .A1(n_746), .A2(n_867), .B(n_884), .Y(n_866) );
INVx1_ASAP7_75t_L g971 ( .A(n_746), .Y(n_971) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_755), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_757), .B(n_1456), .Y(n_1455) );
AOI211xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_767), .B(n_768), .C(n_783), .Y(n_758) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g888 ( .A(n_761), .Y(n_888) );
INVx2_ASAP7_75t_SL g1971 ( .A(n_765), .Y(n_1971) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_767), .Y(n_850) );
NAND3xp33_ASAP7_75t_L g1013 ( .A(n_767), .B(n_1014), .C(n_1017), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_774), .B1(n_775), .B2(n_777), .C(n_778), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_770), .A2(n_846), .B1(n_1159), .B2(n_1174), .Y(n_1184) );
OAI221xp5_ASAP7_75t_L g1432 ( .A1(n_770), .A2(n_837), .B1(n_1433), .B2(n_1434), .C(n_1435), .Y(n_1432) );
INVx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
BUFx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx2_ASAP7_75t_L g835 ( .A(n_773), .Y(n_835) );
BUFx2_ASAP7_75t_L g845 ( .A(n_773), .Y(n_845) );
INVx1_ASAP7_75t_L g982 ( .A(n_773), .Y(n_982) );
INVx1_ASAP7_75t_L g1429 ( .A(n_775), .Y(n_1429) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g1183 ( .A(n_776), .Y(n_1183) );
INVx3_ASAP7_75t_L g849 ( .A(n_779), .Y(n_849) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_779), .Y(n_894) );
OAI33xp33_ASAP7_75t_L g1321 ( .A1(n_781), .A2(n_1185), .A3(n_1322), .B1(n_1329), .B2(n_1332), .B3(n_1335), .Y(n_1321) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND3xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_796), .C(n_828), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
OAI21xp33_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_811), .B(n_827), .Y(n_796) );
OAI211xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B(n_801), .C(n_804), .Y(n_797) );
OAI211xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B(n_809), .C(n_810), .Y(n_804) );
OAI221xp5_ASAP7_75t_L g842 ( .A1(n_805), .A2(n_816), .B1(n_843), .B2(n_846), .C(n_847), .Y(n_842) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g1351 ( .A(n_808), .Y(n_1351) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g924 ( .A1(n_815), .A2(n_819), .B1(n_925), .B2(n_926), .Y(n_924) );
BUFx6f_ASAP7_75t_L g1173 ( .A(n_815), .Y(n_1173) );
OAI22xp33_ASAP7_75t_L g1157 ( .A1(n_817), .A2(n_914), .B1(n_1158), .B2(n_1159), .Y(n_1157) );
OAI22xp33_ASAP7_75t_L g1171 ( .A1(n_817), .A2(n_1172), .B1(n_1173), .B2(n_1174), .Y(n_1171) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OAI22xp33_ASAP7_75t_L g911 ( .A1(n_819), .A2(n_912), .B1(n_913), .B2(n_914), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_823), .B1(n_824), .B2(n_826), .Y(n_821) );
OAI221xp5_ASAP7_75t_L g833 ( .A1(n_823), .A2(n_834), .B1(n_836), .B2(n_837), .C(n_838), .Y(n_833) );
OAI221xp5_ASAP7_75t_L g1490 ( .A1(n_824), .A2(n_967), .B1(n_1475), .B2(n_1491), .C(n_1492), .Y(n_1490) );
CKINVDCx8_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
INVx3_ASAP7_75t_L g1164 ( .A(n_825), .Y(n_1164) );
INVx3_ASAP7_75t_L g1346 ( .A(n_825), .Y(n_1346) );
INVx3_ASAP7_75t_L g1568 ( .A(n_825), .Y(n_1568) );
INVx1_ASAP7_75t_L g1631 ( .A(n_827), .Y(n_1631) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_841), .C(n_852), .Y(n_828) );
INVxp67_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g1181 ( .A1(n_834), .A2(n_1161), .B1(n_1166), .B2(n_1182), .Y(n_1181) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx2_ASAP7_75t_L g1257 ( .A(n_835), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_843), .A2(n_1192), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_843), .A2(n_1254), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g869 ( .A(n_844), .Y(n_869) );
INVx4_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
XNOR2xp5_ASAP7_75t_L g859 ( .A(n_860), .B(n_993), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
XNOR2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_928), .Y(n_861) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
OR2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_895), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_873), .B(n_874), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_878), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_879), .A2(n_881), .B1(n_882), .B2(n_883), .Y(n_878) );
INVx1_ASAP7_75t_L g1144 ( .A(n_879), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_883), .A2(n_899), .B1(n_900), .B2(n_903), .Y(n_898) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_890), .B1(n_891), .B2(n_893), .Y(n_884) );
INVx2_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g1018 ( .A(n_887), .Y(n_1018) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
HB1xp67_ASAP7_75t_L g1643 ( .A(n_894), .Y(n_1643) );
NAND3xp33_ASAP7_75t_SL g895 ( .A(n_896), .B(n_898), .C(n_904), .Y(n_895) );
AND2x2_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
INVx2_ASAP7_75t_L g921 ( .A(n_901), .Y(n_921) );
INVxp67_ASAP7_75t_L g1612 ( .A(n_902), .Y(n_1612) );
NOR2xp33_ASAP7_75t_SL g904 ( .A(n_905), .B(n_908), .Y(n_904) );
OAI33xp33_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_911), .A3(n_915), .B1(n_920), .B2(n_924), .B3(n_927), .Y(n_908) );
BUFx3_ASAP7_75t_L g1342 ( .A(n_909), .Y(n_1342) );
BUFx4f_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
BUFx2_ASAP7_75t_L g1156 ( .A(n_910), .Y(n_1156) );
BUFx8_ASAP7_75t_L g1486 ( .A(n_910), .Y(n_1486) );
HB1xp67_ASAP7_75t_L g1344 ( .A(n_914), .Y(n_1344) );
OAI22xp5_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_917), .B1(n_918), .B2(n_919), .Y(n_915) );
INVx8_ASAP7_75t_L g1029 ( .A(n_917), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_918), .A2(n_921), .B1(n_922), .B2(n_923), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_921), .A2(n_951), .B1(n_1331), .B2(n_1340), .Y(n_1347) );
NAND4xp75_ASAP7_75t_L g929 ( .A(n_930), .B(n_972), .C(n_989), .D(n_990), .Y(n_929) );
OAI21x1_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_945), .B(n_970), .Y(n_930) );
OAI21xp5_ASAP7_75t_L g931 ( .A1(n_932), .A2(n_934), .B(n_940), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_933), .A2(n_1003), .B1(n_1035), .B2(n_1038), .Y(n_1034) );
AOI221xp5_ASAP7_75t_SL g934 ( .A1(n_935), .A2(n_936), .B1(n_937), .B2(n_938), .C(n_939), .Y(n_934) );
A2O1A1Ixp33_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_942), .B(n_943), .C(n_944), .Y(n_940) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_952), .B1(n_958), .B2(n_964), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_947), .A2(n_948), .B1(n_950), .B2(n_951), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g975 ( .A1(n_947), .A2(n_959), .B1(n_976), .B2(n_978), .Y(n_975) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g1942 ( .A1(n_951), .A2(n_1943), .B1(n_1944), .B2(n_1946), .Y(n_1942) );
OAI221xp5_ASAP7_75t_L g1950 ( .A1(n_951), .A2(n_1951), .B1(n_1952), .B2(n_1954), .C(n_1955), .Y(n_1950) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g966 ( .A(n_955), .Y(n_966) );
INVx2_ASAP7_75t_L g1057 ( .A(n_955), .Y(n_1057) );
INVx2_ASAP7_75t_L g1449 ( .A(n_955), .Y(n_1449) );
BUFx4f_ASAP7_75t_SL g960 ( .A(n_961), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g1565 ( .A1(n_961), .A2(n_1566), .B1(n_1567), .B2(n_1568), .Y(n_1565) );
INVx3_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx2_ASAP7_75t_SL g1350 ( .A(n_962), .Y(n_1350) );
INVx2_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
AOI211x1_ASAP7_75t_L g972 ( .A1(n_973), .A2(n_974), .B(n_979), .C(n_985), .Y(n_972) );
INVx1_ASAP7_75t_L g1178 ( .A(n_976), .Y(n_1178) );
BUFx3_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
BUFx3_ASAP7_75t_L g1091 ( .A(n_977), .Y(n_1091) );
INVx2_ASAP7_75t_SL g1264 ( .A(n_977), .Y(n_1264) );
BUFx6f_ASAP7_75t_L g1431 ( .A(n_977), .Y(n_1431) );
BUFx2_ASAP7_75t_L g1354 ( .A(n_978), .Y(n_1354) );
INVx2_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_1044), .B1(n_1045), .B2(n_1094), .Y(n_993) );
INVx1_ASAP7_75t_L g1094 ( .A(n_994), .Y(n_1094) );
OAI21x1_ASAP7_75t_SL g994 ( .A1(n_995), .A2(n_996), .B(n_1043), .Y(n_994) );
NAND4xp25_ASAP7_75t_L g1043 ( .A(n_995), .B(n_998), .C(n_1000), .D(n_1020), .Y(n_1043) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
NAND3xp33_ASAP7_75t_L g997 ( .A(n_998), .B(n_1000), .C(n_1020), .Y(n_997) );
NOR2xp33_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1006), .Y(n_1000) );
NAND3xp33_ASAP7_75t_SL g1006 ( .A(n_1007), .B(n_1010), .C(n_1013), .Y(n_1006) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
NAND3xp33_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1026), .C(n_1034), .Y(n_1021) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_1027), .A2(n_1028), .B1(n_1030), .B2(n_1031), .Y(n_1026) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
OAI21xp5_ASAP7_75t_L g1483 ( .A1(n_1033), .A2(n_1484), .B(n_1485), .Y(n_1483) );
OAI22xp5_ASAP7_75t_L g1572 ( .A1(n_1033), .A2(n_1573), .B1(n_1574), .B2(n_1575), .Y(n_1572) );
INVx1_ASAP7_75t_L g1903 ( .A(n_1033), .Y(n_1903) );
INVx1_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_1040), .B(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
NOR2x1_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1071), .Y(n_1046) );
A2O1A1Ixp33_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1052), .B(n_1068), .C(n_1069), .Y(n_1047) );
NOR3xp33_ASAP7_75t_SL g1052 ( .A(n_1053), .B(n_1061), .C(n_1062), .Y(n_1052) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_1059), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1090) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
O2A1O1Ixp5_ASAP7_75t_L g1250 ( .A1(n_1068), .A2(n_1251), .B(n_1270), .C(n_1278), .Y(n_1250) );
OAI21xp5_ASAP7_75t_L g1912 ( .A1(n_1068), .A2(n_1913), .B(n_1920), .Y(n_1912) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1079), .Y(n_1071) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
OAI33xp33_ASAP7_75t_L g1175 ( .A1(n_1085), .A2(n_1176), .A3(n_1181), .B1(n_1184), .B2(n_1185), .B3(n_1187), .Y(n_1175) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1089), .Y(n_1640) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
NAND2xp67_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1123), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1102), .B1(n_1103), .B2(n_1104), .C(n_1105), .Y(n_1100) );
AOI221xp5_ASAP7_75t_L g1509 ( .A1(n_1101), .A2(n_1103), .B1(n_1510), .B2(n_1511), .C(n_1512), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1280 ( .A(n_1103), .B(n_1281), .Y(n_1280) );
AOI21xp5_ASAP7_75t_L g1499 ( .A1(n_1103), .A2(n_1500), .B(n_1501), .Y(n_1499) );
AOI21xp33_ASAP7_75t_L g1593 ( .A1(n_1103), .A2(n_1594), .B(n_1595), .Y(n_1593) );
AOI21xp5_ASAP7_75t_L g1654 ( .A1(n_1103), .A2(n_1655), .B(n_1656), .Y(n_1654) );
AOI21xp33_ASAP7_75t_SL g1909 ( .A1(n_1103), .A2(n_1910), .B(n_1911), .Y(n_1909) );
AOI21xp5_ASAP7_75t_L g1957 ( .A1(n_1103), .A2(n_1958), .B(n_1959), .Y(n_1957) );
NAND3xp33_ASAP7_75t_SL g1105 ( .A(n_1106), .B(n_1109), .C(n_1110), .Y(n_1105) );
AOI222xp33_ASAP7_75t_L g1136 ( .A1(n_1107), .A2(n_1108), .B1(n_1137), .B2(n_1138), .C1(n_1140), .C2(n_1143), .Y(n_1136) );
NAND3xp33_ASAP7_75t_SL g1512 ( .A(n_1109), .B(n_1513), .C(n_1518), .Y(n_1512) );
INVx2_ASAP7_75t_SL g1672 ( .A(n_1109), .Y(n_1672) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_1111), .A2(n_1115), .B1(n_1119), .B2(n_1121), .Y(n_1110) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1165 ( .A1(n_1113), .A2(n_1166), .B1(n_1167), .B2(n_1168), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1116), .B(n_1118), .Y(n_1115) );
BUFx2_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
BUFx2_ASAP7_75t_L g1170 ( .A(n_1117), .Y(n_1170) );
BUFx2_ASAP7_75t_L g1905 ( .A(n_1117), .Y(n_1905) );
AOI21xp5_ASAP7_75t_L g1123 ( .A1(n_1124), .A2(n_1145), .B(n_1146), .Y(n_1123) );
NAND3xp33_ASAP7_75t_SL g1124 ( .A(n_1125), .B(n_1131), .C(n_1136), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1125 ( .A1(n_1126), .A2(n_1127), .B1(n_1129), .B2(n_1130), .Y(n_1125) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_1128), .A2(n_1130), .B1(n_1276), .B2(n_1277), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1527 ( .A1(n_1128), .A2(n_1130), .B1(n_1528), .B2(n_1529), .Y(n_1527) );
INVx1_ASAP7_75t_L g1975 ( .A(n_1128), .Y(n_1975) );
AOI222xp33_ASAP7_75t_L g1536 ( .A1(n_1137), .A2(n_1143), .B1(n_1514), .B2(n_1517), .C1(n_1537), .C2(n_1538), .Y(n_1536) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
A2O1A1Ixp33_ASAP7_75t_L g1372 ( .A1(n_1145), .A2(n_1373), .B(n_1385), .C(n_1389), .Y(n_1372) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
AOI22xp5_ASAP7_75t_L g1149 ( .A1(n_1150), .A2(n_1415), .B1(n_1673), .B2(n_1674), .Y(n_1149) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1150), .Y(n_1673) );
AO22x2_ASAP7_75t_L g1150 ( .A1(n_1151), .A2(n_1297), .B1(n_1298), .B2(n_1414), .Y(n_1150) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1151), .Y(n_1414) );
XNOR2xp5_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1248), .Y(n_1151) );
NAND3xp33_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1190), .C(n_1218), .Y(n_1153) );
NOR2xp33_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1175), .Y(n_1154) );
OAI33xp33_ASAP7_75t_L g1155 ( .A1(n_1156), .A2(n_1157), .A3(n_1160), .B1(n_1165), .B2(n_1169), .B3(n_1171), .Y(n_1155) );
OAI22xp5_ASAP7_75t_SL g1176 ( .A1(n_1158), .A2(n_1172), .B1(n_1177), .B2(n_1179), .Y(n_1176) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_1161), .A2(n_1162), .B1(n_1163), .B2(n_1164), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_1163), .A2(n_1168), .B1(n_1177), .B2(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
OAI211xp5_ASAP7_75t_L g1425 ( .A1(n_1179), .A2(n_1426), .B(n_1427), .C(n_1428), .Y(n_1425) );
HB1xp67_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1180), .Y(n_1189) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_1180), .A2(n_1384), .B1(n_1403), .B2(n_1404), .Y(n_1402) );
HB1xp67_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
OAI211xp5_ASAP7_75t_SL g1627 ( .A1(n_1183), .A2(n_1628), .B(n_1629), .C(n_1630), .Y(n_1627) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
OAI221xp5_ASAP7_75t_L g1962 ( .A1(n_1188), .A2(n_1263), .B1(n_1946), .B2(n_1954), .C(n_1963), .Y(n_1962) );
OAI221xp5_ASAP7_75t_L g1969 ( .A1(n_1188), .A2(n_1948), .B1(n_1970), .B2(n_1972), .C(n_1973), .Y(n_1969) );
INVx2_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
OAI31xp33_ASAP7_75t_L g1190 ( .A1(n_1191), .A2(n_1204), .A3(n_1211), .B(n_1215), .Y(n_1190) );
INVx3_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_1197), .A2(n_1198), .B1(n_1200), .B2(n_1201), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_1197), .A2(n_1228), .B1(n_1232), .B2(n_1235), .Y(n_1227) );
BUFx3_ASAP7_75t_L g1356 ( .A(n_1198), .Y(n_1356) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
INVx2_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx2_ASAP7_75t_L g1359 ( .A(n_1203), .Y(n_1359) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1206), .Y(n_1362) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx2_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
BUFx2_ASAP7_75t_L g1364 ( .A(n_1210), .Y(n_1364) );
INVx3_ASAP7_75t_SL g1213 ( .A(n_1214), .Y(n_1213) );
CKINVDCx16_ASAP7_75t_R g1366 ( .A(n_1214), .Y(n_1366) );
OAI31xp33_ASAP7_75t_L g1352 ( .A1(n_1215), .A2(n_1353), .A3(n_1360), .B(n_1365), .Y(n_1352) );
BUFx3_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
OAI31xp33_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1224), .A3(n_1236), .B(n_1242), .Y(n_1218) );
INVx2_ASAP7_75t_SL g1307 ( .A(n_1220), .Y(n_1307) );
INVx2_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1222), .Y(n_1308) );
CKINVDCx8_ASAP7_75t_R g1225 ( .A(n_1226), .Y(n_1225) );
BUFx3_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
BUFx3_ASAP7_75t_L g1313 ( .A(n_1229), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1230), .B(n_1231), .Y(n_1229) );
AND2x4_ASAP7_75t_L g1233 ( .A(n_1230), .B(n_1234), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_1232), .A2(n_1313), .B1(n_1314), .B2(n_1315), .Y(n_1312) );
BUFx6f_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx2_ASAP7_75t_SL g1238 ( .A(n_1239), .Y(n_1238) );
BUFx2_ASAP7_75t_L g1317 ( .A(n_1239), .Y(n_1317) );
BUFx3_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx2_ASAP7_75t_L g1319 ( .A(n_1241), .Y(n_1319) );
BUFx2_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
AND2x2_ASAP7_75t_SL g1243 ( .A(n_1244), .B(n_1246), .Y(n_1243) );
AND2x4_ASAP7_75t_L g1303 ( .A(n_1244), .B(n_1246), .Y(n_1303) );
INVx1_ASAP7_75t_SL g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
NAND3x1_ASAP7_75t_L g1249 ( .A(n_1250), .B(n_1280), .C(n_1282), .Y(n_1249) );
OAI221xp5_ASAP7_75t_L g1253 ( .A1(n_1254), .A2(n_1256), .B1(n_1257), .B2(n_1258), .C(n_1259), .Y(n_1253) );
INVx5_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1261 ( .A1(n_1262), .A2(n_1263), .B1(n_1265), .B2(n_1268), .Y(n_1261) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
BUFx2_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
BUFx6f_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVxp33_ASAP7_75t_L g1436 ( .A(n_1267), .Y(n_1436) );
AND4x1_ASAP7_75t_SL g1282 ( .A(n_1283), .B(n_1286), .C(n_1289), .D(n_1296), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1288), .Y(n_1286) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
AOI22xp5_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1300), .B1(n_1369), .B2(n_1370), .Y(n_1298) );
INVx2_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1301), .Y(n_1367) );
OAI211xp5_ASAP7_75t_L g1301 ( .A1(n_1302), .A2(n_1304), .B(n_1320), .C(n_1352), .Y(n_1301) );
CKINVDCx14_ASAP7_75t_R g1302 ( .A(n_1303), .Y(n_1302) );
NOR3xp33_ASAP7_75t_SL g1304 ( .A(n_1305), .B(n_1309), .C(n_1316), .Y(n_1304) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_1314), .A2(n_1356), .B1(n_1357), .B2(n_1358), .Y(n_1355) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
NOR2xp33_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1341), .Y(n_1320) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
OAI22xp5_ASAP7_75t_L g1406 ( .A1(n_1326), .A2(n_1407), .B1(n_1408), .B2(n_1409), .Y(n_1406) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_1328), .A2(n_1334), .B1(n_1350), .B2(n_1351), .Y(n_1349) );
OAI22xp5_ASAP7_75t_L g1335 ( .A1(n_1336), .A2(n_1337), .B1(n_1338), .B2(n_1340), .Y(n_1335) );
BUFx3_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
OAI33xp33_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1343), .A3(n_1345), .B1(n_1347), .B2(n_1348), .B3(n_1349), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1611 ( .A(n_1350), .B(n_1612), .Y(n_1611) );
OR2x6_ASAP7_75t_L g1671 ( .A(n_1350), .B(n_1612), .Y(n_1671) );
INVx2_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
HB1xp67_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1391), .Y(n_1371) );
NOR3xp33_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1375), .C(n_1379), .Y(n_1373) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
NAND4xp25_ASAP7_75t_L g1391 ( .A(n_1392), .B(n_1395), .C(n_1410), .D(n_1412), .Y(n_1391) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
INVx1_ASAP7_75t_L g1964 ( .A(n_1399), .Y(n_1964) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1415), .Y(n_1674) );
XNOR2xp5_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1546), .Y(n_1415) );
AOI22xp5_ASAP7_75t_L g1416 ( .A1(n_1417), .A2(n_1458), .B1(n_1543), .B2(n_1545), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
HB1xp67_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1419), .Y(n_1544) );
XOR2x2_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1457), .Y(n_1419) );
NOR2x1_ASAP7_75t_SL g1420 ( .A(n_1421), .B(n_1441), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1432), .Y(n_1424) );
INVx2_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
NOR3xp33_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1451), .C(n_1454), .Y(n_1445) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1458), .Y(n_1545) );
AOI22xp5_ASAP7_75t_L g1458 ( .A1(n_1459), .A2(n_1505), .B1(n_1506), .B2(n_1542), .Y(n_1458) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1459), .Y(n_1542) );
HB1xp67_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
AND4x1_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1481), .C(n_1499), .D(n_1503), .Y(n_1461) );
INVx2_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
OAI211xp5_ASAP7_75t_L g1474 ( .A1(n_1475), .A2(n_1476), .B(n_1477), .C(n_1478), .Y(n_1474) );
OAI22xp5_ASAP7_75t_L g1482 ( .A1(n_1483), .A2(n_1487), .B1(n_1490), .B2(n_1493), .Y(n_1482) );
CKINVDCx20_ASAP7_75t_R g1485 ( .A(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
BUFx3_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1509), .B(n_1525), .Y(n_1508) );
INVx2_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
AOI21xp5_ASAP7_75t_SL g1525 ( .A1(n_1526), .A2(n_1539), .B(n_1540), .Y(n_1525) );
NAND3xp33_ASAP7_75t_SL g1526 ( .A(n_1527), .B(n_1530), .C(n_1536), .Y(n_1526) );
INVx2_ASAP7_75t_L g1532 ( .A(n_1533), .Y(n_1532) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
OAI31xp33_ASAP7_75t_L g1960 ( .A1(n_1539), .A2(n_1961), .A3(n_1966), .B(n_1974), .Y(n_1960) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
XNOR2xp5_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1632), .Y(n_1546) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
XNOR2xp5_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1591), .Y(n_1548) );
XOR2x2_ASAP7_75t_L g1549 ( .A(n_1550), .B(n_1590), .Y(n_1549) );
NOR2xp33_ASAP7_75t_L g1550 ( .A(n_1551), .B(n_1577), .Y(n_1550) );
OAI22xp5_ASAP7_75t_L g1561 ( .A1(n_1562), .A2(n_1565), .B1(n_1569), .B2(n_1572), .Y(n_1561) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
NAND4xp25_ASAP7_75t_SL g1577 ( .A(n_1578), .B(n_1579), .C(n_1581), .D(n_1584), .Y(n_1577) );
NAND3xp33_ASAP7_75t_SL g1592 ( .A(n_1593), .B(n_1596), .C(n_1614), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g1597 ( .A(n_1598), .B(n_1602), .Y(n_1597) );
INVx1_ASAP7_75t_L g1939 ( .A(n_1600), .Y(n_1939) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
OAI21xp5_ASAP7_75t_L g1614 ( .A1(n_1615), .A2(n_1625), .B(n_1631), .Y(n_1614) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1633), .Y(n_1632) );
NAND3xp33_ASAP7_75t_SL g1634 ( .A(n_1635), .B(n_1654), .C(n_1657), .Y(n_1634) );
OAI21xp33_ASAP7_75t_L g1635 ( .A1(n_1636), .A2(n_1647), .B(n_1653), .Y(n_1635) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
NOR3xp33_ASAP7_75t_L g1657 ( .A(n_1658), .B(n_1670), .C(n_1672), .Y(n_1657) );
NAND2xp5_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1662), .Y(n_1658) );
INVx1_ASAP7_75t_L g1666 ( .A(n_1667), .Y(n_1666) );
NOR3xp33_ASAP7_75t_L g1895 ( .A(n_1672), .B(n_1896), .C(n_1907), .Y(n_1895) );
OAI221xp5_ASAP7_75t_L g1675 ( .A1(n_1676), .A2(n_1890), .B1(n_1893), .B2(n_1925), .C(n_1928), .Y(n_1675) );
AOI21xp5_ASAP7_75t_L g1676 ( .A1(n_1677), .A2(n_1816), .B(n_1864), .Y(n_1676) );
NAND5xp2_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1766), .C(n_1782), .D(n_1795), .E(n_1808), .Y(n_1677) );
AOI211xp5_ASAP7_75t_L g1678 ( .A1(n_1679), .A2(n_1710), .B(n_1725), .C(n_1750), .Y(n_1678) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1680), .B(n_1696), .Y(n_1679) );
AND2x2_ASAP7_75t_L g1842 ( .A(n_1680), .B(n_1777), .Y(n_1842) );
CKINVDCx5p33_ASAP7_75t_R g1680 ( .A(n_1681), .Y(n_1680) );
OR2x2_ASAP7_75t_L g1768 ( .A(n_1681), .B(n_1734), .Y(n_1768) );
AND2x2_ASAP7_75t_L g1776 ( .A(n_1681), .B(n_1777), .Y(n_1776) );
AOI322xp5_ASAP7_75t_L g1795 ( .A1(n_1681), .A2(n_1752), .A3(n_1796), .B1(n_1800), .B2(n_1801), .C1(n_1805), .C2(n_1806), .Y(n_1795) );
NAND2xp5_ASAP7_75t_L g1834 ( .A(n_1681), .B(n_1835), .Y(n_1834) );
NAND2xp5_ASAP7_75t_L g1851 ( .A(n_1681), .B(n_1852), .Y(n_1851) );
NAND2xp5_ASAP7_75t_L g1880 ( .A(n_1681), .B(n_1742), .Y(n_1880) );
O2A1O1Ixp33_ASAP7_75t_SL g1886 ( .A1(n_1681), .A2(n_1736), .B(n_1751), .C(n_1836), .Y(n_1886) );
INVx4_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx4_ASAP7_75t_L g1732 ( .A(n_1682), .Y(n_1732) );
NAND2xp5_ASAP7_75t_SL g1741 ( .A(n_1682), .B(n_1698), .Y(n_1741) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1682), .B(n_1770), .Y(n_1769) );
NOR2xp33_ASAP7_75t_L g1785 ( .A(n_1682), .B(n_1717), .Y(n_1785) );
OR2x2_ASAP7_75t_L g1804 ( .A(n_1682), .B(n_1698), .Y(n_1804) );
NOR2xp33_ASAP7_75t_L g1805 ( .A(n_1682), .B(n_1703), .Y(n_1805) );
NAND2xp5_ASAP7_75t_L g1831 ( .A(n_1682), .B(n_1811), .Y(n_1831) );
AND2x2_ASAP7_75t_L g1863 ( .A(n_1682), .B(n_1771), .Y(n_1863) );
AOI321xp33_ASAP7_75t_R g1875 ( .A1(n_1682), .A2(n_1710), .A3(n_1769), .B1(n_1781), .B2(n_1800), .C(n_1876), .Y(n_1875) );
AND2x4_ASAP7_75t_SL g1682 ( .A(n_1683), .B(n_1691), .Y(n_1682) );
AND2x4_ASAP7_75t_L g1684 ( .A(n_1685), .B(n_1686), .Y(n_1684) );
AND2x6_ASAP7_75t_L g1689 ( .A(n_1685), .B(n_1690), .Y(n_1689) );
AND2x6_ASAP7_75t_L g1692 ( .A(n_1685), .B(n_1693), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1685), .B(n_1695), .Y(n_1694) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_1685), .B(n_1695), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1716 ( .A(n_1685), .B(n_1695), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1761 ( .A(n_1685), .B(n_1686), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1688), .Y(n_1686) );
INVx2_ASAP7_75t_L g1763 ( .A(n_1689), .Y(n_1763) );
INVx2_ASAP7_75t_L g1892 ( .A(n_1692), .Y(n_1892) );
OAI21xp5_ASAP7_75t_L g1978 ( .A1(n_1693), .A2(n_1979), .B(n_1980), .Y(n_1978) );
AOI221xp5_ASAP7_75t_L g1884 ( .A1(n_1696), .A2(n_1826), .B1(n_1849), .B2(n_1885), .C(n_1886), .Y(n_1884) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1702), .Y(n_1696) );
OR2x2_ASAP7_75t_L g1746 ( .A(n_1697), .B(n_1703), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1770 ( .A(n_1697), .B(n_1771), .Y(n_1770) );
OR2x2_ASAP7_75t_L g1836 ( .A(n_1697), .B(n_1736), .Y(n_1836) );
AND2x2_ASAP7_75t_L g1866 ( .A(n_1697), .B(n_1815), .Y(n_1866) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
NAND2xp5_ASAP7_75t_L g1784 ( .A(n_1698), .B(n_1707), .Y(n_1784) );
OR2x2_ASAP7_75t_L g1788 ( .A(n_1698), .B(n_1704), .Y(n_1788) );
AND2x2_ASAP7_75t_L g1790 ( .A(n_1698), .B(n_1742), .Y(n_1790) );
AND2x2_ASAP7_75t_L g1793 ( .A(n_1698), .B(n_1794), .Y(n_1793) );
AND2x2_ASAP7_75t_L g1847 ( .A(n_1698), .B(n_1772), .Y(n_1847) );
OR2x2_ASAP7_75t_L g1883 ( .A(n_1698), .B(n_1772), .Y(n_1883) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1699), .B(n_1700), .Y(n_1698) );
AND2x2_ASAP7_75t_L g1735 ( .A(n_1699), .B(n_1700), .Y(n_1735) );
NAND2xp5_ASAP7_75t_L g1775 ( .A(n_1702), .B(n_1776), .Y(n_1775) );
NAND3xp33_ASAP7_75t_L g1829 ( .A(n_1702), .B(n_1821), .C(n_1830), .Y(n_1829) );
NAND2xp5_ASAP7_75t_L g1843 ( .A(n_1702), .B(n_1828), .Y(n_1843) );
AND2x2_ASAP7_75t_L g1874 ( .A(n_1702), .B(n_1740), .Y(n_1874) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1703), .Y(n_1702) );
OR2x2_ASAP7_75t_L g1824 ( .A(n_1703), .B(n_1804), .Y(n_1824) );
OR2x2_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1707), .Y(n_1703) );
NAND2xp5_ASAP7_75t_L g1736 ( .A(n_1704), .B(n_1737), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_1704), .B(n_1707), .Y(n_1742) );
INVx2_ASAP7_75t_L g1772 ( .A(n_1704), .Y(n_1772) );
NAND2x1p5_ASAP7_75t_L g1704 ( .A(n_1705), .B(n_1706), .Y(n_1704) );
INVx1_ASAP7_75t_L g1737 ( .A(n_1707), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1707), .B(n_1772), .Y(n_1771) );
INVx1_ASAP7_75t_L g1794 ( .A(n_1707), .Y(n_1794) );
OR2x2_ASAP7_75t_L g1853 ( .A(n_1707), .B(n_1735), .Y(n_1853) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1709), .Y(n_1707) );
AOI221xp5_ASAP7_75t_L g1865 ( .A1(n_1710), .A2(n_1755), .B1(n_1866), .B2(n_1867), .C(n_1868), .Y(n_1865) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
OR2x2_ASAP7_75t_L g1711 ( .A(n_1712), .B(n_1717), .Y(n_1711) );
AOI221xp5_ASAP7_75t_L g1766 ( .A1(n_1712), .A2(n_1752), .B1(n_1767), .B2(n_1769), .C(n_1773), .Y(n_1766) );
AOI221xp5_ASAP7_75t_L g1782 ( .A1(n_1712), .A2(n_1783), .B1(n_1785), .B2(n_1786), .C(n_1791), .Y(n_1782) );
OAI322xp33_ASAP7_75t_L g1840 ( .A1(n_1712), .A2(n_1735), .A3(n_1841), .B1(n_1843), .B2(n_1844), .C1(n_1845), .C2(n_1846), .Y(n_1840) );
AND2x2_ASAP7_75t_L g1862 ( .A(n_1712), .B(n_1828), .Y(n_1862) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
INVx3_ASAP7_75t_L g1728 ( .A(n_1713), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1713), .B(n_1745), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1780 ( .A(n_1713), .B(n_1721), .Y(n_1780) );
OR2x2_ASAP7_75t_L g1812 ( .A(n_1713), .B(n_1721), .Y(n_1812) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1714), .B(n_1715), .Y(n_1713) );
AOI21xp33_ASAP7_75t_L g1889 ( .A1(n_1717), .A2(n_1768), .B(n_1789), .Y(n_1889) );
OR2x2_ASAP7_75t_L g1717 ( .A(n_1718), .B(n_1721), .Y(n_1717) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1718), .Y(n_1733) );
INVx1_ASAP7_75t_L g1749 ( .A(n_1718), .Y(n_1749) );
NAND2xp5_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1720), .Y(n_1718) );
A2O1A1Ixp33_ASAP7_75t_L g1738 ( .A1(n_1721), .A2(n_1739), .B(n_1743), .C(n_1747), .Y(n_1738) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1721), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1752 ( .A(n_1721), .B(n_1728), .Y(n_1752) );
OR2x2_ASAP7_75t_L g1778 ( .A(n_1721), .B(n_1749), .Y(n_1778) );
OAI22xp5_ASAP7_75t_L g1786 ( .A1(n_1721), .A2(n_1787), .B1(n_1788), .B2(n_1789), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1800 ( .A(n_1721), .B(n_1733), .Y(n_1800) );
INVx2_ASAP7_75t_L g1821 ( .A(n_1721), .Y(n_1821) );
INVx2_ASAP7_75t_L g1721 ( .A(n_1722), .Y(n_1721) );
OR2x2_ASAP7_75t_L g1814 ( .A(n_1722), .B(n_1749), .Y(n_1814) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1723), .B(n_1724), .Y(n_1722) );
NAND2xp5_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1738), .Y(n_1725) );
NAND2xp5_ASAP7_75t_L g1726 ( .A(n_1727), .B(n_1729), .Y(n_1726) );
CKINVDCx14_ASAP7_75t_R g1727 ( .A(n_1728), .Y(n_1727) );
NAND2xp5_ASAP7_75t_L g1807 ( .A(n_1728), .B(n_1733), .Y(n_1807) );
OR2x2_ASAP7_75t_L g1839 ( .A(n_1728), .B(n_1748), .Y(n_1839) );
OR2x2_ASAP7_75t_L g1844 ( .A(n_1728), .B(n_1733), .Y(n_1844) );
OR2x2_ASAP7_75t_L g1845 ( .A(n_1728), .B(n_1778), .Y(n_1845) );
AND2x2_ASAP7_75t_L g1849 ( .A(n_1728), .B(n_1777), .Y(n_1849) );
O2A1O1Ixp33_ASAP7_75t_SL g1868 ( .A1(n_1728), .A2(n_1799), .B(n_1869), .C(n_1871), .Y(n_1868) );
OR2x2_ASAP7_75t_L g1882 ( .A(n_1728), .B(n_1814), .Y(n_1882) );
A2O1A1Ixp33_ASAP7_75t_R g1887 ( .A1(n_1728), .A2(n_1842), .B(n_1888), .C(n_1889), .Y(n_1887) );
AOI221xp5_ASAP7_75t_L g1817 ( .A1(n_1729), .A2(n_1752), .B1(n_1778), .B2(n_1818), .C(n_1823), .Y(n_1817) );
NOR2xp33_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1734), .Y(n_1729) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1731), .Y(n_1730) );
OAI21xp33_ASAP7_75t_L g1779 ( .A1(n_1731), .A2(n_1780), .B(n_1781), .Y(n_1779) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1732), .B(n_1733), .Y(n_1731) );
AND2x2_ASAP7_75t_L g1755 ( .A(n_1732), .B(n_1756), .Y(n_1755) );
NOR2x1_ASAP7_75t_L g1815 ( .A(n_1732), .B(n_1798), .Y(n_1815) );
NAND2x1_ASAP7_75t_L g1819 ( .A(n_1732), .B(n_1790), .Y(n_1819) );
CKINVDCx5p33_ASAP7_75t_R g1828 ( .A(n_1732), .Y(n_1828) );
NOR2xp33_ASAP7_75t_L g1870 ( .A(n_1732), .B(n_1745), .Y(n_1870) );
INVx2_ASAP7_75t_L g1811 ( .A(n_1733), .Y(n_1811) );
AND2x2_ASAP7_75t_L g1827 ( .A(n_1733), .B(n_1828), .Y(n_1827) );
NAND2xp5_ASAP7_75t_L g1783 ( .A(n_1734), .B(n_1784), .Y(n_1783) );
OR2x2_ASAP7_75t_L g1734 ( .A(n_1735), .B(n_1736), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1781 ( .A(n_1735), .B(n_1771), .Y(n_1781) );
OR2x2_ASAP7_75t_L g1797 ( .A(n_1735), .B(n_1798), .Y(n_1797) );
AOI321xp33_ASAP7_75t_L g1859 ( .A1(n_1735), .A2(n_1757), .A3(n_1806), .B1(n_1860), .B2(n_1862), .C(n_1863), .Y(n_1859) );
OAI221xp5_ASAP7_75t_L g1750 ( .A1(n_1736), .A2(n_1751), .B1(n_1753), .B2(n_1754), .C(n_1757), .Y(n_1750) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1736), .Y(n_1756) );
NAND2xp5_ASAP7_75t_L g1860 ( .A(n_1736), .B(n_1861), .Y(n_1860) );
INVx1_ASAP7_75t_L g1774 ( .A(n_1739), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1740), .B(n_1742), .Y(n_1739) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1798 ( .A(n_1742), .Y(n_1798) );
NAND2xp5_ASAP7_75t_L g1802 ( .A(n_1742), .B(n_1803), .Y(n_1802) );
OAI31xp33_ASAP7_75t_L g1808 ( .A1(n_1743), .A2(n_1809), .A3(n_1813), .B(n_1815), .Y(n_1808) );
NOR2xp33_ASAP7_75t_L g1743 ( .A(n_1744), .B(n_1746), .Y(n_1743) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1744), .Y(n_1753) );
AOI221xp5_ASAP7_75t_L g1848 ( .A1(n_1744), .A2(n_1849), .B1(n_1850), .B2(n_1854), .C(n_1855), .Y(n_1848) );
OAI22xp5_ASAP7_75t_L g1818 ( .A1(n_1745), .A2(n_1819), .B1(n_1820), .B2(n_1822), .Y(n_1818) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1746), .Y(n_1858) );
OAI211xp5_ASAP7_75t_L g1773 ( .A1(n_1747), .A2(n_1774), .B(n_1775), .C(n_1779), .Y(n_1773) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1751 ( .A(n_1748), .B(n_1752), .Y(n_1751) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
NOR2xp33_ASAP7_75t_L g1872 ( .A(n_1749), .B(n_1873), .Y(n_1872) );
A2O1A1Ixp33_ASAP7_75t_L g1877 ( .A1(n_1749), .A2(n_1780), .B(n_1815), .C(n_1837), .Y(n_1877) );
AND2x2_ASAP7_75t_L g1885 ( .A(n_1752), .B(n_1827), .Y(n_1885) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1755), .Y(n_1754) );
INVx2_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1759), .Y(n_1758) );
INVx1_ASAP7_75t_L g1759 ( .A(n_1760), .Y(n_1759) );
OAI221xp5_ASAP7_75t_L g1760 ( .A1(n_1761), .A2(n_1762), .B1(n_1763), .B2(n_1764), .C(n_1765), .Y(n_1760) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1768), .Y(n_1767) );
NAND2xp5_ASAP7_75t_L g1822 ( .A(n_1771), .B(n_1803), .Y(n_1822) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1771), .Y(n_1861) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1776), .Y(n_1787) );
NAND2xp5_ASAP7_75t_L g1792 ( .A(n_1776), .B(n_1793), .Y(n_1792) );
CKINVDCx5p33_ASAP7_75t_R g1777 ( .A(n_1778), .Y(n_1777) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1784), .Y(n_1888) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1788), .Y(n_1826) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
INVxp67_ASAP7_75t_L g1791 ( .A(n_1792), .Y(n_1791) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1793), .Y(n_1799) );
NAND2xp5_ASAP7_75t_SL g1796 ( .A(n_1797), .B(n_1799), .Y(n_1796) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1797), .Y(n_1854) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1802), .Y(n_1801) );
OAI211xp5_ASAP7_75t_L g1878 ( .A1(n_1803), .A2(n_1879), .B(n_1881), .C(n_1883), .Y(n_1878) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1804), .Y(n_1803) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
OR2x2_ASAP7_75t_L g1810 ( .A(n_1811), .B(n_1812), .Y(n_1810) );
CKINVDCx5p33_ASAP7_75t_R g1813 ( .A(n_1814), .Y(n_1813) );
OAI211xp5_ASAP7_75t_L g1823 ( .A1(n_1814), .A2(n_1824), .B(n_1825), .C(n_1829), .Y(n_1823) );
NAND4xp25_ASAP7_75t_L g1816 ( .A(n_1817), .B(n_1832), .C(n_1848), .D(n_1859), .Y(n_1816) );
NAND3xp33_ASAP7_75t_L g1825 ( .A(n_1820), .B(n_1826), .C(n_1827), .Y(n_1825) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1821), .Y(n_1820) );
INVx1_ASAP7_75t_L g1837 ( .A(n_1824), .Y(n_1837) );
INVx1_ASAP7_75t_L g1830 ( .A(n_1831), .Y(n_1830) );
O2A1O1Ixp33_ASAP7_75t_L g1832 ( .A1(n_1833), .A2(n_1837), .B(n_1838), .C(n_1840), .Y(n_1832) );
INVxp67_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1836), .Y(n_1835) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1839), .Y(n_1838) );
INVx1_ASAP7_75t_L g1841 ( .A(n_1842), .Y(n_1841) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1844), .Y(n_1857) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1845), .Y(n_1867) );
CKINVDCx14_ASAP7_75t_R g1846 ( .A(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g1850 ( .A(n_1851), .Y(n_1850) );
INVxp67_ASAP7_75t_L g1852 ( .A(n_1853), .Y(n_1852) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1856), .Y(n_1855) );
NAND2xp5_ASAP7_75t_L g1856 ( .A(n_1857), .B(n_1858), .Y(n_1856) );
NAND4xp25_ASAP7_75t_L g1864 ( .A(n_1865), .B(n_1875), .C(n_1884), .D(n_1887), .Y(n_1864) );
INVx1_ASAP7_75t_L g1869 ( .A(n_1870), .Y(n_1869) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1872), .Y(n_1871) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1874), .Y(n_1873) );
NAND2xp5_ASAP7_75t_SL g1876 ( .A(n_1877), .B(n_1878), .Y(n_1876) );
INVxp67_ASAP7_75t_SL g1879 ( .A(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1882), .Y(n_1881) );
CKINVDCx20_ASAP7_75t_R g1890 ( .A(n_1891), .Y(n_1890) );
CKINVDCx20_ASAP7_75t_R g1891 ( .A(n_1892), .Y(n_1891) );
NAND3xp33_ASAP7_75t_L g1894 ( .A(n_1895), .B(n_1909), .C(n_1912), .Y(n_1894) );
NAND2xp5_ASAP7_75t_L g1896 ( .A(n_1897), .B(n_1900), .Y(n_1896) );
INVxp67_ASAP7_75t_L g1937 ( .A(n_1908), .Y(n_1937) );
INVx3_ASAP7_75t_L g1925 ( .A(n_1926), .Y(n_1925) );
HB1xp67_ASAP7_75t_L g1929 ( .A(n_1930), .Y(n_1929) );
BUFx3_ASAP7_75t_L g1930 ( .A(n_1931), .Y(n_1930) );
INVx1_ASAP7_75t_L g1933 ( .A(n_1934), .Y(n_1933) );
AND3x2_ASAP7_75t_L g1934 ( .A(n_1935), .B(n_1957), .C(n_1960), .Y(n_1934) );
AOI211xp5_ASAP7_75t_SL g1935 ( .A1(n_1936), .A2(n_1937), .B(n_1938), .C(n_1941), .Y(n_1935) );
INVx1_ASAP7_75t_L g1944 ( .A(n_1945), .Y(n_1944) );
INVx2_ASAP7_75t_L g1952 ( .A(n_1953), .Y(n_1952) );
INVxp67_ASAP7_75t_L g1967 ( .A(n_1968), .Y(n_1967) );
INVx2_ASAP7_75t_L g1970 ( .A(n_1971), .Y(n_1970) );
HB1xp67_ASAP7_75t_L g1977 ( .A(n_1978), .Y(n_1977) );
INVx1_ASAP7_75t_L g1980 ( .A(n_1981), .Y(n_1980) );
endmodule