module fake_jpeg_2883_n_171 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_44),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_1),
.C(n_4),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_55),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_48),
.B1(n_43),
.B2(n_38),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_15),
.B1(n_22),
.B2(n_6),
.Y(n_83)
);

NAND2x1_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_28),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_58),
.B(n_59),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_33),
.B(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_24),
.Y(n_72)
);

MAJx2_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_28),
.C(n_22),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_16),
.B1(n_28),
.B2(n_26),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_28),
.B1(n_26),
.B2(n_15),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_10),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_12),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_99),
.B(n_62),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_73),
.Y(n_114)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_85),
.B1(n_89),
.B2(n_98),
.Y(n_117)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_5),
.C(n_7),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_88),
.C(n_57),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_5),
.C(n_7),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_7),
.B1(n_9),
.B2(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_9),
.B1(n_66),
.B2(n_63),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_50),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_65),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_109),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_115),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_114),
.B(n_95),
.Y(n_129)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_75),
.B1(n_67),
.B2(n_74),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_79),
.B1(n_100),
.B2(n_80),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_78),
.C(n_67),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_78),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_122),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_125),
.Y(n_140)
);

OAI22x1_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_87),
.B1(n_95),
.B2(n_93),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_115),
.B(n_109),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_88),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_127),
.B(n_123),
.Y(n_135)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_129),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_117),
.B1(n_104),
.B2(n_119),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_126),
.B1(n_125),
.B2(n_131),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_112),
.B(n_105),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_118),
.B(n_113),
.Y(n_153)
);

OAI21x1_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_140),
.B(n_143),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_148),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_112),
.B(n_134),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_150),
.B(n_152),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_145),
.B(n_90),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_96),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_132),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_90),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_153),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_158),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_140),
.C(n_144),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_86),
.C(n_137),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_163),
.C(n_159),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_155),
.A2(n_141),
.B1(n_117),
.B2(n_139),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_121),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_139),
.C(n_84),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_154),
.C(n_92),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_165),
.A2(n_166),
.B(n_160),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_91),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_168),
.C(n_68),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_60),
.Y(n_171)
);


endmodule