module fake_netlist_6_4273_n_1817 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1817);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1817;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_27),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_72),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_100),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_134),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_13),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_89),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_63),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_84),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_92),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_68),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_124),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_59),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_60),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_3),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_61),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_160),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_10),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_150),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_8),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_76),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_30),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_148),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_6),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_69),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_107),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_102),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_70),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_83),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_91),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_157),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_18),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_22),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_71),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_166),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_56),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_110),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_142),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_147),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_109),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_88),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_30),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_51),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_93),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_106),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_23),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_78),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_179),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_1),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_21),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_39),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_73),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_50),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_90),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_57),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_103),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_96),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_54),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_81),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_132),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_20),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_164),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_127),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_114),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_20),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_118),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_67),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_1),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_37),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_98),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_13),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_3),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_32),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_44),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_75),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_63),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_133),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_121),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_29),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_165),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_29),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_46),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_2),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_23),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_87),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_125),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_35),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_138),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_34),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_168),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_31),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_19),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_141),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_111),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_174),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_173),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_6),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_116),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_26),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_32),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_167),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_16),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_95),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_14),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_156),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_42),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_17),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_10),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_178),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_82),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_16),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_41),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_151),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_60),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_26),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_74),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_113),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_80),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_45),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_175),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_94),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_41),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_40),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_119),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_62),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_155),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_11),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_131),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_50),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_145),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_108),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_104),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_44),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_56),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_27),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_7),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_11),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_55),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_62),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_85),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_0),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_172),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_24),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_144),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_171),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_137),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_54),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_105),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_40),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_65),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_101),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_99),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_115),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_163),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_31),
.Y(n_345)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_143),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_135),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_79),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_176),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_47),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_52),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_45),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_58),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_21),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_34),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_46),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_19),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_161),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_152),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_15),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_24),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_36),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_36),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_53),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_180),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_182),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_261),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_183),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_262),
.B(n_4),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_221),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_184),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_267),
.B(n_4),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_188),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_261),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_244),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_244),
.B(n_5),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_261),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_199),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_261),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_228),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_330),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_338),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_261),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_261),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_200),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_190),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_237),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_5),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_191),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_200),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_193),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_195),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_238),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_238),
.Y(n_394)
);

INVxp33_ASAP7_75t_L g395 ( 
.A(n_199),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_181),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_330),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_301),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_213),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_357),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_196),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_185),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_226),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_202),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_267),
.B(n_7),
.Y(n_406)
);

INVxp33_ASAP7_75t_SL g407 ( 
.A(n_201),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_357),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_187),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_215),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_203),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_288),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_288),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_288),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_282),
.B(n_8),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_255),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_347),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_282),
.B(n_9),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_204),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_302),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_192),
.B(n_9),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_302),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_215),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_208),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_192),
.B(n_194),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_213),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_302),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_210),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_337),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_211),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_189),
.B(n_12),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_337),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_337),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_217),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_227),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_227),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_220),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_230),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_341),
.B(n_12),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_R g440 ( 
.A(n_341),
.B(n_15),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_230),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_224),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_231),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_231),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_234),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_225),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_232),
.Y(n_447)
);

BUFx2_ASAP7_75t_SL g448 ( 
.A(n_326),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_194),
.B(n_17),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_236),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_234),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_246),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_239),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_197),
.B(n_206),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_239),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_205),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_248),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_242),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_242),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_384),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_365),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_367),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_367),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_374),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_374),
.Y(n_467)
);

AND2x2_ASAP7_75t_SL g468 ( 
.A(n_406),
.B(n_300),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_377),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_375),
.A2(n_309),
.B1(n_363),
.B2(n_305),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_410),
.B(n_240),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_404),
.B(n_226),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_377),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_366),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_371),
.B(n_226),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_373),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_386),
.B(n_336),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_389),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_404),
.B(n_336),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_404),
.B(n_336),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_368),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_379),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_383),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_391),
.B(n_275),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_392),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_370),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_388),
.B(n_439),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_376),
.B(n_341),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_402),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_380),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_405),
.B(n_419),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_430),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_396),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_385),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_434),
.Y(n_499)
);

AND2x2_ASAP7_75t_SL g500 ( 
.A(n_372),
.B(n_300),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_442),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_446),
.B(n_275),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_385),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_436),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_293),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_381),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_R g508 ( 
.A(n_409),
.B(n_249),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_447),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_390),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_417),
.B(n_311),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_436),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_412),
.B(n_293),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_457),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_390),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_411),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_393),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_413),
.B(n_240),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_387),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_393),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_407),
.B(n_214),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_424),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_394),
.B(n_266),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_456),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_394),
.Y(n_527)
);

NOR2xp67_ASAP7_75t_L g528 ( 
.A(n_398),
.B(n_279),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_398),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_399),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_438),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_397),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_441),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_428),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_416),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_413),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_538),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_476),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_538),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_369),
.C(n_415),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_468),
.B(n_186),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_538),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_489),
.B(n_382),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_483),
.B(n_431),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_460),
.Y(n_547)
);

NOR2x1p5_ASAP7_75t_L g548 ( 
.A(n_463),
.B(n_376),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_472),
.B(n_448),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_493),
.B(n_448),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_460),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_469),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_490),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_476),
.Y(n_554)
);

INVx5_ASAP7_75t_L g555 ( 
.A(n_490),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_468),
.A2(n_500),
.B1(n_490),
.B2(n_454),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_470),
.B(n_326),
.Y(n_557)
);

INVx4_ASAP7_75t_SL g558 ( 
.A(n_490),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_473),
.B(n_300),
.Y(n_559)
);

BUFx4f_ASAP7_75t_L g560 ( 
.A(n_468),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_461),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_477),
.B(n_437),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_476),
.Y(n_564)
);

AND3x2_ASAP7_75t_L g565 ( 
.A(n_509),
.B(n_418),
.C(n_421),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_470),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_470),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_473),
.B(n_414),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_523),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_523),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_488),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_489),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_462),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_479),
.B(n_450),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_496),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_500),
.B(n_186),
.Y(n_576)
);

AO22x2_ASAP7_75t_L g577 ( 
.A1(n_471),
.A2(n_353),
.B1(n_304),
.B2(n_328),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_462),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_490),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_489),
.B(n_425),
.Y(n_580)
);

NAND3xp33_ASAP7_75t_L g581 ( 
.A(n_472),
.B(n_440),
.C(n_449),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_496),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_500),
.A2(n_329),
.B1(n_278),
.B2(n_354),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_498),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_486),
.B(n_452),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_490),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_490),
.A2(n_329),
.B1(n_278),
.B2(n_354),
.Y(n_587)
);

INVx4_ASAP7_75t_SL g588 ( 
.A(n_473),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_489),
.B(n_253),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_498),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_492),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_507),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_481),
.A2(n_360),
.B1(n_247),
.B2(n_353),
.Y(n_593)
);

AO22x2_ASAP7_75t_L g594 ( 
.A1(n_512),
.A2(n_247),
.B1(n_290),
.B2(n_294),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_523),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_496),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_508),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_502),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_464),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_520),
.B(n_431),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_SL g601 ( 
.A(n_503),
.B(n_198),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_495),
.B(n_395),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_469),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_464),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_466),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_466),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_481),
.B(n_295),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_467),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_481),
.B(n_420),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_469),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_469),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_517),
.B(n_420),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_502),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_L g614 ( 
.A1(n_526),
.A2(n_297),
.B1(n_324),
.B2(n_325),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_506),
.B(n_422),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_482),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_475),
.B(n_422),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_469),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_482),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_505),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_467),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_484),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_482),
.B(n_427),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_469),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_484),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_513),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_474),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_482),
.B(n_212),
.Y(n_629)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_474),
.Y(n_630)
);

INVx8_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_506),
.B(n_429),
.Y(n_632)
);

OAI22xp33_ASAP7_75t_L g633 ( 
.A1(n_507),
.A2(n_312),
.B1(n_339),
.B2(n_361),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_504),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_537),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_506),
.B(n_429),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_514),
.B(n_432),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_474),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_514),
.B(n_432),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_504),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_480),
.B(n_487),
.Y(n_641)
);

BUFx4f_ASAP7_75t_L g642 ( 
.A(n_474),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_513),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_531),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_531),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_514),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_514),
.B(n_433),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_491),
.B(n_212),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_504),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_504),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_519),
.B(n_433),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_504),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_465),
.B(n_252),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_532),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_532),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_494),
.B(n_378),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_519),
.B(n_534),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_524),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_499),
.A2(n_283),
.B1(n_269),
.B2(n_259),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_533),
.B(n_400),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_534),
.B(n_399),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_501),
.B(n_233),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_535),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_510),
.B(n_233),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_515),
.B(n_426),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_535),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_504),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_511),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_525),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_527),
.A2(n_298),
.B1(n_294),
.B2(n_360),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_525),
.B(n_453),
.C(n_444),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_474),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_527),
.A2(n_290),
.B1(n_351),
.B2(n_333),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_537),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_528),
.B(n_197),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_465),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_485),
.Y(n_677)
);

AND2x6_ASAP7_75t_L g678 ( 
.A(n_527),
.B(n_300),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_485),
.Y(n_679)
);

NAND2x1p5_ASAP7_75t_L g680 ( 
.A(n_528),
.B(n_206),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_485),
.B(n_256),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_485),
.Y(n_682)
);

AND2x6_ASAP7_75t_L g683 ( 
.A(n_527),
.B(n_300),
.Y(n_683)
);

INVx8_ASAP7_75t_L g684 ( 
.A(n_485),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_602),
.B(n_536),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_560),
.A2(n_274),
.B1(n_264),
.B2(n_277),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_599),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_556),
.B(n_529),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_560),
.A2(n_298),
.B(n_304),
.C(n_328),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_R g690 ( 
.A(n_658),
.B(n_592),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_599),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_572),
.B(n_529),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_566),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_572),
.B(n_529),
.Y(n_694)
);

AND2x6_ASAP7_75t_SL g695 ( 
.A(n_641),
.B(n_333),
.Y(n_695)
);

NOR2x1p5_ASAP7_75t_L g696 ( 
.A(n_542),
.B(n_207),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_617),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_549),
.B(n_580),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_549),
.B(n_529),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_617),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_560),
.B(n_300),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_601),
.A2(n_285),
.B1(n_287),
.B2(n_291),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_656),
.B(n_222),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_543),
.A2(n_245),
.B1(n_284),
.B2(n_303),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_618),
.B(n_362),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_576),
.A2(n_543),
.B(n_684),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_620),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_665),
.B(n_222),
.Y(n_708)
);

CKINVDCx11_ASAP7_75t_R g709 ( 
.A(n_592),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_566),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_620),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_555),
.B(n_320),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_568),
.B(n_511),
.Y(n_713)
);

NOR3x1_ASAP7_75t_L g714 ( 
.A(n_648),
.B(n_351),
.C(n_345),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_571),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_563),
.B(n_209),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_604),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_581),
.B(n_443),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_545),
.B(n_589),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_574),
.B(n_218),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_624),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_604),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_576),
.A2(n_485),
.B(n_497),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_624),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_646),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_555),
.B(n_320),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_612),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_555),
.B(n_553),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_583),
.A2(n_245),
.B1(n_284),
.B2(n_303),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_600),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_646),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_585),
.B(n_648),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_544),
.B(n_615),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_661),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_615),
.B(n_521),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_609),
.A2(n_345),
.B(n_216),
.C(n_335),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_607),
.A2(n_332),
.B(n_223),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_555),
.B(n_553),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_662),
.B(n_219),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_658),
.Y(n_740)
);

INVx8_ASAP7_75t_L g741 ( 
.A(n_550),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_657),
.B(n_597),
.Y(n_742)
);

NAND2x1p5_ASAP7_75t_L g743 ( 
.A(n_555),
.B(n_553),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_662),
.B(n_235),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_SL g745 ( 
.A(n_631),
.B(n_331),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_L g746 ( 
.A(n_633),
.B(n_265),
.C(n_271),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_605),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_639),
.B(n_216),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_629),
.A2(n_223),
.B(n_229),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_579),
.B(n_320),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_569),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_L g752 ( 
.A(n_601),
.B(n_268),
.C(n_270),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_647),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_657),
.B(n_222),
.Y(n_754)
);

AND2x6_ASAP7_75t_SL g755 ( 
.A(n_660),
.B(n_443),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_647),
.B(n_229),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_579),
.B(n_320),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_657),
.B(n_241),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_587),
.A2(n_332),
.B1(n_241),
.B2(n_243),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_584),
.B(n_243),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_590),
.B(n_251),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_651),
.A2(n_321),
.B1(n_251),
.B2(n_259),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_664),
.B(n_250),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_598),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_539),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_579),
.B(n_320),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_613),
.B(n_269),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_605),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_606),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_586),
.A2(n_318),
.B1(n_283),
.B2(n_321),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_616),
.B(n_308),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_586),
.B(n_320),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_621),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_664),
.B(n_570),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_627),
.B(n_308),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_643),
.B(n_318),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_586),
.B(n_346),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_L g778 ( 
.A(n_593),
.B(n_260),
.C(n_257),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_559),
.B(n_346),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_606),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_651),
.B(n_222),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_651),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_569),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_669),
.B(n_254),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_644),
.B(n_335),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_558),
.B(n_346),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_645),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_654),
.B(n_342),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_655),
.B(n_342),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_550),
.B(n_445),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_608),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_567),
.B(n_343),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_663),
.B(n_343),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_629),
.A2(n_349),
.B(n_344),
.C(n_451),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_666),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_550),
.B(n_258),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_632),
.B(n_344),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_636),
.B(n_349),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_558),
.B(n_539),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_539),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_637),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_550),
.A2(n_299),
.B1(n_306),
.B2(n_307),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_547),
.B(n_516),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_631),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_594),
.A2(n_346),
.B1(n_311),
.B2(n_516),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_595),
.A2(n_310),
.B1(n_314),
.B2(n_316),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_539),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_660),
.B(n_565),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_558),
.B(n_346),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_614),
.B(n_263),
.C(n_272),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_594),
.A2(n_346),
.B1(n_311),
.B2(n_518),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_557),
.A2(n_364),
.B1(n_276),
.B2(n_280),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_551),
.B(n_530),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_561),
.B(n_322),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_608),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_548),
.A2(n_334),
.B1(n_348),
.B2(n_358),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_541),
.B(n_346),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_660),
.B(n_445),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_562),
.B(n_359),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_622),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_631),
.B(n_451),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_573),
.B(n_346),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_622),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_578),
.B(n_455),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_541),
.B(n_311),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_541),
.B(n_653),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_623),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_L g828 ( 
.A(n_671),
.B(n_66),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_623),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_660),
.B(n_273),
.Y(n_830)
);

O2A1O1Ixp5_ASAP7_75t_L g831 ( 
.A1(n_676),
.A2(n_459),
.B(n_458),
.C(n_455),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_594),
.A2(n_323),
.B1(n_286),
.B2(n_289),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_557),
.B(n_659),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_681),
.A2(n_459),
.B(n_458),
.C(n_408),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_L g835 ( 
.A(n_559),
.B(n_327),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_SL g836 ( 
.A(n_631),
.B(n_591),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_626),
.A2(n_408),
.B(n_401),
.C(n_356),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_626),
.B(n_355),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_675),
.B(n_352),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_557),
.B(n_350),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_688),
.A2(n_619),
.B(n_642),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_826),
.A2(n_684),
.B(n_642),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_698),
.B(n_594),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_706),
.A2(n_642),
.B(n_649),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_SL g845 ( 
.A(n_740),
.B(n_635),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_732),
.B(n_675),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_716),
.A2(n_675),
.B1(n_559),
.B2(n_557),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_705),
.B(n_577),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_742),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_743),
.A2(n_684),
.B(n_603),
.Y(n_850)
);

INVx4_ASAP7_75t_L g851 ( 
.A(n_725),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_701),
.A2(n_634),
.B(n_667),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_725),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_720),
.A2(n_670),
.B(n_673),
.C(n_640),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_743),
.A2(n_611),
.B(n_630),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_701),
.A2(n_699),
.B(n_750),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_715),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_728),
.A2(n_611),
.B(n_630),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_719),
.B(n_680),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_801),
.B(n_680),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_687),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_690),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_687),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_728),
.A2(n_611),
.B(n_603),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_739),
.A2(n_652),
.B(n_650),
.C(n_667),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_693),
.B(n_588),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_725),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_691),
.Y(n_868)
);

NAND2x1_ASAP7_75t_L g869 ( 
.A(n_800),
.B(n_807),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_777),
.A2(n_677),
.B(n_682),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_744),
.A2(n_650),
.B(n_649),
.C(n_652),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_703),
.B(n_708),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_801),
.B(n_552),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_689),
.A2(n_554),
.B(n_582),
.C(n_540),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_763),
.A2(n_668),
.B(n_634),
.C(n_679),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_738),
.A2(n_628),
.B(n_630),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_738),
.A2(n_628),
.B(n_603),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_721),
.A2(n_577),
.B1(n_610),
.B2(n_625),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_735),
.A2(n_628),
.B(n_672),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_727),
.B(n_610),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_734),
.B(n_577),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_713),
.A2(n_625),
.B(n_638),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_757),
.A2(n_564),
.B(n_540),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_685),
.B(n_546),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_689),
.A2(n_564),
.B(n_554),
.C(n_575),
.Y(n_885)
);

NOR2x1_ASAP7_75t_L g886 ( 
.A(n_804),
.B(n_635),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_721),
.A2(n_577),
.B1(n_575),
.B2(n_582),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_725),
.B(n_724),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_753),
.B(n_559),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_724),
.B(n_596),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_765),
.A2(n_596),
.B(n_559),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_733),
.B(n_559),
.Y(n_892)
);

AO32x2_ASAP7_75t_L g893 ( 
.A1(n_770),
.A2(n_832),
.A3(n_782),
.B1(n_783),
.B2(n_802),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_690),
.Y(n_894)
);

NOR2x1_ASAP7_75t_L g895 ( 
.A(n_804),
.B(n_674),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_709),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_737),
.A2(n_315),
.B(n_292),
.C(n_340),
.Y(n_897)
);

AO21x1_ASAP7_75t_L g898 ( 
.A1(n_766),
.A2(n_22),
.B(n_25),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_812),
.B(n_281),
.C(n_296),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_692),
.A2(n_694),
.B(n_766),
.Y(n_900)
);

OAI21xp5_ASAP7_75t_L g901 ( 
.A1(n_772),
.A2(n_683),
.B(n_678),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_792),
.B(n_678),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_777),
.A2(n_799),
.B(n_707),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_799),
.A2(n_678),
.B(n_319),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_707),
.A2(n_317),
.B(n_313),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_790),
.B(n_25),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_800),
.A2(n_77),
.B(n_170),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_800),
.A2(n_177),
.B(n_169),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_792),
.B(n_28),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_800),
.A2(n_162),
.B(n_158),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_723),
.A2(n_149),
.B(n_140),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_807),
.A2(n_136),
.B(n_130),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_729),
.A2(n_28),
.B1(n_33),
.B2(n_35),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_748),
.A2(n_129),
.B(n_128),
.Y(n_914)
);

OR2x6_ASAP7_75t_SL g915 ( 
.A(n_740),
.B(n_33),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_807),
.A2(n_123),
.B(n_122),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_792),
.B(n_764),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_773),
.B(n_37),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_SL g919 ( 
.A1(n_807),
.A2(n_120),
.B(n_112),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_787),
.B(n_38),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_L g921 ( 
.A(n_774),
.B(n_38),
.C(n_39),
.Y(n_921)
);

AO21x1_ASAP7_75t_L g922 ( 
.A1(n_749),
.A2(n_42),
.B(n_43),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_718),
.B(n_43),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_833),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_818),
.B(n_48),
.Y(n_925)
);

BUFx4f_ASAP7_75t_L g926 ( 
.A(n_821),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_754),
.B(n_49),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_782),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_795),
.B(n_55),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_758),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_783),
.B(n_61),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_691),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_717),
.B(n_722),
.Y(n_933)
);

AO21x1_ASAP7_75t_L g934 ( 
.A1(n_817),
.A2(n_64),
.B(n_65),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_696),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_L g936 ( 
.A(n_796),
.B(n_64),
.C(n_86),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_756),
.A2(n_831),
.B(n_736),
.C(n_797),
.Y(n_937)
);

OAI22x1_ASAP7_75t_L g938 ( 
.A1(n_808),
.A2(n_730),
.B1(n_830),
.B2(n_840),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_709),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_731),
.A2(n_711),
.B1(n_697),
.B2(n_700),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_693),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_786),
.A2(n_809),
.B(n_814),
.Y(n_942)
);

NAND3xp33_ASAP7_75t_L g943 ( 
.A(n_784),
.B(n_746),
.C(n_810),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_820),
.B(n_823),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_717),
.B(n_768),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_722),
.A2(n_769),
.B(n_791),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_747),
.Y(n_947)
);

O2A1O1Ixp5_ASAP7_75t_L g948 ( 
.A1(n_834),
.A2(n_798),
.B(n_789),
.C(n_788),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_736),
.A2(n_785),
.B(n_761),
.C(n_767),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_747),
.B(n_768),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_760),
.A2(n_793),
.B(n_776),
.C(n_775),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_780),
.B(n_829),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_819),
.A2(n_817),
.B(n_726),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_L g954 ( 
.A(n_704),
.B(n_741),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_712),
.A2(n_726),
.B(n_813),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_815),
.B(n_827),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_712),
.A2(n_803),
.B(n_822),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_781),
.B(n_838),
.Y(n_958)
);

BUFx4f_ASAP7_75t_L g959 ( 
.A(n_821),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_839),
.A2(n_686),
.B(n_771),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_762),
.B(n_759),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_779),
.A2(n_825),
.B(n_824),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_710),
.B(n_751),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_710),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_779),
.A2(n_825),
.B(n_751),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_805),
.B(n_811),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_835),
.A2(n_794),
.B(n_828),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_702),
.A2(n_778),
.B(n_752),
.C(n_741),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_837),
.A2(n_741),
.B(n_835),
.C(n_816),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_755),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_806),
.A2(n_741),
.B(n_821),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_745),
.B(n_821),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_836),
.A2(n_714),
.B(n_695),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_687),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_826),
.A2(n_743),
.B(n_738),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_732),
.A2(n_560),
.B(n_720),
.C(n_716),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_826),
.A2(n_743),
.B(n_738),
.Y(n_977)
);

OAI22xp33_ASAP7_75t_L g978 ( 
.A1(n_698),
.A2(n_560),
.B1(n_719),
.B2(n_734),
.Y(n_978)
);

O2A1O1Ixp5_ASAP7_75t_L g979 ( 
.A1(n_701),
.A2(n_543),
.B(n_576),
.C(n_737),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_727),
.B(n_698),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_698),
.B(n_732),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_698),
.B(n_732),
.Y(n_982)
);

OAI21xp33_ASAP7_75t_L g983 ( 
.A1(n_705),
.A2(n_720),
.B(n_716),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_701),
.A2(n_543),
.B(n_576),
.C(n_737),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_L g985 ( 
.A(n_740),
.B(n_658),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_L g986 ( 
.A(n_705),
.B(n_732),
.C(n_720),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_698),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_732),
.A2(n_560),
.B1(n_556),
.B2(n_698),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_698),
.B(n_732),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_777),
.A2(n_757),
.B(n_750),
.Y(n_990)
);

OR2x2_ASAP7_75t_SL g991 ( 
.A(n_685),
.B(n_537),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_698),
.B(n_732),
.Y(n_992)
);

AO21x1_ASAP7_75t_L g993 ( 
.A1(n_701),
.A2(n_543),
.B(n_576),
.Y(n_993)
);

NAND2x1p5_ASAP7_75t_L g994 ( 
.A(n_707),
.B(n_804),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_826),
.A2(n_743),
.B(n_738),
.Y(n_995)
);

NAND2x1p5_ASAP7_75t_L g996 ( 
.A(n_707),
.B(n_804),
.Y(n_996)
);

AO22x1_ASAP7_75t_L g997 ( 
.A1(n_732),
.A2(n_705),
.B1(n_720),
.B2(n_716),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_826),
.A2(n_743),
.B(n_738),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_687),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_826),
.A2(n_743),
.B(n_738),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_698),
.B(n_732),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_693),
.B(n_710),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_826),
.A2(n_743),
.B(n_738),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_727),
.B(n_698),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_732),
.A2(n_560),
.B1(n_556),
.B2(n_698),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_687),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_698),
.B(n_732),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_698),
.B(n_732),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_690),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_732),
.A2(n_560),
.B1(n_698),
.B2(n_716),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_980),
.B(n_1004),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_975),
.A2(n_995),
.B(n_977),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_980),
.B(n_1004),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_1002),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_983),
.A2(n_986),
.B(n_923),
.C(n_976),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_SL g1016 ( 
.A1(n_896),
.A2(n_884),
.B1(n_970),
.B2(n_991),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_998),
.A2(n_1003),
.B(n_1000),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_872),
.B(n_849),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_979),
.A2(n_984),
.B(n_988),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_844),
.A2(n_903),
.B(n_879),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_850),
.A2(n_954),
.B(n_855),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_979),
.A2(n_984),
.B(n_1005),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_856),
.A2(n_1010),
.B(n_982),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_SL g1024 ( 
.A1(n_843),
.A2(n_958),
.B(n_892),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_981),
.A2(n_992),
.B1(n_1001),
.B2(n_1008),
.Y(n_1025)
);

AOI21x1_ASAP7_75t_L g1026 ( 
.A1(n_888),
.A2(n_842),
.B(n_900),
.Y(n_1026)
);

AOI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_943),
.A2(n_1007),
.B(n_989),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_997),
.B(n_987),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_1002),
.Y(n_1029)
);

OAI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_948),
.A2(n_937),
.B(n_966),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_987),
.A2(n_923),
.B1(n_848),
.B2(n_972),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_863),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_913),
.A2(n_925),
.B(n_914),
.C(n_961),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_894),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_948),
.A2(n_937),
.B(n_846),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_857),
.Y(n_1036)
);

OAI22x1_ASAP7_75t_L g1037 ( 
.A1(n_972),
.A2(n_935),
.B1(n_925),
.B2(n_881),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_841),
.A2(n_858),
.B(n_864),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_867),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_859),
.B(n_917),
.Y(n_1040)
);

AO21x1_ASAP7_75t_L g1041 ( 
.A1(n_978),
.A2(n_911),
.B(n_960),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_913),
.A2(n_921),
.B(n_924),
.C(n_936),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_932),
.Y(n_1043)
);

NAND2x1_ASAP7_75t_L g1044 ( 
.A(n_851),
.B(n_867),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_876),
.A2(n_877),
.B(n_883),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_990),
.A2(n_852),
.B(n_874),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_962),
.A2(n_854),
.B(n_942),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_985),
.B(n_862),
.Y(n_1048)
);

AOI21x1_ASAP7_75t_L g1049 ( 
.A1(n_888),
.A2(n_967),
.B(n_945),
.Y(n_1049)
);

AOI221xp5_ASAP7_75t_L g1050 ( 
.A1(n_899),
.A2(n_973),
.B1(n_938),
.B2(n_897),
.C(n_936),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_880),
.B(n_927),
.Y(n_1051)
);

NAND2x1_ASAP7_75t_L g1052 ( 
.A(n_851),
.B(n_867),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_906),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_944),
.Y(n_1054)
);

NAND2x1p5_ASAP7_75t_L g1055 ( 
.A(n_866),
.B(n_867),
.Y(n_1055)
);

INVxp67_ASAP7_75t_SL g1056 ( 
.A(n_853),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_885),
.A2(n_953),
.B(n_957),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_963),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_866),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_963),
.B(n_845),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_965),
.A2(n_860),
.B(n_951),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_886),
.B(n_895),
.Y(n_1062)
);

AND3x4_ASAP7_75t_L g1063 ( 
.A(n_899),
.B(n_915),
.C(n_939),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_978),
.B(n_847),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_964),
.B(n_909),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_SL g1066 ( 
.A(n_964),
.B(n_941),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_918),
.B(n_920),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_869),
.Y(n_1068)
);

OA22x2_ASAP7_75t_L g1069 ( 
.A1(n_1009),
.A2(n_878),
.B1(n_887),
.B2(n_929),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_941),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_902),
.A2(n_873),
.B(n_956),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_952),
.A2(n_955),
.B(n_993),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_853),
.B(n_868),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_889),
.A2(n_891),
.B(n_890),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_890),
.A2(n_969),
.B(n_933),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_947),
.B(n_999),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_931),
.Y(n_1077)
);

BUFx12f_ASAP7_75t_L g1078 ( 
.A(n_994),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_974),
.B(n_1006),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_922),
.A2(n_875),
.A3(n_871),
.B(n_865),
.Y(n_1080)
);

OAI22x1_ASAP7_75t_L g1081 ( 
.A1(n_994),
.A2(n_996),
.B1(n_959),
.B2(n_926),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_940),
.B(n_905),
.Y(n_1082)
);

NOR4xp25_ASAP7_75t_L g1083 ( 
.A(n_930),
.B(n_928),
.C(n_968),
.D(n_949),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_950),
.B(n_968),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_996),
.B(n_971),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_959),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_893),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_934),
.B(n_898),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_926),
.B(n_904),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_893),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_919),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_901),
.A2(n_907),
.B(n_908),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_910),
.A2(n_916),
.B(n_912),
.C(n_893),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_893),
.B(n_980),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_975),
.A2(n_743),
.B(n_579),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_849),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_975),
.A2(n_743),
.B(n_579),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_983),
.A2(n_560),
.B(n_986),
.C(n_923),
.Y(n_1098)
);

O2A1O1Ixp5_ASAP7_75t_L g1099 ( 
.A1(n_997),
.A2(n_976),
.B(n_701),
.C(n_986),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_867),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1002),
.B(n_941),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_983),
.A2(n_560),
.B(n_986),
.C(n_923),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_863),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_863),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_946),
.A2(n_870),
.B(n_882),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_946),
.A2(n_870),
.B(n_882),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_983),
.A2(n_560),
.B(n_986),
.C(n_923),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_983),
.A2(n_560),
.B(n_986),
.C(n_923),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_851),
.B(n_866),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_946),
.A2(n_870),
.B(n_882),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_986),
.A2(n_984),
.B(n_979),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_867),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_975),
.A2(n_743),
.B(n_579),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_861),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1010),
.B(n_560),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_983),
.A2(n_560),
.B(n_986),
.C(n_923),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_946),
.A2(n_870),
.B(n_882),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_861),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_980),
.B(n_1004),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_857),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_986),
.B(n_983),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_980),
.B(n_1004),
.Y(n_1122)
);

INVx1_ASAP7_75t_SL g1123 ( 
.A(n_857),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_851),
.B(n_866),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_975),
.A2(n_743),
.B(n_579),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_975),
.A2(n_743),
.B(n_579),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_975),
.A2(n_743),
.B(n_579),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_986),
.A2(n_984),
.B(n_979),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_946),
.A2(n_870),
.B(n_882),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1002),
.B(n_866),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_975),
.A2(n_743),
.B(n_579),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_946),
.A2(n_870),
.B(n_882),
.Y(n_1132)
);

NAND2xp33_ASAP7_75t_L g1133 ( 
.A(n_976),
.B(n_556),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_L g1134 ( 
.A1(n_888),
.A2(n_701),
.B(n_1003),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_975),
.A2(n_743),
.B(n_579),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_983),
.A2(n_560),
.B(n_986),
.C(n_923),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_993),
.A2(n_1005),
.A3(n_988),
.B(n_937),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_863),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_986),
.B(n_983),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1010),
.B(n_560),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_946),
.A2(n_870),
.B(n_882),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_980),
.B(n_1004),
.Y(n_1142)
);

NOR3xp33_ASAP7_75t_L g1143 ( 
.A(n_997),
.B(n_983),
.C(n_986),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_986),
.A2(n_560),
.B1(n_976),
.B2(n_1010),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_980),
.B(n_1004),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_946),
.A2(n_870),
.B(n_882),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1010),
.B(n_560),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_980),
.B(n_1004),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_946),
.A2(n_870),
.B(n_882),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_888),
.A2(n_701),
.B(n_1003),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_975),
.A2(n_743),
.B(n_579),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_980),
.B(n_1004),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1018),
.B(n_1053),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1119),
.A2(n_1152),
.B1(n_1122),
.B2(n_1148),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1025),
.B(n_1142),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1032),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1043),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1038),
.A2(n_1021),
.B(n_1017),
.Y(n_1159)
);

NOR2xp67_ASAP7_75t_L g1160 ( 
.A(n_1034),
.B(n_1036),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_L g1161 ( 
.A(n_1143),
.B(n_1139),
.C(n_1121),
.Y(n_1161)
);

AOI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1115),
.A2(n_1147),
.B(n_1140),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1145),
.B(n_1120),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1060),
.B(n_1031),
.Y(n_1164)
);

INVx6_ASAP7_75t_L g1165 ( 
.A(n_1078),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_1058),
.B(n_1123),
.Y(n_1166)
);

OA22x2_ASAP7_75t_L g1167 ( 
.A1(n_1063),
.A2(n_1096),
.B1(n_1037),
.B2(n_1016),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_1094),
.B2(n_1015),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_1015),
.B2(n_1102),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1012),
.A2(n_1047),
.B(n_1061),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1133),
.A2(n_1023),
.B(n_1035),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1096),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1078),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1098),
.A2(n_1136),
.B1(n_1102),
.B2(n_1116),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1133),
.A2(n_1115),
.B(n_1147),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1098),
.A2(n_1108),
.B1(n_1107),
.B2(n_1116),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1027),
.B(n_1040),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1103),
.Y(n_1178)
);

INVx1_ASAP7_75t_SL g1179 ( 
.A(n_1130),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1014),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1054),
.B(n_1143),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1130),
.B(n_1101),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1028),
.B(n_1077),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1028),
.B(n_1130),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1100),
.Y(n_1185)
);

CKINVDCx6p67_ASAP7_75t_R g1186 ( 
.A(n_1048),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1151),
.A2(n_1097),
.B(n_1135),
.Y(n_1187)
);

OR2x6_ASAP7_75t_L g1188 ( 
.A(n_1048),
.B(n_1109),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_1034),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1107),
.A2(n_1108),
.B(n_1136),
.C(n_1099),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1014),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1067),
.B(n_1051),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1048),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1062),
.B(n_1086),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_1111),
.A2(n_1128),
.B(n_1089),
.C(n_1030),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1100),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1029),
.B(n_1059),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1029),
.B(n_1059),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1050),
.B(n_1065),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1114),
.B(n_1118),
.Y(n_1200)
);

NAND2x1p5_ASAP7_75t_L g1201 ( 
.A(n_1039),
.B(n_1066),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1069),
.A2(n_1088),
.B1(n_1090),
.B2(n_1064),
.Y(n_1202)
);

NAND2x1p5_ASAP7_75t_L g1203 ( 
.A(n_1039),
.B(n_1100),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1091),
.A2(n_1144),
.B1(n_1041),
.B2(n_1089),
.Y(n_1204)
);

NOR2x1_ASAP7_75t_L g1205 ( 
.A(n_1070),
.B(n_1112),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1095),
.A2(n_1113),
.B(n_1125),
.Y(n_1206)
);

BUFx10_ASAP7_75t_L g1207 ( 
.A(n_1068),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1126),
.A2(n_1127),
.B(n_1131),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1081),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1104),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1085),
.A2(n_1072),
.B(n_1075),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1055),
.Y(n_1212)
);

AO21x1_ASAP7_75t_L g1213 ( 
.A1(n_1064),
.A2(n_1084),
.B(n_1082),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_1099),
.B(n_1083),
.C(n_1093),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1138),
.B(n_1118),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1055),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1056),
.B(n_1068),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1069),
.B(n_1137),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1076),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1073),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1079),
.B(n_1124),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1056),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1105),
.A2(n_1132),
.B(n_1110),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1071),
.A2(n_1074),
.B(n_1046),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1137),
.B(n_1052),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1044),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1057),
.A2(n_1020),
.B(n_1045),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1063),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_SL g1229 ( 
.A1(n_1087),
.A2(n_1024),
.B(n_1080),
.C(n_1092),
.Y(n_1229)
);

INVx3_ASAP7_75t_SL g1230 ( 
.A(n_1068),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1068),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1137),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1106),
.A2(n_1129),
.B(n_1149),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1137),
.B(n_1087),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1080),
.B(n_1049),
.Y(n_1235)
);

AOI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1134),
.A2(n_1150),
.B(n_1026),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1080),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1117),
.B(n_1146),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1024),
.A2(n_983),
.B(n_732),
.C(n_1011),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_SL g1240 ( 
.A(n_1141),
.B(n_983),
.C(n_986),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1011),
.B(n_983),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1036),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1036),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1011),
.B(n_1013),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1036),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1036),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1130),
.B(n_1101),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1048),
.B(n_1078),
.Y(n_1248)
);

BUFx3_ASAP7_75t_L g1249 ( 
.A(n_1036),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1123),
.Y(n_1250)
);

OAI21xp33_ASAP7_75t_L g1251 ( 
.A1(n_1011),
.A2(n_705),
.B(n_983),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1143),
.A2(n_983),
.B1(n_986),
.B2(n_732),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1143),
.A2(n_983),
.B1(n_986),
.B2(n_997),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1100),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1036),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1018),
.B(n_1053),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1011),
.B(n_983),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1078),
.Y(n_1258)
);

OA21x2_ASAP7_75t_L g1259 ( 
.A1(n_1030),
.A2(n_1022),
.B(n_1019),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1078),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1038),
.A2(n_1021),
.B(n_1017),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1018),
.B(n_1053),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1036),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_1034),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1011),
.A2(n_560),
.B1(n_1119),
.B2(n_1013),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1036),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1038),
.A2(n_1021),
.B(n_1017),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1018),
.B(n_1053),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1025),
.B(n_981),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1021),
.A2(n_560),
.B(n_1095),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1036),
.Y(n_1271)
);

AOI22x1_ASAP7_75t_L g1272 ( 
.A1(n_1037),
.A2(n_872),
.B1(n_1061),
.B2(n_960),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1036),
.Y(n_1273)
);

OR2x6_ASAP7_75t_L g1274 ( 
.A(n_1048),
.B(n_1078),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1018),
.B(n_1053),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1018),
.B(n_1053),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1011),
.B(n_983),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1025),
.B(n_981),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1100),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1130),
.B(n_1101),
.Y(n_1280)
);

NOR2xp67_ASAP7_75t_L g1281 ( 
.A(n_1034),
.B(n_1036),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1038),
.A2(n_1021),
.B(n_1017),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1130),
.B(n_1101),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1032),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1034),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1025),
.B(n_981),
.Y(n_1286)
);

AND2x4_ASAP7_75t_L g1287 ( 
.A(n_1130),
.B(n_1101),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1038),
.A2(n_1021),
.B(n_1017),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1011),
.A2(n_983),
.B(n_732),
.C(n_1013),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1036),
.Y(n_1290)
);

BUFx4f_ASAP7_75t_SL g1291 ( 
.A(n_1263),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1162),
.B(n_1225),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1161),
.A2(n_1251),
.B1(n_1252),
.B2(n_1277),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1167),
.A2(n_1241),
.B1(n_1257),
.B2(n_1169),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1157),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1164),
.A2(n_1253),
.B1(n_1169),
.B2(n_1199),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1158),
.Y(n_1297)
);

BUFx4f_ASAP7_75t_SL g1298 ( 
.A(n_1189),
.Y(n_1298)
);

CKINVDCx6p67_ASAP7_75t_R g1299 ( 
.A(n_1264),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1192),
.B(n_1244),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1156),
.B(n_1177),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1167),
.A2(n_1204),
.B1(n_1272),
.B2(n_1181),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1165),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1156),
.B(n_1177),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1181),
.A2(n_1214),
.B1(n_1168),
.B2(n_1154),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1223),
.A2(n_1233),
.B(n_1236),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1178),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1210),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1200),
.B(n_1184),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1155),
.A2(n_1168),
.B1(n_1174),
.B2(n_1176),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1155),
.B(n_1289),
.Y(n_1311)
);

AO21x1_ASAP7_75t_L g1312 ( 
.A1(n_1174),
.A2(n_1176),
.B(n_1171),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1265),
.B(n_1269),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1203),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1153),
.B(n_1256),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1265),
.A2(n_1183),
.B1(n_1213),
.B2(n_1171),
.Y(n_1316)
);

INVx6_ASAP7_75t_L g1317 ( 
.A(n_1207),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1245),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1278),
.A2(n_1286),
.B1(n_1268),
.B2(n_1262),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1166),
.Y(n_1320)
);

NOR2xp67_ASAP7_75t_SL g1321 ( 
.A(n_1286),
.B(n_1165),
.Y(n_1321)
);

INVx6_ASAP7_75t_L g1322 ( 
.A(n_1207),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1275),
.A2(n_1276),
.B1(n_1240),
.B2(n_1163),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_1285),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1215),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1209),
.A2(n_1172),
.B1(n_1191),
.B2(n_1193),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1228),
.Y(n_1327)
);

INVx4_ASAP7_75t_SL g1328 ( 
.A(n_1230),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1284),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1222),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1165),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1219),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1264),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1220),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1220),
.Y(n_1335)
);

CKINVDCx11_ASAP7_75t_R g1336 ( 
.A(n_1250),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1250),
.B(n_1179),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1172),
.Y(n_1338)
);

INVx8_ASAP7_75t_L g1339 ( 
.A(n_1188),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1191),
.A2(n_1274),
.B1(n_1248),
.B2(n_1188),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1221),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1234),
.B(n_1232),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1186),
.A2(n_1160),
.B1(n_1281),
.B2(n_1248),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1235),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1202),
.A2(n_1248),
.B1(n_1274),
.B2(n_1175),
.Y(n_1345)
);

AO21x1_ASAP7_75t_L g1346 ( 
.A1(n_1175),
.A2(n_1202),
.B(n_1239),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1179),
.B(n_1283),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1218),
.B(n_1195),
.Y(n_1348)
);

OAI21xp33_ASAP7_75t_L g1349 ( 
.A1(n_1190),
.A2(n_1249),
.B(n_1246),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1259),
.A2(n_1280),
.B1(n_1283),
.B2(n_1247),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1271),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1242),
.B(n_1273),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1243),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1212),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1259),
.Y(n_1355)
);

BUFx12f_ASAP7_75t_L g1356 ( 
.A(n_1290),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1185),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1217),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1274),
.A2(n_1258),
.B1(n_1260),
.B2(n_1173),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1217),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1182),
.A2(n_1247),
.B1(n_1280),
.B2(n_1287),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1196),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1182),
.A2(n_1287),
.B1(n_1218),
.B2(n_1255),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1197),
.A2(n_1180),
.B1(n_1266),
.B2(n_1201),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1201),
.A2(n_1258),
.B1(n_1173),
.B2(n_1260),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1198),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1237),
.B(n_1216),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1170),
.A2(n_1270),
.B1(n_1288),
.B2(n_1261),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1224),
.A2(n_1226),
.B1(n_1288),
.B2(n_1159),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1254),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1224),
.A2(n_1282),
.B1(n_1267),
.B2(n_1261),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1238),
.Y(n_1372)
);

CKINVDCx11_ASAP7_75t_R g1373 ( 
.A(n_1254),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1231),
.A2(n_1205),
.B1(n_1187),
.B2(n_1206),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1279),
.B(n_1267),
.Y(n_1375)
);

AO21x2_ASAP7_75t_L g1376 ( 
.A1(n_1227),
.A2(n_1208),
.B(n_1238),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_1227),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1229),
.A2(n_983),
.B1(n_986),
.B2(n_1143),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1253),
.A2(n_745),
.B1(n_986),
.B2(n_1011),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1167),
.A2(n_745),
.B1(n_986),
.B2(n_732),
.Y(n_1380)
);

BUFx2_ASAP7_75t_R g1381 ( 
.A(n_1285),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1157),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1223),
.A2(n_1233),
.B(n_1236),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1161),
.A2(n_983),
.B1(n_986),
.B2(n_1143),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1218),
.B(n_1168),
.Y(n_1385)
);

BUFx8_ASAP7_75t_SL g1386 ( 
.A(n_1189),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1162),
.B(n_1115),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1223),
.A2(n_1233),
.B(n_1236),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1161),
.B(n_368),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1162),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1192),
.B(n_1011),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_1185),
.Y(n_1392)
);

CKINVDCx9p33_ASAP7_75t_R g1393 ( 
.A(n_1194),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1170),
.A2(n_1211),
.B(n_1159),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1166),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1162),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1250),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1166),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1223),
.A2(n_1233),
.B(n_1236),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1157),
.Y(n_1400)
);

INVx4_ASAP7_75t_SL g1401 ( 
.A(n_1375),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1348),
.B(n_1385),
.Y(n_1402)
);

INVxp33_ASAP7_75t_L g1403 ( 
.A(n_1315),
.Y(n_1403)
);

AO21x1_ASAP7_75t_SL g1404 ( 
.A1(n_1311),
.A2(n_1302),
.B(n_1316),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1342),
.B(n_1313),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1348),
.B(n_1385),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1372),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1372),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1342),
.B(n_1313),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1375),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1355),
.Y(n_1411)
);

OR2x6_ASAP7_75t_L g1412 ( 
.A(n_1339),
.B(n_1312),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1391),
.B(n_1379),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1344),
.B(n_1301),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1292),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1301),
.B(n_1304),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1292),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1390),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1304),
.B(n_1344),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1338),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1371),
.A2(n_1346),
.B(n_1369),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1309),
.B(n_1310),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1294),
.A2(n_1293),
.B1(n_1380),
.B2(n_1389),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1390),
.Y(n_1424)
);

CKINVDCx6p67_ASAP7_75t_R g1425 ( 
.A(n_1336),
.Y(n_1425)
);

AOI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1321),
.A2(n_1374),
.B(n_1306),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1396),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1384),
.A2(n_1378),
.B(n_1300),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1394),
.Y(n_1429)
);

CKINVDCx16_ASAP7_75t_R g1430 ( 
.A(n_1333),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1341),
.B(n_1305),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1346),
.Y(n_1432)
);

AOI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1321),
.A2(n_1383),
.B(n_1306),
.Y(n_1433)
);

AO21x1_ASAP7_75t_SL g1434 ( 
.A1(n_1296),
.A2(n_1319),
.B(n_1323),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1398),
.B(n_1387),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1377),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1309),
.B(n_1367),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1387),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1387),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1330),
.Y(n_1440)
);

BUFx2_ASAP7_75t_L g1441 ( 
.A(n_1377),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1338),
.Y(n_1442)
);

AOI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1383),
.A2(n_1388),
.B(n_1399),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1376),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1334),
.B(n_1335),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1325),
.B(n_1358),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1320),
.B(n_1395),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1325),
.B(n_1358),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1295),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1297),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1307),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1308),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1340),
.B(n_1365),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_1397),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1329),
.A2(n_1400),
.B(n_1382),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1337),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1366),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1366),
.Y(n_1458)
);

AO21x2_ASAP7_75t_L g1459 ( 
.A1(n_1332),
.A2(n_1368),
.B(n_1360),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1317),
.Y(n_1460)
);

INVx4_ASAP7_75t_L g1461 ( 
.A(n_1328),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1353),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1345),
.A2(n_1349),
.B1(n_1347),
.B2(n_1363),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1336),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1317),
.Y(n_1465)
);

NAND2x1_ASAP7_75t_L g1466 ( 
.A(n_1350),
.B(n_1314),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1393),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1354),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1317),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1459),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1411),
.B(n_1347),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1427),
.B(n_1362),
.Y(n_1472)
);

OR2x2_ASAP7_75t_SL g1473 ( 
.A(n_1430),
.B(n_1402),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1459),
.Y(n_1474)
);

AOI222xp33_ASAP7_75t_L g1475 ( 
.A1(n_1428),
.A2(n_1298),
.B1(n_1326),
.B2(n_1291),
.C1(n_1343),
.C2(n_1352),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1429),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1402),
.B(n_1406),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1459),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1405),
.B(n_1370),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1435),
.Y(n_1480)
);

NOR2x1p5_ASAP7_75t_L g1481 ( 
.A(n_1461),
.B(n_1299),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1406),
.B(n_1364),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1423),
.A2(n_1333),
.B1(n_1359),
.B2(n_1327),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1409),
.B(n_1392),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1401),
.B(n_1328),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1432),
.B(n_1351),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1432),
.B(n_1351),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1409),
.B(n_1392),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1444),
.B(n_1331),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1416),
.B(n_1303),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1455),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1418),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1423),
.A2(n_1356),
.B1(n_1361),
.B2(n_1327),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1418),
.B(n_1392),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1455),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1435),
.B(n_1303),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1413),
.A2(n_1356),
.B1(n_1318),
.B2(n_1299),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1424),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1455),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1434),
.A2(n_1318),
.B1(n_1386),
.B2(n_1324),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1463),
.A2(n_1403),
.B1(n_1422),
.B2(n_1431),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1449),
.Y(n_1502)
);

INVx5_ASAP7_75t_L g1503 ( 
.A(n_1412),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1430),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1401),
.B(n_1328),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1420),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1416),
.B(n_1438),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1439),
.B(n_1357),
.Y(n_1508)
);

AOI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1443),
.A2(n_1426),
.B(n_1433),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1407),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1507),
.B(n_1410),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1507),
.B(n_1410),
.Y(n_1512)
);

AND2x2_ASAP7_75t_SL g1513 ( 
.A(n_1485),
.B(n_1436),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1477),
.B(n_1480),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1506),
.B(n_1456),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1500),
.B(n_1467),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_SL g1517 ( 
.A(n_1485),
.B(n_1461),
.Y(n_1517)
);

OAI21xp33_ASAP7_75t_L g1518 ( 
.A1(n_1483),
.A2(n_1431),
.B(n_1422),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1477),
.B(n_1415),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1476),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1477),
.B(n_1442),
.Y(n_1521)
);

OAI21xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1483),
.A2(n_1436),
.B(n_1441),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_L g1523 ( 
.A(n_1475),
.B(n_1454),
.C(n_1462),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1480),
.B(n_1419),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1509),
.A2(n_1495),
.B(n_1491),
.Y(n_1525)
);

NAND4xp25_ASAP7_75t_L g1526 ( 
.A(n_1475),
.B(n_1493),
.C(n_1500),
.D(n_1501),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1493),
.A2(n_1441),
.B1(n_1425),
.B2(n_1447),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1504),
.B(n_1464),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1506),
.B(n_1419),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_SL g1530 ( 
.A1(n_1501),
.A2(n_1467),
.B(n_1434),
.Y(n_1530)
);

OAI221xp5_ASAP7_75t_SL g1531 ( 
.A1(n_1497),
.A2(n_1453),
.B1(n_1412),
.B2(n_1447),
.C(n_1425),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1484),
.B(n_1488),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1471),
.B(n_1479),
.Y(n_1533)
);

OAI21xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1481),
.A2(n_1412),
.B(n_1461),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1497),
.A2(n_1404),
.B1(n_1453),
.B2(n_1412),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1471),
.B(n_1417),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1482),
.A2(n_1404),
.B1(n_1453),
.B2(n_1412),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1490),
.B(n_1468),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1482),
.A2(n_1453),
.B1(n_1466),
.B2(n_1458),
.Y(n_1539)
);

NAND3xp33_ASAP7_75t_L g1540 ( 
.A(n_1470),
.B(n_1421),
.C(n_1445),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1502),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1482),
.A2(n_1453),
.B1(n_1504),
.B2(n_1466),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1471),
.B(n_1437),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1470),
.B(n_1421),
.C(n_1445),
.Y(n_1544)
);

AOI211xp5_ASAP7_75t_L g1545 ( 
.A1(n_1474),
.A2(n_1451),
.B(n_1450),
.C(n_1452),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1496),
.B(n_1324),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1510),
.B(n_1440),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1479),
.B(n_1324),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1510),
.B(n_1440),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1479),
.B(n_1446),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1508),
.B(n_1494),
.Y(n_1551)
);

OAI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1486),
.A2(n_1457),
.B1(n_1458),
.B2(n_1465),
.C(n_1469),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1486),
.B(n_1448),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1486),
.B(n_1487),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1502),
.Y(n_1555)
);

OAI221xp5_ASAP7_75t_SL g1556 ( 
.A1(n_1474),
.A2(n_1414),
.B1(n_1457),
.B2(n_1458),
.C(n_1450),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1510),
.B(n_1408),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1487),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1472),
.B(n_1414),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1514),
.B(n_1491),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1514),
.B(n_1473),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1551),
.B(n_1503),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1519),
.B(n_1495),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1554),
.B(n_1473),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1532),
.B(n_1503),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1520),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1521),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1521),
.B(n_1473),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1532),
.B(n_1503),
.Y(n_1569)
);

BUFx2_ASAP7_75t_SL g1570 ( 
.A(n_1516),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1541),
.Y(n_1571)
);

AND2x4_ASAP7_75t_SL g1572 ( 
.A(n_1519),
.B(n_1485),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1541),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1558),
.B(n_1489),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1533),
.B(n_1503),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1555),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1555),
.Y(n_1577)
);

NAND2x1_ASAP7_75t_SL g1578 ( 
.A(n_1536),
.B(n_1478),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1525),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1545),
.B(n_1499),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1528),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1499),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1547),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1547),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1529),
.B(n_1492),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1549),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1524),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1549),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1557),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1525),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1529),
.B(n_1498),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1571),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1571),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1579),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1578),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1579),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1574),
.B(n_1515),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1575),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1588),
.B(n_1543),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1575),
.B(n_1543),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1575),
.B(n_1511),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1575),
.B(n_1511),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1579),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1573),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1573),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1590),
.Y(n_1606)
);

OAI32xp33_ASAP7_75t_L g1607 ( 
.A1(n_1580),
.A2(n_1526),
.A3(n_1518),
.B1(n_1523),
.B2(n_1540),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1576),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1588),
.B(n_1538),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1590),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1574),
.B(n_1540),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1590),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1576),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1561),
.B(n_1544),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1577),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1577),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1565),
.B(n_1512),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1565),
.B(n_1512),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1565),
.B(n_1478),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1567),
.B(n_1544),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1583),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1580),
.B(n_1525),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1583),
.B(n_1550),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_SL g1624 ( 
.A1(n_1570),
.A2(n_1527),
.B1(n_1548),
.B2(n_1505),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1565),
.B(n_1536),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1584),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1584),
.B(n_1553),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1586),
.Y(n_1628)
);

OAI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1561),
.A2(n_1526),
.B1(n_1522),
.B2(n_1530),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1566),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1569),
.B(n_1513),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1560),
.B(n_1559),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1594),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1631),
.B(n_1569),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1599),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1620),
.B(n_1582),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1609),
.B(n_1568),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1609),
.B(n_1568),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1592),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1620),
.B(n_1582),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1592),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1614),
.B(n_1560),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1593),
.Y(n_1643)
);

OR2x2_ASAP7_75t_SL g1644 ( 
.A(n_1614),
.B(n_1564),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1629),
.A2(n_1530),
.B1(n_1522),
.B2(n_1517),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1631),
.B(n_1569),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1629),
.B(n_1564),
.Y(n_1649)
);

NAND2x2_ASAP7_75t_L g1650 ( 
.A(n_1595),
.B(n_1481),
.Y(n_1650)
);

AOI21xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1607),
.A2(n_1581),
.B(n_1518),
.Y(n_1651)
);

NAND2xp67_ASAP7_75t_L g1652 ( 
.A(n_1631),
.B(n_1572),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1600),
.B(n_1569),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1523),
.C(n_1531),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1598),
.A2(n_1570),
.B1(n_1513),
.B2(n_1535),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1594),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1597),
.B(n_1585),
.Y(n_1657)
);

AOI222xp33_ASAP7_75t_L g1658 ( 
.A1(n_1607),
.A2(n_1527),
.B1(n_1542),
.B2(n_1537),
.C1(n_1513),
.C2(n_1539),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1594),
.Y(n_1659)
);

OAI21xp33_ASAP7_75t_L g1660 ( 
.A1(n_1611),
.A2(n_1556),
.B(n_1578),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1600),
.B(n_1562),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1611),
.B(n_1599),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1632),
.B(n_1597),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1624),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1596),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1600),
.B(n_1562),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1632),
.B(n_1563),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1627),
.B(n_1546),
.Y(n_1668)
);

NOR2x1_ASAP7_75t_L g1669 ( 
.A(n_1622),
.B(n_1589),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1627),
.B(n_1585),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1596),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1593),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1598),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1596),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1622),
.B(n_1563),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1601),
.B(n_1591),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1649),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1639),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1641),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1651),
.B(n_1668),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1643),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1644),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1672),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1647),
.A2(n_1598),
.B1(n_1595),
.B2(n_1619),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1663),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1668),
.B(n_1601),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1633),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1664),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1662),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1633),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1673),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1673),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1656),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1636),
.B(n_1601),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1634),
.B(n_1595),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1634),
.B(n_1625),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1663),
.B(n_1621),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1648),
.B(n_1625),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1656),
.Y(n_1700)
);

INVx3_ASAP7_75t_SL g1701 ( 
.A(n_1636),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1659),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1659),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1648),
.B(n_1625),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1665),
.A2(n_1674),
.B(n_1671),
.Y(n_1705)
);

AOI222xp33_ASAP7_75t_L g1706 ( 
.A1(n_1654),
.A2(n_1619),
.B1(n_1628),
.B2(n_1626),
.C1(n_1621),
.C2(n_1602),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1665),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1653),
.B(n_1598),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1637),
.B(n_1386),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1658),
.A2(n_1660),
.B1(n_1650),
.B2(n_1638),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1640),
.Y(n_1711)
);

NOR2x1_ASAP7_75t_L g1712 ( 
.A(n_1640),
.B(n_1604),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1696),
.B(n_1698),
.Y(n_1713)
);

OAI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1680),
.A2(n_1677),
.B1(n_1682),
.B2(n_1710),
.C(n_1688),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1684),
.A2(n_1655),
.B1(n_1624),
.B2(n_1650),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1685),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1696),
.B(n_1653),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1699),
.A2(n_1662),
.B1(n_1635),
.B2(n_1676),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1701),
.B(n_1670),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1701),
.B(n_1645),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1698),
.B(n_1661),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_R g1722 ( 
.A(n_1701),
.B(n_1381),
.Y(n_1722)
);

OAI21xp33_ASAP7_75t_L g1723 ( 
.A1(n_1706),
.A2(n_1642),
.B(n_1646),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1689),
.B(n_1657),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1678),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1695),
.B(n_1661),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1695),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1711),
.B(n_1642),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1695),
.A2(n_1517),
.B1(n_1534),
.B2(n_1666),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1678),
.Y(n_1730)
);

AOI32xp33_ASAP7_75t_L g1731 ( 
.A1(n_1699),
.A2(n_1666),
.A3(n_1619),
.B1(n_1617),
.B2(n_1618),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1679),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1679),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1712),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1681),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1709),
.B(n_1652),
.Y(n_1736)
);

NAND2x1p5_ASAP7_75t_L g1737 ( 
.A(n_1712),
.B(n_1461),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1686),
.B(n_1667),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1714),
.A2(n_1694),
.B1(n_1695),
.B2(n_1704),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1722),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1713),
.B(n_1704),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1719),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1719),
.Y(n_1743)
);

NAND2x1_ASAP7_75t_L g1744 ( 
.A(n_1726),
.B(n_1691),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1726),
.B(n_1708),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1727),
.B(n_1692),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1714),
.B(n_1697),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1737),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1717),
.B(n_1708),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1736),
.B(n_1716),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1737),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1734),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1725),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1724),
.B(n_1697),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1728),
.B(n_1681),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1720),
.B(n_1683),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1730),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1720),
.B(n_1683),
.Y(n_1758)
);

AOI211xp5_ASAP7_75t_L g1759 ( 
.A1(n_1747),
.A2(n_1715),
.B(n_1718),
.C(n_1723),
.Y(n_1759)
);

A2O1A1Ixp33_ASAP7_75t_L g1760 ( 
.A1(n_1739),
.A2(n_1738),
.B(n_1731),
.C(n_1728),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1740),
.B(n_1729),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1754),
.Y(n_1762)
);

AOI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1742),
.A2(n_1735),
.B1(n_1733),
.B2(n_1732),
.C(n_1721),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1750),
.A2(n_1691),
.B(n_1690),
.Y(n_1764)
);

AOI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1743),
.A2(n_1692),
.B(n_1687),
.C(n_1690),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1745),
.A2(n_1692),
.B1(n_1693),
.B2(n_1687),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1745),
.A2(n_1693),
.B1(n_1702),
.B2(n_1700),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1744),
.A2(n_1705),
.B(n_1702),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1746),
.B(n_1700),
.Y(n_1769)
);

OAI211xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1756),
.A2(n_1707),
.B(n_1703),
.C(n_1675),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1762),
.B(n_1758),
.Y(n_1771)
);

NAND4xp25_ASAP7_75t_L g1772 ( 
.A(n_1759),
.B(n_1752),
.C(n_1755),
.D(n_1753),
.Y(n_1772)
);

OAI211xp5_ASAP7_75t_L g1773 ( 
.A1(n_1760),
.A2(n_1744),
.B(n_1755),
.C(n_1757),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1765),
.B(n_1746),
.C(n_1754),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1769),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1763),
.B(n_1746),
.Y(n_1776)
);

AOI211x1_ASAP7_75t_L g1777 ( 
.A1(n_1761),
.A2(n_1749),
.B(n_1741),
.C(n_1628),
.Y(n_1777)
);

AOI22x1_ASAP7_75t_SL g1778 ( 
.A1(n_1764),
.A2(n_1751),
.B1(n_1748),
.B2(n_1707),
.Y(n_1778)
);

NOR2x1_ASAP7_75t_L g1779 ( 
.A(n_1770),
.B(n_1748),
.Y(n_1779)
);

NOR3xp33_ASAP7_75t_L g1780 ( 
.A(n_1766),
.B(n_1751),
.C(n_1741),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1767),
.B(n_1749),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1768),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_SL g1783 ( 
.A(n_1773),
.B(n_1707),
.C(n_1675),
.Y(n_1783)
);

AOI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1772),
.A2(n_1705),
.B(n_1703),
.C(n_1674),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1780),
.B(n_1667),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1776),
.B(n_1671),
.C(n_1552),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1775),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1774),
.Y(n_1788)
);

NOR4xp25_ASAP7_75t_L g1789 ( 
.A(n_1782),
.B(n_1771),
.C(n_1781),
.D(n_1778),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1785),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1788),
.B(n_1777),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1789),
.B(n_1779),
.Y(n_1792)
);

CKINVDCx16_ASAP7_75t_R g1793 ( 
.A(n_1783),
.Y(n_1793)
);

BUFx2_ASAP7_75t_L g1794 ( 
.A(n_1787),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1784),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1786),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1792),
.B(n_1703),
.Y(n_1797)
);

XNOR2xp5_ASAP7_75t_L g1798 ( 
.A(n_1792),
.B(n_1703),
.Y(n_1798)
);

XOR2xp5_ASAP7_75t_L g1799 ( 
.A(n_1793),
.B(n_1602),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1796),
.A2(n_1317),
.B1(n_1322),
.B2(n_1626),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1790),
.A2(n_1322),
.B1(n_1603),
.B2(n_1606),
.Y(n_1801)
);

NAND4xp75_ASAP7_75t_L g1802 ( 
.A(n_1791),
.B(n_1534),
.C(n_1603),
.D(n_1610),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1799),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1798),
.B(n_1794),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1797),
.Y(n_1805)
);

AOI22x1_ASAP7_75t_L g1806 ( 
.A1(n_1803),
.A2(n_1795),
.B1(n_1800),
.B2(n_1802),
.Y(n_1806)
);

OAI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1806),
.A2(n_1795),
.B1(n_1803),
.B2(n_1805),
.C(n_1804),
.Y(n_1807)
);

OAI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1807),
.A2(n_1801),
.B1(n_1610),
.B2(n_1603),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1807),
.A2(n_1606),
.B1(n_1610),
.B2(n_1612),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1808),
.A2(n_1606),
.B1(n_1612),
.B2(n_1373),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1809),
.Y(n_1811)
);

AOI222xp33_ASAP7_75t_L g1812 ( 
.A1(n_1811),
.A2(n_1612),
.B1(n_1605),
.B2(n_1608),
.C1(n_1604),
.C2(n_1616),
.Y(n_1812)
);

AOI21xp33_ASAP7_75t_SL g1813 ( 
.A1(n_1810),
.A2(n_1465),
.B(n_1460),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1813),
.A2(n_1812),
.B(n_1617),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1814),
.A2(n_1373),
.B1(n_1630),
.B2(n_1608),
.Y(n_1815)
);

OAI221xp5_ASAP7_75t_R g1816 ( 
.A1(n_1815),
.A2(n_1630),
.B1(n_1328),
.B2(n_1616),
.C(n_1615),
.Y(n_1816)
);

AOI211xp5_ASAP7_75t_L g1817 ( 
.A1(n_1816),
.A2(n_1615),
.B(n_1605),
.C(n_1613),
.Y(n_1817)
);


endmodule