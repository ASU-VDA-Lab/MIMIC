module fake_netlist_1_8555_n_20 (n_1, n_2, n_4, n_3, n_5, n_0, n_20);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_6;
wire n_7;
INVx1_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_5), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_0), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_4), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_1), .Y(n_10) );
OAI21x1_ASAP7_75t_L g11 ( .A1(n_7), .A2(n_0), .B(n_1), .Y(n_11) );
OAI22xp33_ASAP7_75t_L g12 ( .A1(n_8), .A2(n_2), .B1(n_3), .B2(n_6), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_13), .B(n_8), .Y(n_14) );
INVx4_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
A2O1A1Ixp33_ASAP7_75t_L g16 ( .A1(n_14), .A2(n_11), .B(n_10), .C(n_12), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_15), .B(n_11), .Y(n_17) );
O2A1O1Ixp33_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_2), .B(n_15), .C(n_17), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
XOR2xp5_ASAP7_75t_L g20 ( .A(n_19), .B(n_15), .Y(n_20) );
endmodule