module real_aes_6809_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_119;
wire n_504;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g178 ( .A1(n_0), .A2(n_179), .B(n_180), .C(n_184), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_1), .B(n_173), .Y(n_186) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g126 ( .A(n_2), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_3), .B(n_158), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_4), .A2(n_167), .B(n_479), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_5), .A2(n_147), .B(n_164), .C(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_6), .A2(n_167), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_7), .B(n_173), .Y(n_485) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_8), .A2(n_139), .B(n_261), .Y(n_260) );
AND2x6_ASAP7_75t_L g164 ( .A(n_9), .B(n_165), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_10), .A2(n_147), .B(n_164), .C(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g576 ( .A(n_11), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_39), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_13), .B(n_183), .Y(n_525) );
INVx1_ASAP7_75t_L g144 ( .A(n_14), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_15), .B(n_158), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_16), .A2(n_159), .B(n_534), .C(n_536), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_17), .B(n_173), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_18), .B(n_201), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_19), .A2(n_147), .B(n_193), .C(n_200), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g542 ( .A1(n_20), .A2(n_182), .B(n_235), .C(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_21), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_22), .B(n_183), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_23), .B(n_183), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_24), .Y(n_503) );
INVx1_ASAP7_75t_L g473 ( .A(n_25), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_26), .A2(n_147), .B(n_200), .C(n_264), .Y(n_263) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_27), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_28), .Y(n_521) );
INVx1_ASAP7_75t_L g497 ( .A(n_29), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_30), .A2(n_167), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g149 ( .A(n_31), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_32), .A2(n_162), .B(n_216), .C(n_217), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_33), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_34), .A2(n_182), .B(n_482), .C(n_484), .Y(n_481) );
INVxp67_ASAP7_75t_L g498 ( .A(n_35), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_36), .B(n_266), .Y(n_265) );
CKINVDCx14_ASAP7_75t_R g480 ( .A(n_37), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_38), .A2(n_147), .B(n_200), .C(n_472), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_40), .A2(n_184), .B(n_574), .C(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_41), .B(n_191), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_42), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_43), .B(n_158), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_44), .B(n_167), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_45), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_46), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_47), .A2(n_104), .B1(n_115), .B2(n_730), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_48), .A2(n_162), .B(n_216), .C(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g181 ( .A(n_49), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_50), .A2(n_128), .B1(n_442), .B2(n_443), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_50), .Y(n_442) );
INVx1_ASAP7_75t_L g245 ( .A(n_51), .Y(n_245) );
INVx1_ASAP7_75t_L g541 ( .A(n_52), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_53), .B(n_167), .Y(n_242) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_54), .A2(n_72), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_54), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_55), .Y(n_205) );
AOI222xp33_ASAP7_75t_SL g448 ( .A1(n_56), .A2(n_449), .B1(n_455), .B2(n_724), .C1(n_725), .C2(n_726), .Y(n_448) );
CKINVDCx14_ASAP7_75t_R g572 ( .A(n_57), .Y(n_572) );
INVx1_ASAP7_75t_L g165 ( .A(n_58), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_59), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_60), .B(n_173), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_61), .A2(n_154), .B(n_199), .C(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_62), .A2(n_71), .B1(n_453), .B2(n_454), .Y(n_452) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_62), .Y(n_453) );
INVx1_ASAP7_75t_L g143 ( .A(n_63), .Y(n_143) );
INVx1_ASAP7_75t_SL g483 ( .A(n_64), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_65), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_66), .B(n_158), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_67), .B(n_173), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_68), .B(n_159), .Y(n_232) );
INVx1_ASAP7_75t_L g506 ( .A(n_69), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g176 ( .A(n_70), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_71), .Y(n_454) );
INVx1_ASAP7_75t_L g131 ( .A(n_72), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_73), .B(n_195), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_74), .A2(n_147), .B(n_152), .C(n_162), .Y(n_146) );
CKINVDCx16_ASAP7_75t_R g254 ( .A(n_75), .Y(n_254) );
INVx1_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_77), .A2(n_167), .B(n_571), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_78), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_79), .A2(n_167), .B(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_80), .A2(n_191), .B(n_493), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_81), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_82), .A2(n_450), .B1(n_451), .B2(n_452), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_82), .Y(n_450) );
INVx1_ASAP7_75t_L g532 ( .A(n_83), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_84), .B(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_85), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_86), .A2(n_167), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g535 ( .A(n_87), .Y(n_535) );
INVx2_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
INVx1_ASAP7_75t_L g524 ( .A(n_89), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_90), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_91), .B(n_183), .Y(n_233) );
INVx2_ASAP7_75t_L g109 ( .A(n_92), .Y(n_109) );
OR2x2_ASAP7_75t_L g123 ( .A(n_92), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g459 ( .A(n_92), .B(n_125), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_93), .A2(n_147), .B(n_162), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_94), .B(n_167), .Y(n_214) );
INVx1_ASAP7_75t_L g218 ( .A(n_95), .Y(n_218) );
INVxp67_ASAP7_75t_L g257 ( .A(n_96), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_97), .B(n_139), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g153 ( .A(n_99), .Y(n_153) );
INVx1_ASAP7_75t_L g228 ( .A(n_100), .Y(n_228) );
INVx2_ASAP7_75t_L g544 ( .A(n_101), .Y(n_544) );
AND2x2_ASAP7_75t_L g247 ( .A(n_102), .B(n_203), .Y(n_247) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_106), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_113), .Y(n_107) );
OR2x2_ASAP7_75t_L g723 ( .A(n_109), .B(n_125), .Y(n_723) );
NOR2x2_ASAP7_75t_L g724 ( .A(n_109), .B(n_124), .Y(n_724) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g125 ( .A(n_114), .B(n_126), .Y(n_125) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_447), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_117), .B(n_444), .C(n_448), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_127), .B(n_444), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_123), .Y(n_446) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g443 ( .A(n_128), .Y(n_443) );
XNOR2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_132), .Y(n_128) );
INVx1_ASAP7_75t_L g456 ( .A(n_132), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_132), .A2(n_461), .B1(n_727), .B2(n_728), .Y(n_726) );
OR3x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_350), .C(n_399), .Y(n_132) );
NAND5xp2_ASAP7_75t_L g133 ( .A(n_134), .B(n_284), .C(n_313), .D(n_321), .E(n_336), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_207), .B(n_223), .C(n_268), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_187), .Y(n_135) );
AND2x2_ASAP7_75t_L g279 ( .A(n_136), .B(n_276), .Y(n_279) );
AND2x2_ASAP7_75t_L g312 ( .A(n_136), .B(n_188), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_136), .B(n_211), .Y(n_405) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_172), .Y(n_136) );
INVx2_ASAP7_75t_L g210 ( .A(n_137), .Y(n_210) );
BUFx2_ASAP7_75t_L g379 ( .A(n_137), .Y(n_379) );
AO21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_145), .B(n_170), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_138), .B(n_171), .Y(n_170) );
INVx3_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_138), .B(n_222), .Y(n_221) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_138), .A2(n_227), .B(n_237), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_138), .B(n_476), .Y(n_475) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_138), .A2(n_502), .B(n_509), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_138), .B(n_527), .Y(n_526) );
INVx4_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_139), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_139), .A2(n_262), .B(n_263), .Y(n_261) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g239 ( .A(n_140), .Y(n_239) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g203 ( .A(n_141), .B(n_142), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_166), .Y(n_145) );
INVx5_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
BUFx3_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
INVx1_ASAP7_75t_L g236 ( .A(n_149), .Y(n_236) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_151), .Y(n_156) );
INVx3_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
AND2x2_ASAP7_75t_L g168 ( .A(n_151), .B(n_169), .Y(n_168) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
INVx1_ASAP7_75t_L g266 ( .A(n_151), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_157), .C(n_160), .Y(n_152) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
OAI22xp33_ASAP7_75t_L g496 ( .A1(n_155), .A2(n_158), .B1(n_497), .B2(n_498), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_155), .B(n_535), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_155), .B(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
INVx2_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_158), .B(n_257), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_158), .A2(n_198), .B(n_473), .C(n_474), .Y(n_472) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_159), .B(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g484 ( .A(n_161), .Y(n_484) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_SL g175 ( .A1(n_163), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_163), .A2(n_177), .B(n_254), .C(n_255), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_163), .A2(n_177), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_163), .A2(n_177), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_163), .A2(n_177), .B(n_532), .C(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g540 ( .A1(n_163), .A2(n_177), .B(n_541), .C(n_542), .Y(n_540) );
O2A1O1Ixp33_ASAP7_75t_SL g571 ( .A1(n_163), .A2(n_177), .B(n_572), .C(n_573), .Y(n_571) );
INVx4_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g167 ( .A(n_164), .B(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
NAND2x1p5_ASAP7_75t_L g229 ( .A(n_164), .B(n_168), .Y(n_229) );
BUFx2_ASAP7_75t_L g191 ( .A(n_167), .Y(n_191) );
INVx1_ASAP7_75t_L g199 ( .A(n_169), .Y(n_199) );
AND2x2_ASAP7_75t_L g187 ( .A(n_172), .B(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g277 ( .A(n_172), .Y(n_277) );
AND2x2_ASAP7_75t_L g363 ( .A(n_172), .B(n_276), .Y(n_363) );
AND2x2_ASAP7_75t_L g418 ( .A(n_172), .B(n_210), .Y(n_418) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_186), .Y(n_172) );
INVx2_ASAP7_75t_L g216 ( .A(n_177), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_182), .B(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g574 ( .A(n_183), .Y(n_574) );
INVx2_ASAP7_75t_L g508 ( .A(n_184), .Y(n_508) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_185), .Y(n_220) );
INVx1_ASAP7_75t_L g536 ( .A(n_185), .Y(n_536) );
INVx1_ASAP7_75t_L g335 ( .A(n_187), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_187), .B(n_211), .Y(n_382) );
INVx5_ASAP7_75t_L g276 ( .A(n_188), .Y(n_276) );
AND2x4_ASAP7_75t_L g297 ( .A(n_188), .B(n_277), .Y(n_297) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_188), .Y(n_319) );
AND2x2_ASAP7_75t_L g394 ( .A(n_188), .B(n_379), .Y(n_394) );
AND2x2_ASAP7_75t_L g397 ( .A(n_188), .B(n_212), .Y(n_397) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_204), .Y(n_188) );
AOI21xp5_ASAP7_75t_SL g189 ( .A1(n_190), .A2(n_192), .B(n_201), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_196), .B(n_198), .Y(n_193) );
INVx2_ASAP7_75t_L g197 ( .A(n_195), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_197), .A2(n_218), .B(n_219), .C(n_220), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_197), .A2(n_220), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_197), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
O2A1O1Ixp5_ASAP7_75t_L g523 ( .A1(n_197), .A2(n_508), .B(n_524), .C(n_525), .Y(n_523) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_199), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_202), .B(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g206 ( .A(n_203), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_203), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_203), .A2(n_242), .B(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_203), .A2(n_229), .B(n_470), .C(n_471), .Y(n_469) );
OA21x2_ASAP7_75t_L g569 ( .A1(n_203), .A2(n_570), .B(n_577), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_206), .A2(n_520), .B(n_526), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_207), .B(n_277), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_207), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
AND2x2_ASAP7_75t_L g302 ( .A(n_209), .B(n_277), .Y(n_302) );
AND2x2_ASAP7_75t_L g320 ( .A(n_209), .B(n_212), .Y(n_320) );
INVx1_ASAP7_75t_L g340 ( .A(n_209), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_209), .B(n_276), .Y(n_385) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_209), .Y(n_427) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_210), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_211), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_211), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_211), .A2(n_272), .B(n_333), .C(n_335), .Y(n_332) );
AND2x2_ASAP7_75t_L g339 ( .A(n_211), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g348 ( .A(n_211), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g352 ( .A(n_211), .B(n_276), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_211), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g367 ( .A(n_211), .B(n_277), .Y(n_367) );
AND2x2_ASAP7_75t_L g417 ( .A(n_211), .B(n_418), .Y(n_417) );
INVx5_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
BUFx2_ASAP7_75t_L g281 ( .A(n_212), .Y(n_281) );
AND2x2_ASAP7_75t_L g322 ( .A(n_212), .B(n_275), .Y(n_322) );
AND2x2_ASAP7_75t_L g334 ( .A(n_212), .B(n_309), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_212), .B(n_363), .Y(n_381) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_221), .Y(n_212) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_248), .Y(n_223) );
INVx1_ASAP7_75t_L g270 ( .A(n_224), .Y(n_270) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_240), .Y(n_224) );
OR2x2_ASAP7_75t_L g272 ( .A(n_225), .B(n_240), .Y(n_272) );
NAND3xp33_ASAP7_75t_L g278 ( .A(n_225), .B(n_279), .C(n_280), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_225), .B(n_250), .Y(n_289) );
OR2x2_ASAP7_75t_L g304 ( .A(n_225), .B(n_292), .Y(n_304) );
AND2x2_ASAP7_75t_L g310 ( .A(n_225), .B(n_259), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_225), .B(n_441), .Y(n_440) );
INVx5_ASAP7_75t_SL g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_226), .B(n_250), .Y(n_307) );
AND2x2_ASAP7_75t_L g346 ( .A(n_226), .B(n_260), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_226), .B(n_259), .Y(n_374) );
OR2x2_ASAP7_75t_L g377 ( .A(n_226), .B(n_259), .Y(n_377) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_230), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_229), .A2(n_503), .B(n_504), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_229), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_234), .A2(n_265), .B(n_267), .Y(n_264) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g491 ( .A(n_239), .Y(n_491) );
INVx5_ASAP7_75t_SL g292 ( .A(n_240), .Y(n_292) );
OR2x2_ASAP7_75t_L g298 ( .A(n_240), .B(n_249), .Y(n_298) );
AND2x2_ASAP7_75t_L g314 ( .A(n_240), .B(n_315), .Y(n_314) );
AOI321xp33_ASAP7_75t_L g321 ( .A1(n_240), .A2(n_322), .A3(n_323), .B1(n_324), .B2(n_330), .C(n_332), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_240), .B(n_248), .Y(n_331) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_240), .Y(n_344) );
OR2x2_ASAP7_75t_L g391 ( .A(n_240), .B(n_289), .Y(n_391) );
AND2x2_ASAP7_75t_L g413 ( .A(n_240), .B(n_310), .Y(n_413) );
AND2x2_ASAP7_75t_L g432 ( .A(n_240), .B(n_250), .Y(n_432) );
OR2x6_ASAP7_75t_L g240 ( .A(n_241), .B(n_247), .Y(n_240) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_259), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_250), .B(n_259), .Y(n_273) );
AND2x2_ASAP7_75t_L g282 ( .A(n_250), .B(n_283), .Y(n_282) );
INVx3_ASAP7_75t_L g309 ( .A(n_250), .Y(n_309) );
AND2x2_ASAP7_75t_L g315 ( .A(n_250), .B(n_310), .Y(n_315) );
INVxp67_ASAP7_75t_L g345 ( .A(n_250), .Y(n_345) );
OR2x2_ASAP7_75t_L g387 ( .A(n_250), .B(n_292), .Y(n_387) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_258), .Y(n_250) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_251), .A2(n_478), .B(n_485), .Y(n_477) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_251), .A2(n_530), .B(n_537), .Y(n_529) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_251), .A2(n_539), .B(n_545), .Y(n_538) );
OR2x2_ASAP7_75t_L g269 ( .A(n_259), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_SL g283 ( .A(n_259), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_259), .B(n_272), .Y(n_316) );
AND2x2_ASAP7_75t_L g365 ( .A(n_259), .B(n_309), .Y(n_365) );
AND2x2_ASAP7_75t_L g403 ( .A(n_259), .B(n_292), .Y(n_403) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_260), .B(n_292), .Y(n_291) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_271), .B(n_274), .C(n_278), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_269), .A2(n_271), .B1(n_396), .B2(n_398), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_271), .A2(n_294), .B1(n_349), .B2(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_SL g423 ( .A(n_272), .Y(n_423) );
INVx1_ASAP7_75t_SL g323 ( .A(n_273), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_275), .B(n_295), .Y(n_325) );
AOI222xp33_ASAP7_75t_L g336 ( .A1(n_275), .A2(n_316), .B1(n_323), .B2(n_337), .C1(n_341), .C2(n_347), .Y(n_336) );
AND2x2_ASAP7_75t_L g426 ( .A(n_275), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx2_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_276), .B(n_296), .Y(n_371) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_276), .Y(n_408) );
AND2x2_ASAP7_75t_L g411 ( .A(n_276), .B(n_320), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_276), .B(n_427), .Y(n_437) );
INVx1_ASAP7_75t_L g328 ( .A(n_277), .Y(n_328) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_277), .Y(n_356) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_279), .A2(n_420), .B(n_421), .C(n_424), .Y(n_419) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_281), .B(n_343), .C(n_346), .Y(n_342) );
OR2x2_ASAP7_75t_L g370 ( .A(n_281), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_281), .B(n_297), .Y(n_398) );
OR2x2_ASAP7_75t_L g303 ( .A(n_283), .B(n_304), .Y(n_303) );
AOI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_287), .B(n_293), .C(n_305), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_286), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g392 ( .A(n_287), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_288), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g306 ( .A(n_291), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_292), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g360 ( .A(n_292), .B(n_310), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_292), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_292), .B(n_309), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_298), .B1(n_299), .B2(n_303), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_295), .B(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_297), .B(n_339), .Y(n_338) );
OAI221xp5_ASAP7_75t_SL g361 ( .A1(n_298), .A2(n_362), .B1(n_364), .B2(n_366), .C(n_368), .Y(n_361) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g416 ( .A(n_301), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g429 ( .A(n_301), .B(n_418), .Y(n_429) );
INVx1_ASAP7_75t_L g349 ( .A(n_302), .Y(n_349) );
INVx1_ASAP7_75t_L g420 ( .A(n_303), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_304), .A2(n_387), .B(n_410), .Y(n_409) );
AOI21xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_308), .B(n_311), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI21xp5_ASAP7_75t_SL g313 ( .A1(n_314), .A2(n_316), .B(n_317), .Y(n_313) );
INVx1_ASAP7_75t_L g353 ( .A(n_314), .Y(n_353) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_315), .A2(n_401), .B1(n_404), .B2(n_406), .C(n_409), .Y(n_400) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_323), .A2(n_413), .B1(n_414), .B2(n_416), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g389 ( .A(n_325), .Y(n_389) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NOR2xp67_ASAP7_75t_SL g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g393 ( .A(n_329), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g358 ( .A(n_334), .Y(n_358) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_339), .B(n_363), .Y(n_415) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_345), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g431 ( .A(n_346), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g438 ( .A(n_346), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI211xp5_ASAP7_75t_SL g350 ( .A1(n_351), .A2(n_353), .B(n_354), .C(n_388), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI211xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B(n_361), .C(n_380), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g441 ( .A(n_365), .Y(n_441) );
AND2x2_ASAP7_75t_L g378 ( .A(n_367), .B(n_379), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B1(n_376), .B2(n_378), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
OR2x2_ASAP7_75t_L g386 ( .A(n_374), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g439 ( .A(n_375), .Y(n_439) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI31xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .A3(n_383), .B(n_386), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI211xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B(n_392), .C(n_395), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g396 ( .A(n_397), .Y(n_396) );
NAND5xp2_ASAP7_75t_L g399 ( .A(n_400), .B(n_412), .C(n_419), .D(n_433), .E(n_436), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_411), .A2(n_437), .B1(n_438), .B2(n_440), .Y(n_436) );
INVx1_ASAP7_75t_SL g435 ( .A(n_413), .Y(n_435) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_428), .B(n_430), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g725 ( .A(n_449), .Y(n_725) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_457), .B1(n_460), .B2(n_723), .Y(n_455) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g727 ( .A(n_458), .Y(n_727) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR3x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_634), .C(n_681), .Y(n_461) );
NAND3xp33_ASAP7_75t_SL g462 ( .A(n_463), .B(n_580), .C(n_605), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_518), .B1(n_546), .B2(n_549), .C(n_557), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_486), .B(n_511), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_466), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_466), .B(n_562), .Y(n_678) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .Y(n_466) );
AND2x2_ASAP7_75t_L g548 ( .A(n_467), .B(n_517), .Y(n_548) );
AND2x2_ASAP7_75t_L g598 ( .A(n_467), .B(n_516), .Y(n_598) );
AND2x2_ASAP7_75t_L g619 ( .A(n_467), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g624 ( .A(n_467), .B(n_591), .Y(n_624) );
OR2x2_ASAP7_75t_L g632 ( .A(n_467), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g704 ( .A(n_467), .B(n_500), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_467), .B(n_653), .Y(n_718) );
INVx3_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g563 ( .A(n_468), .B(n_477), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_468), .B(n_500), .Y(n_564) );
AND2x4_ASAP7_75t_L g586 ( .A(n_468), .B(n_517), .Y(n_586) );
AND2x2_ASAP7_75t_L g616 ( .A(n_468), .B(n_488), .Y(n_616) );
AND2x2_ASAP7_75t_L g625 ( .A(n_468), .B(n_615), .Y(n_625) );
AND2x2_ASAP7_75t_L g641 ( .A(n_468), .B(n_501), .Y(n_641) );
OR2x2_ASAP7_75t_L g650 ( .A(n_468), .B(n_633), .Y(n_650) );
AND2x2_ASAP7_75t_L g656 ( .A(n_468), .B(n_591), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_468), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g670 ( .A(n_468), .B(n_513), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_468), .B(n_559), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_468), .B(n_620), .Y(n_709) );
OR2x6_ASAP7_75t_L g468 ( .A(n_469), .B(n_475), .Y(n_468) );
INVx2_ASAP7_75t_L g517 ( .A(n_477), .Y(n_517) );
AND2x2_ASAP7_75t_L g615 ( .A(n_477), .B(n_500), .Y(n_615) );
AND2x2_ASAP7_75t_L g620 ( .A(n_477), .B(n_501), .Y(n_620) );
INVx1_ASAP7_75t_L g676 ( .A(n_477), .Y(n_676) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g585 ( .A(n_487), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_500), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_488), .B(n_548), .Y(n_547) );
BUFx3_ASAP7_75t_L g562 ( .A(n_488), .Y(n_562) );
OR2x2_ASAP7_75t_L g633 ( .A(n_488), .B(n_500), .Y(n_633) );
OR2x2_ASAP7_75t_L g694 ( .A(n_488), .B(n_601), .Y(n_694) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_492), .B(n_499), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_490), .A2(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g514 ( .A(n_492), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_499), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_500), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g653 ( .A(n_500), .B(n_513), .Y(n_653) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g592 ( .A(n_501), .Y(n_592) );
INVx1_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_512), .A2(n_698), .B1(n_702), .B2(n_705), .C(n_706), .Y(n_697) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
INVx1_ASAP7_75t_SL g560 ( .A(n_513), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_513), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g692 ( .A(n_513), .B(n_548), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_516), .B(n_562), .Y(n_684) );
AND2x2_ASAP7_75t_L g591 ( .A(n_517), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g595 ( .A(n_518), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_518), .B(n_601), .Y(n_631) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
AND2x2_ASAP7_75t_L g556 ( .A(n_519), .B(n_529), .Y(n_556) );
INVx4_ASAP7_75t_L g568 ( .A(n_519), .Y(n_568) );
BUFx3_ASAP7_75t_L g611 ( .A(n_519), .Y(n_611) );
AND3x2_ASAP7_75t_L g626 ( .A(n_519), .B(n_627), .C(n_628), .Y(n_626) );
AND2x2_ASAP7_75t_L g708 ( .A(n_528), .B(n_622), .Y(n_708) );
AND2x2_ASAP7_75t_L g716 ( .A(n_528), .B(n_601), .Y(n_716) );
INVx1_ASAP7_75t_SL g721 ( .A(n_528), .Y(n_721) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
INVx1_ASAP7_75t_SL g579 ( .A(n_529), .Y(n_579) );
AND2x2_ASAP7_75t_L g602 ( .A(n_529), .B(n_568), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_529), .B(n_552), .Y(n_604) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_529), .Y(n_644) );
OR2x2_ASAP7_75t_L g649 ( .A(n_529), .B(n_568), .Y(n_649) );
INVx2_ASAP7_75t_L g554 ( .A(n_538), .Y(n_554) );
AND2x2_ASAP7_75t_L g589 ( .A(n_538), .B(n_569), .Y(n_589) );
OR2x2_ASAP7_75t_L g609 ( .A(n_538), .B(n_569), .Y(n_609) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_538), .Y(n_629) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AOI21xp33_ASAP7_75t_L g679 ( .A1(n_547), .A2(n_588), .B(n_680), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g715 ( .A1(n_549), .A2(n_559), .A3(n_586), .B1(n_716), .B2(n_717), .C1(n_719), .C2(n_722), .Y(n_715) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_555), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_551), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_552), .B(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g578 ( .A(n_553), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g646 ( .A(n_554), .B(n_568), .Y(n_646) );
AND2x2_ASAP7_75t_L g713 ( .A(n_554), .B(n_569), .Y(n_713) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g654 ( .A(n_556), .B(n_608), .Y(n_654) );
AOI31xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .A3(n_564), .B(n_565), .Y(n_557) );
AND2x2_ASAP7_75t_L g613 ( .A(n_559), .B(n_591), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_559), .B(n_583), .Y(n_695) );
AND2x2_ASAP7_75t_L g714 ( .A(n_559), .B(n_619), .Y(n_714) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_562), .B(n_591), .Y(n_603) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_562), .B(n_620), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_562), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_562), .B(n_704), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_563), .B(n_620), .Y(n_652) );
INVx1_ASAP7_75t_L g696 ( .A(n_563), .Y(n_696) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_578), .Y(n_566) );
INVxp67_ASAP7_75t_L g648 ( .A(n_567), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_568), .B(n_579), .Y(n_584) );
INVx1_ASAP7_75t_L g690 ( .A(n_568), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_568), .B(n_667), .Y(n_701) );
BUFx3_ASAP7_75t_L g601 ( .A(n_569), .Y(n_601) );
AND2x2_ASAP7_75t_L g627 ( .A(n_569), .B(n_579), .Y(n_627) );
INVx2_ASAP7_75t_L g667 ( .A(n_569), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_578), .B(n_700), .Y(n_699) );
AOI211xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_585), .B(n_587), .C(n_596), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI21xp33_ASAP7_75t_L g630 ( .A1(n_582), .A2(n_631), .B(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_583), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_583), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g663 ( .A(n_584), .B(n_609), .Y(n_663) );
INVx3_ASAP7_75t_L g594 ( .A(n_586), .Y(n_594) );
OAI22xp5_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_590), .B1(n_593), .B2(n_595), .Y(n_587) );
OAI21xp5_ASAP7_75t_SL g612 ( .A1(n_589), .A2(n_613), .B(n_614), .Y(n_612) );
AND2x2_ASAP7_75t_L g638 ( .A(n_589), .B(n_602), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_589), .B(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g593 ( .A(n_592), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g662 ( .A(n_592), .Y(n_662) );
OAI21xp5_ASAP7_75t_SL g606 ( .A1(n_593), .A2(n_607), .B(n_612), .Y(n_606) );
OAI22xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_599), .B1(n_603), .B2(n_604), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_598), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g622 ( .A(n_601), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_601), .B(n_644), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_617), .C(n_630), .Y(n_605) );
OAI22xp5_ASAP7_75t_SL g672 ( .A1(n_607), .A2(n_673), .B1(n_677), .B2(n_678), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g677 ( .A(n_609), .B(n_610), .Y(n_677) );
AND2x2_ASAP7_75t_L g685 ( .A(n_610), .B(n_666), .Y(n_685) );
CKINVDCx16_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_SL g693 ( .A1(n_611), .A2(n_694), .B(n_695), .C(n_696), .Y(n_693) );
OR2x2_ASAP7_75t_L g720 ( .A(n_611), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B(n_623), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_619), .A2(n_656), .B(n_657), .C(n_660), .Y(n_655) );
OAI21xp33_ASAP7_75t_SL g623 ( .A1(n_624), .A2(n_625), .B(n_626), .Y(n_623) );
AND2x2_ASAP7_75t_L g688 ( .A(n_627), .B(n_646), .Y(n_688) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g666 ( .A(n_629), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g671 ( .A(n_631), .Y(n_671) );
NAND3xp33_ASAP7_75t_SL g634 ( .A(n_635), .B(n_655), .C(n_668), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B(n_639), .C(n_647), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g705 ( .A(n_642), .Y(n_705) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g665 ( .A(n_644), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_644), .B(n_713), .Y(n_712) );
INVxp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B(n_650), .C(n_651), .Y(n_647) );
INVx2_ASAP7_75t_SL g659 ( .A(n_649), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_650), .A2(n_661), .B1(n_663), .B2(n_664), .Y(n_660) );
OAI21xp33_ASAP7_75t_SL g651 ( .A1(n_652), .A2(n_653), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B(n_672), .C(n_679), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
INVxp33_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g722 ( .A(n_676), .Y(n_722) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_682), .B(n_697), .C(n_710), .D(n_715), .Y(n_681) );
AOI211xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_685), .B(n_686), .C(n_693), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_691), .Y(n_686) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_687), .A2(n_707), .B(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_694), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_714), .Y(n_710) );
INVxp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g729 ( .A(n_723), .Y(n_729) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
endmodule