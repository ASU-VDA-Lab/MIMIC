module fake_ariane_43_n_186 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_186);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;

output n_186;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_178;
wire n_42;
wire n_31;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_144;
wire n_130;
wire n_85;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_28;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVxp33_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_7),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_43),
.B(n_0),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_4),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_6),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_8),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

AO22x2_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_42),
.B1(n_35),
.B2(n_38),
.Y(n_67)
);

AO22x2_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_38),
.B1(n_28),
.B2(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2x1p5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_27),
.Y(n_74)
);

NAND2x1p5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_45),
.Y(n_75)
);

AO22x2_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_10),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_21),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

AND3x1_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_66),
.C(n_63),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_54),
.B1(n_56),
.B2(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_59),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_81),
.B(n_56),
.C(n_77),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_67),
.B1(n_54),
.B2(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_68),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AND2x4_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_63),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_67),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_93),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_95),
.B(n_89),
.C(n_60),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_53),
.B(n_93),
.C(n_90),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_88),
.Y(n_108)
);

NOR2x1_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_91),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

OR2x6_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_91),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_103),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_98),
.B1(n_74),
.B2(n_68),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_106),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_112),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_112),
.A2(n_104),
.B(n_105),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_103),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_108),
.B1(n_76),
.B2(n_102),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_108),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_74),
.B1(n_80),
.B2(n_76),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_108),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_121),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_116),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_120),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_119),
.C(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_118),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_132),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_80),
.B(n_52),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_140),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_65),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_132),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_10),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_118),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_120),
.Y(n_152)
);

NOR2x1p5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_139),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_151),
.B(n_124),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_51),
.C(n_62),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_69),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_80),
.B1(n_117),
.B2(n_108),
.Y(n_158)
);

NAND2x1p5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_125),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_65),
.Y(n_161)
);

NOR2x1p5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_59),
.Y(n_162)
);

AOI221x1_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_151),
.B1(n_51),
.B2(n_62),
.C(n_65),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_62),
.Y(n_165)
);

NOR3x1_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_52),
.C(n_66),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_158),
.A2(n_49),
.B(n_102),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_49),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_155),
.B1(n_157),
.B2(n_125),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_49),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_109),
.Y(n_173)
);

AOI211xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_49),
.B(n_13),
.C(n_14),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_11),
.Y(n_175)
);

OAI211xp5_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_11),
.B(n_14),
.C(n_15),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_167),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_162),
.B1(n_169),
.B2(n_167),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_177),
.A3(n_176),
.B1(n_174),
.B2(n_166),
.C1(n_175),
.C2(n_85),
.Y(n_179)
);

AOI221xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_61),
.B1(n_108),
.B2(n_163),
.C(n_94),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_107),
.B1(n_100),
.B2(n_61),
.Y(n_181)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_90),
.C(n_87),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_109),
.B(n_92),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_61),
.B1(n_17),
.B2(n_16),
.Y(n_184)
);

OR2x6_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_179),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_183),
.B1(n_182),
.B2(n_24),
.Y(n_186)
);


endmodule