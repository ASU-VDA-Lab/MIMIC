module real_jpeg_26186_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx6_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_0),
.Y(n_158)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_0),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_4),
.A2(n_113),
.B(n_115),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_77),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_53),
.C(n_63),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_31),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_4),
.A2(n_80),
.B1(n_172),
.B2(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_68),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_68),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_7),
.A2(n_36),
.B1(n_109),
.B2(n_110),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_7),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_8),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_57),
.Y(n_122)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_14),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_72),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_15),
.A2(n_28),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_15),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_128),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_19),
.B(n_88),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_59),
.C(n_73),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_20),
.A2(n_21),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_22),
.B(n_41),
.C(n_47),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_23),
.A2(n_37),
.B1(n_39),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_24),
.A2(n_31),
.B1(n_35),
.B2(n_76),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_26),
.B(n_32),
.Y(n_78)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI32xp33_ASAP7_75t_L g75 ( 
.A1(n_27),
.A2(n_30),
.A3(n_33),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g76 ( 
.A(n_28),
.B(n_77),
.CON(n_76),
.SN(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_28),
.A2(n_45),
.B(n_92),
.C(n_95),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_30),
.B(n_44),
.C(n_93),
.Y(n_95)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_32),
.A2(n_33),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_33),
.B(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_44),
.A2(n_45),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_55),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_52),
.Y(n_58)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_50),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_53),
.B1(n_63),
.B2(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_52),
.B(n_179),
.Y(n_178)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_86),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_58),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_59),
.A2(n_60),
.B1(n_73),
.B2(n_74),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_67),
.B(n_69),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_61),
.A2(n_71),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_61),
.A2(n_67),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_61),
.A2(n_135),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_61),
.A2(n_134),
.B1(n_135),
.B2(n_145),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_66),
.B(n_77),
.Y(n_170)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_75),
.B(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_77),
.B(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_83),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_80),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_80),
.A2(n_163),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_82),
.B(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_87),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_103),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_102),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_96),
.B1(n_100),
.B2(n_101),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_118),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_107),
.B1(n_112),
.B2(n_116),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_139),
.B(n_190),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_130),
.B(n_136),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.C(n_133),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_132),
.B(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_185),
.B(n_189),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_159),
.B(n_184),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_142),
.B(n_148),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_146),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_153),
.C(n_154),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_168),
.B(n_183),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_167),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_175),
.B(n_182),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_170),
.B(n_171),
.Y(n_182)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_178),
.Y(n_175)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_187),
.Y(n_189)
);


endmodule