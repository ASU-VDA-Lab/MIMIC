module fake_aes_3878_n_26 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_26);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
AOI22x1_ASAP7_75t_SL g10 ( .A1(n_8), .A2(n_6), .B1(n_3), .B2(n_7), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
HB1xp67_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
INVx5_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
OR2x6_ASAP7_75t_L g17 ( .A(n_14), .B(n_11), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_17), .B(n_15), .Y(n_18) );
OR2x2_ASAP7_75t_L g19 ( .A(n_18), .B(n_17), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_17), .B1(n_16), .B2(n_10), .Y(n_21) );
OAI211xp5_ASAP7_75t_SL g22 ( .A1(n_21), .A2(n_16), .B(n_1), .C(n_2), .Y(n_22) );
OR5x1_ASAP7_75t_L g23 ( .A(n_21), .B(n_0), .C(n_3), .D(n_4), .E(n_5), .Y(n_23) );
OAI22xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_22), .B1(n_16), .B2(n_6), .Y(n_24) );
AOI22xp5_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_16), .B1(n_5), .B2(n_9), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
endmodule