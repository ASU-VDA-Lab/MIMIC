module fake_jpeg_19220_n_201 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_201);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_39),
.Y(n_51)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_14),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_45),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_3),
.C(n_4),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_40),
.B1(n_39),
.B2(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_25),
.B1(n_15),
.B2(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_60),
.B1(n_57),
.B2(n_53),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_54),
.B1(n_40),
.B2(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_25),
.B1(n_26),
.B2(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_18),
.B1(n_15),
.B2(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_76),
.B1(n_80),
.B2(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_72),
.Y(n_105)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_33),
.B1(n_45),
.B2(n_35),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_64),
.B1(n_43),
.B2(n_58),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_38),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_38),
.Y(n_76)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_37),
.B(n_42),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_81),
.C(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_44),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_42),
.B1(n_37),
.B2(n_33),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_43),
.B(n_24),
.C(n_28),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_49),
.A2(n_31),
.B1(n_30),
.B2(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_90),
.Y(n_97)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_24),
.CI(n_31),
.CON(n_87),
.SN(n_87)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_81),
.B1(n_77),
.B2(n_87),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_43),
.B1(n_30),
.B2(n_29),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_94),
.B1(n_29),
.B2(n_19),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_27),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_52),
.B(n_3),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_79),
.C(n_66),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_106),
.C(n_104),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_73),
.A2(n_29),
.B1(n_19),
.B2(n_16),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_19),
.C(n_16),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_27),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_86),
.A2(n_17),
.B1(n_21),
.B2(n_6),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_113),
.B1(n_82),
.B2(n_5),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_113)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_120),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_106),
.Y(n_137)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_123),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_85),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_88),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_111),
.B1(n_109),
.B2(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_65),
.B(n_85),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_100),
.B(n_70),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_132),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_78),
.B1(n_84),
.B2(n_7),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_131),
.B1(n_112),
.B2(n_97),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_78),
.B1(n_84),
.B2(n_7),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_117),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_116),
.C(n_133),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_114),
.B(n_110),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_149),
.B(n_4),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_140),
.B(n_135),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_141),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_121),
.B(n_125),
.C(n_119),
.D(n_123),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_17),
.B(n_21),
.C(n_8),
.D(n_10),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_147),
.A2(n_117),
.B1(n_129),
.B2(n_118),
.Y(n_156)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_154),
.C(n_136),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_130),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_156),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_150),
.B1(n_141),
.B2(n_149),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_120),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_159),
.B(n_162),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_115),
.Y(n_160)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_168),
.C(n_171),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_136),
.C(n_145),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_148),
.C(n_146),
.Y(n_182)
);

OAI321xp33_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_142),
.A3(n_138),
.B1(n_139),
.B2(n_141),
.C(n_147),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_153),
.B(n_160),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_171),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_153),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_174),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_167),
.A2(n_158),
.B(n_162),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_175),
.B(n_176),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_151),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_178),
.C(n_179),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_161),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_182),
.C(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_187),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_172),
.C(n_159),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_169),
.C(n_146),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_152),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_190),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_180),
.B1(n_179),
.B2(n_152),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_183),
.B(n_115),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_6),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_191),
.A2(n_70),
.B(n_8),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_190),
.B(n_8),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_193),
.B(n_11),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_11),
.B(n_12),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_12),
.Y(n_201)
);


endmodule