module real_jpeg_1626_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_0),
.A2(n_42),
.B1(n_60),
.B2(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_0),
.A2(n_42),
.B1(n_71),
.B2(n_73),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_0),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_2),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_37),
.B1(n_39),
.B2(n_143),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_2),
.A2(n_71),
.B1(n_73),
.B2(n_143),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_2),
.A2(n_60),
.B1(n_66),
.B2(n_143),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_4),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_4),
.A2(n_37),
.B1(n_39),
.B2(n_87),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_71),
.B1(n_73),
.B2(n_87),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g213 ( 
.A1(n_4),
.A2(n_60),
.B1(n_66),
.B2(n_87),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_6),
.A2(n_45),
.B1(n_71),
.B2(n_73),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_6),
.A2(n_37),
.B1(n_39),
.B2(n_45),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_45),
.B1(n_60),
.B2(n_66),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_7),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_7),
.A2(n_37),
.B1(n_39),
.B2(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_70),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_7),
.A2(n_60),
.B1(n_66),
.B2(n_70),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_8),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_8),
.A2(n_37),
.B1(n_39),
.B2(n_85),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_8),
.A2(n_71),
.B1(n_73),
.B2(n_85),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_8),
.A2(n_60),
.B1(n_66),
.B2(n_85),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_9),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_9),
.A2(n_37),
.B1(n_39),
.B2(n_177),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_9),
.A2(n_71),
.B1(n_73),
.B2(n_177),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_9),
.A2(n_60),
.B1(n_66),
.B2(n_177),
.Y(n_279)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_14),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_14),
.A2(n_37),
.B1(n_39),
.B2(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_14),
.A2(n_71),
.B1(n_73),
.B2(n_196),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_14),
.A2(n_60),
.B1(n_66),
.B2(n_196),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_15),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_16),
.A2(n_37),
.B1(n_39),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_16),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_93),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_16),
.A2(n_71),
.B1(n_73),
.B2(n_93),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_16),
.A2(n_60),
.B1(n_66),
.B2(n_93),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_17),
.B(n_30),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_17),
.B(n_40),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_17),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_17),
.A2(n_30),
.B(n_186),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_17),
.B(n_96),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g254 ( 
.A1(n_17),
.A2(n_39),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_17),
.B(n_60),
.C(n_76),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_17),
.A2(n_71),
.B1(n_73),
.B2(n_222),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_17),
.B(n_63),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_17),
.B(n_80),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_46),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_47),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_40),
.B(n_41),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_28),
.A2(n_40),
.B1(n_142),
.B2(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_28),
.A2(n_40),
.B1(n_44),
.B2(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI32xp33_ASAP7_75t_L g185 ( 
.A1(n_31),
.A2(n_35),
.A3(n_39),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_33),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_33),
.B(n_37),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_36),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_36),
.A2(n_83),
.B1(n_86),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_36),
.A2(n_83),
.B1(n_84),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_36),
.A2(n_83),
.B1(n_106),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_36),
.A2(n_83),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_36),
.A2(n_83),
.B1(n_195),
.B2(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_37),
.A2(n_39),
.B1(n_97),
.B2(n_98),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_37),
.B(n_222),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g220 ( 
.A1(n_39),
.A2(n_71),
.A3(n_97),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_43),
.B(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_47),
.B(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_327),
.B(n_329),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_315),
.B(n_326),
.Y(n_49)
);

AO21x1_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_157),
.B(n_312),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_144),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_117),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_53),
.B(n_117),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_88),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_54),
.B(n_103),
.C(n_115),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_81),
.B(n_82),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_55),
.A2(n_56),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_67),
.Y(n_56)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_57),
.A2(n_81),
.B1(n_82),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_57),
.A2(n_67),
.B1(n_68),
.B2(n_81),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_64),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_58),
.A2(n_62),
.B1(n_131),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_58),
.A2(n_62),
.B1(n_225),
.B2(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_58),
.A2(n_62),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_59),
.A2(n_63),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_59),
.A2(n_63),
.B1(n_189),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_59),
.A2(n_63),
.B1(n_226),
.B2(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_59),
.A2(n_63),
.B1(n_222),
.B2(n_275),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_59),
.A2(n_63),
.B1(n_275),
.B2(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_66),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_60),
.B(n_273),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_69),
.A2(n_74),
.B1(n_80),
.B2(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_71),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

AO22x2_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_73),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_71),
.B(n_263),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_73),
.B(n_98),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_80),
.B(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_74),
.A2(n_80),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_74),
.A2(n_80),
.B1(n_218),
.B2(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_74),
.A2(n_80),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_74),
.A2(n_80),
.B1(n_245),
.B2(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_78),
.A2(n_135),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_78),
.A2(n_170),
.B1(n_217),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_103),
.B1(n_115),
.B2(n_116),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_90),
.B(n_101),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_101),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_94),
.B1(n_96),
.B2(n_100),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_92),
.A2(n_95),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_96),
.B1(n_100),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_94),
.A2(n_96),
.B1(n_138),
.B2(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_94),
.A2(n_96),
.B(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_95),
.A2(n_113),
.B1(n_139),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_95),
.A2(n_139),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_95),
.A2(n_139),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_95),
.A2(n_139),
.B1(n_192),
.B2(n_208),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_95),
.A2(n_139),
.B1(n_207),
.B2(n_254),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_107),
.B2(n_108),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_104),
.A2(n_105),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_109),
.C(n_111),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_105),
.B(n_148),
.C(n_155),
.Y(n_316)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_114),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_109),
.B(n_151),
.C(n_153),
.Y(n_325)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.C(n_125),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_118),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_136),
.C(n_140),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_127),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_198)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_140),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_144),
.A2(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_156),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_145),
.B(n_156),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_152),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_154),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_178),
.B(n_311),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_159),
.B(n_161),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_166),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_173),
.C(n_175),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_168),
.B(n_171),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_175),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_174),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_201),
.B(n_310),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_199),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_180),
.B(n_199),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_198),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_181),
.B(n_198),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_183),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_191),
.C(n_194),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_184),
.B(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_188),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_191),
.B(n_194),
.Y(n_301)
);

AOI31xp33_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_295),
.A3(n_304),
.B(n_307),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_240),
.B(n_294),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_228),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_204),
.B(n_228),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_215),
.C(n_219),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_205),
.B(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_210),
.C(n_214),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_215),
.B(n_219),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_228),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_228),
.B(n_305),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_230),
.CI(n_231),
.CON(n_228),
.SN(n_228)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_232),
.B(n_235),
.C(n_239),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_289),
.B(n_293),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_258),
.B(n_288),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_250),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.C(n_248),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_247),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_253),
.C(n_256),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_269),
.B(n_287),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_267),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_281),
.B(n_286),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_276),
.B(n_280),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_278),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_279),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_285),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_285),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_292),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_299),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_303),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_317),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_321),
.B1(n_323),
.B2(n_324),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_321),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_323),
.C(n_325),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_328),
.Y(n_331)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule