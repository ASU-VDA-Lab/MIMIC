module fake_jpeg_27775_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_11),
.B1(n_13),
.B2(n_7),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_17),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_1),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_19),
.Y(n_23)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_20),
.B(n_10),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_20),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_14),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_16),
.B1(n_19),
.B2(n_11),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_31),
.Y(n_33)
);

NOR4xp25_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_17),
.C(n_16),
.D(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_15),
.B1(n_19),
.B2(n_13),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_22),
.C(n_23),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_21),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_16),
.B(n_2),
.Y(n_37)
);

OAI211xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_39),
.B(n_12),
.C(n_8),
.Y(n_41)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_41),
.C2(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_42),
.Y(n_43)
);


endmodule