module fake_jpeg_27_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_55),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g59 ( 
.A(n_56),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_64),
.A2(n_49),
.B1(n_54),
.B2(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_93),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_51),
.C(n_48),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_41),
.Y(n_85)
);

OR2x2_ASAP7_75t_SL g87 ( 
.A(n_69),
.B(n_49),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_89),
.B(n_92),
.Y(n_96)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_72),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

OR2x6_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_73),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_18),
.C(n_38),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_42),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_42),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_61),
.B1(n_54),
.B2(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_70),
.B1(n_57),
.B2(n_2),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_92),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_4),
.Y(n_129)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_121),
.B(n_20),
.Y(n_135)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_119),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_17),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_13),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_125),
.C(n_27),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_1),
.B(n_3),
.Y(n_121)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_123),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_19),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_102),
.C(n_109),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_4),
.CI(n_5),
.CON(n_127),
.SN(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_128),
.B(n_8),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_25),
.B1(n_37),
.B2(n_36),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_133),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_5),
.B(n_7),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_136),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_SL g142 ( 
.A(n_137),
.B(n_138),
.C(n_112),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_144),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_117),
.B1(n_113),
.B2(n_127),
.Y(n_144)
);

OAI321xp33_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_123),
.A3(n_119),
.B1(n_120),
.B2(n_111),
.C(n_29),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_145),
.B(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_141),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_137),
.C(n_132),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_146),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_151),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_147),
.B(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_131),
.A3(n_134),
.B1(n_11),
.B2(n_12),
.C1(n_31),
.C2(n_34),
.Y(n_156)
);

NAND2x1_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_40),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_10),
.Y(n_158)
);


endmodule