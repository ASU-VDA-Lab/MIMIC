module fake_ariane_205_n_1546 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_424, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_350, n_291, n_344, n_381, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_420, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_417, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_418, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_1546);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_424;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_420;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_417;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_418;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_1546;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_1495;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_512;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_436;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_1521;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_519;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_917;
wire n_1271;
wire n_1530;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_946;
wire n_757;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_849;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_392),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_122),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_274),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_391),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_48),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_68),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_199),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_111),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_163),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_414),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_231),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_417),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_343),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_270),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_240),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_222),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_410),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_25),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_309),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_339),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_359),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_116),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_64),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_156),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_157),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_331),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_201),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_88),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_114),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_219),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_4),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_29),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_64),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_397),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_246),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_404),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_265),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_119),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_155),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_177),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_356),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_161),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_205),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_140),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_269),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_194),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_136),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_217),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_372),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_225),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_382),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_182),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_210),
.Y(n_478)
);

BUFx5_ASAP7_75t_L g479 ( 
.A(n_1),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_191),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_393),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_267),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_345),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_268),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_17),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_32),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_310),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_102),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_236),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_136),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_282),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_164),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_376),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_127),
.Y(n_494)
);

INVxp33_ASAP7_75t_L g495 ( 
.A(n_48),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_70),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_26),
.B(n_56),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_31),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_232),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_144),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_299),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_132),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_321),
.Y(n_503)
);

CKINVDCx14_ASAP7_75t_R g504 ( 
.A(n_167),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_327),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_348),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_314),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_301),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_78),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_63),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_370),
.Y(n_511)
);

CKINVDCx14_ASAP7_75t_R g512 ( 
.A(n_303),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_195),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_354),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_351),
.B(n_334),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_227),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_237),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_371),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_365),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_87),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_317),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_377),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_316),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_27),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_400),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_95),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_9),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_69),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_6),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_36),
.Y(n_530)
);

BUFx2_ASAP7_75t_SL g531 ( 
.A(n_329),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_151),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_171),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_37),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_8),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_289),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_120),
.B(n_313),
.Y(n_537)
);

BUFx5_ASAP7_75t_L g538 ( 
.A(n_203),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_364),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_10),
.Y(n_540)
);

CKINVDCx14_ASAP7_75t_R g541 ( 
.A(n_78),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_273),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_153),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_190),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_87),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_322),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_390),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_180),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_165),
.B(n_352),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_271),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_242),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_253),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_202),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_162),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_101),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_415),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_91),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_52),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_173),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_277),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_0),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_149),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_9),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_234),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_295),
.Y(n_565)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_315),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_319),
.B(n_196),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_412),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_204),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_130),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_389),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_394),
.Y(n_572)
);

NOR2xp67_ASAP7_75t_L g573 ( 
.A(n_402),
.B(n_85),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_398),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_257),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_85),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_375),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_251),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_342),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_387),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_58),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_27),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_41),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_422),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_129),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_381),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_388),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_367),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_170),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_386),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_383),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_198),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_408),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_26),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_57),
.Y(n_595)
);

CKINVDCx16_ASAP7_75t_R g596 ( 
.A(n_275),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_6),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_291),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_223),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_211),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_332),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_235),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_403),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_46),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_226),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_52),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_272),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_298),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_147),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_337),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_456),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_479),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_496),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_479),
.Y(n_614)
);

OAI22x1_ASAP7_75t_SL g615 ( 
.A1(n_430),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_541),
.B(n_2),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_482),
.B(n_3),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_479),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_479),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_479),
.B(n_3),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_464),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_479),
.B(n_5),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_440),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_464),
.Y(n_624)
);

NOR2x1_ASAP7_75t_L g625 ( 
.A(n_536),
.B(n_137),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_464),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_546),
.B(n_5),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_486),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_529),
.A2(n_495),
.B1(n_528),
.B2(n_602),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_442),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_525),
.Y(n_631)
);

OA21x2_ASAP7_75t_L g632 ( 
.A1(n_431),
.A2(n_7),
.B(n_8),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_606),
.A2(n_12),
.B1(n_7),
.B2(n_11),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_446),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_545),
.B(n_11),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_454),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_559),
.B(n_12),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_494),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_453),
.Y(n_640)
);

OA21x2_ASAP7_75t_L g641 ( 
.A1(n_433),
.A2(n_13),
.B(n_14),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_462),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_485),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_563),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_488),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_490),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_498),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_509),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_510),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_520),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_526),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_530),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_534),
.Y(n_653)
);

OA21x2_ASAP7_75t_L g654 ( 
.A1(n_434),
.A2(n_13),
.B(n_14),
.Y(n_654)
);

BUFx8_ASAP7_75t_L g655 ( 
.A(n_507),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_528),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_656)
);

OAI21x1_ASAP7_75t_L g657 ( 
.A1(n_428),
.A2(n_139),
.B(n_138),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_535),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_592),
.B(n_16),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_525),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_438),
.B(n_18),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_540),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_525),
.Y(n_663)
);

AND2x2_ASAP7_75t_SL g664 ( 
.A(n_596),
.B(n_18),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_548),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_555),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_551),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_558),
.B(n_19),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_561),
.B(n_581),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_576),
.Y(n_670)
);

OA21x2_ASAP7_75t_L g671 ( 
.A1(n_445),
.A2(n_19),
.B(n_20),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_448),
.B(n_20),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_449),
.B(n_458),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_551),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_460),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_551),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_583),
.B(n_21),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_585),
.Y(n_678)
);

AOI22x1_ASAP7_75t_SL g679 ( 
.A1(n_475),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_553),
.B(n_141),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_463),
.B(n_22),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_594),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_595),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_597),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_468),
.B(n_23),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_469),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_604),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_471),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_467),
.Y(n_689)
);

CKINVDCx8_ASAP7_75t_R g690 ( 
.A(n_531),
.Y(n_690)
);

CKINVDCx16_ASAP7_75t_R g691 ( 
.A(n_467),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_554),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_553),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_474),
.B(n_24),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_553),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_476),
.B(n_25),
.Y(n_696)
);

CKINVDCx11_ASAP7_75t_R g697 ( 
.A(n_554),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_580),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_617),
.B(n_537),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_629),
.A2(n_502),
.B1(n_527),
.B2(n_576),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_616),
.B(n_538),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_665),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_623),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_614),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_617),
.B(n_537),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_668),
.A2(n_497),
.B1(n_512),
.B2(n_504),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_619),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_612),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_621),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_665),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_621),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_627),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_691),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_655),
.B(n_483),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_690),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_668),
.A2(n_497),
.B1(n_505),
.B2(n_425),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_689),
.B(n_427),
.Y(n_717)
);

BUFx10_ASAP7_75t_L g718 ( 
.A(n_627),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_629),
.A2(n_600),
.B1(n_603),
.B2(n_539),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_636),
.B(n_427),
.Y(n_720)
);

INVx5_ASAP7_75t_L g721 ( 
.A(n_680),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_656),
.B(n_573),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_618),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_693),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_656),
.B(n_439),
.Y(n_725)
);

AND2x2_ASAP7_75t_SL g726 ( 
.A(n_664),
.B(n_549),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_680),
.Y(n_727)
);

OAI22x1_ASAP7_75t_L g728 ( 
.A1(n_628),
.A2(n_426),
.B1(n_432),
.B2(n_429),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_675),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_636),
.B(n_439),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_677),
.A2(n_505),
.B1(n_566),
.B2(n_425),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_664),
.B(n_470),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_621),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_638),
.B(n_452),
.C(n_447),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_634),
.A2(n_670),
.B1(n_633),
.B2(n_659),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_633),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_697),
.Y(n_737)
);

INVx6_ASAP7_75t_L g738 ( 
.A(n_693),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_670),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_621),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_624),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_640),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_680),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_611),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_643),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_624),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_677),
.B(n_470),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_692),
.B(n_489),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_624),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_624),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_611),
.B(n_499),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_697),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_630),
.B(n_491),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_626),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_724),
.B(n_744),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_SL g756 ( 
.A1(n_719),
.A2(n_726),
.B1(n_637),
.B2(n_725),
.Y(n_756)
);

OAI21xp5_ASAP7_75t_L g757 ( 
.A1(n_708),
.A2(n_723),
.B(n_701),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_720),
.B(n_686),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_702),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_742),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_720),
.B(n_688),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_730),
.B(n_673),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_731),
.B(n_716),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_702),
.B(n_669),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_715),
.B(n_613),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_730),
.B(n_673),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_739),
.B(n_613),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_699),
.B(n_681),
.Y(n_768)
);

O2A1O1Ixp5_ASAP7_75t_L g769 ( 
.A1(n_699),
.A2(n_620),
.B(n_622),
.C(n_661),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_705),
.B(n_681),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_704),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_738),
.B(n_638),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_731),
.B(n_500),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_716),
.B(n_513),
.Y(n_774)
);

AND2x6_ASAP7_75t_L g775 ( 
.A(n_715),
.B(n_625),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_710),
.B(n_669),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_704),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_705),
.B(n_661),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_706),
.B(n_514),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_703),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_747),
.B(n_672),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_701),
.A2(n_622),
.B(n_620),
.Y(n_782)
);

BUFx12f_ASAP7_75t_L g783 ( 
.A(n_713),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_738),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_710),
.Y(n_785)
);

OAI221xp5_ASAP7_75t_L g786 ( 
.A1(n_706),
.A2(n_634),
.B1(n_735),
.B2(n_732),
.C(n_659),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_751),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_725),
.B(n_722),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_738),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_717),
.B(n_685),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_712),
.B(n_517),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_717),
.B(n_685),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_736),
.B(n_639),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_707),
.B(n_694),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_712),
.B(n_694),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_732),
.A2(n_726),
.B1(n_725),
.B2(n_753),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_718),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_718),
.B(n_696),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_750),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_753),
.B(n_645),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_745),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_714),
.B(n_696),
.Y(n_802)
);

AND2x2_ASAP7_75t_SL g803 ( 
.A(n_734),
.B(n_632),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_750),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_729),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_709),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_748),
.B(n_648),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_727),
.B(n_518),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_753),
.B(n_639),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_727),
.B(n_521),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_709),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_743),
.B(n_523),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_743),
.B(n_721),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_711),
.B(n_649),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_SL g815 ( 
.A1(n_722),
.A2(n_637),
.B1(n_615),
.B2(n_567),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_737),
.B(n_644),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_733),
.B(n_652),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_733),
.B(n_658),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_740),
.B(n_662),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_741),
.B(n_682),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_746),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_752),
.B(n_644),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_728),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_722),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_746),
.B(n_683),
.Y(n_825)
);

OAI21x1_ASAP7_75t_L g826 ( 
.A1(n_782),
.A2(n_657),
.B(n_515),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_804),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_795),
.B(n_798),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_755),
.A2(n_566),
.B(n_721),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_786),
.A2(n_700),
.B1(n_568),
.B2(n_588),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_790),
.A2(n_568),
.B1(n_588),
.B2(n_491),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_792),
.A2(n_684),
.B(n_607),
.C(n_642),
.Y(n_832)
);

BUFx4f_ASAP7_75t_L g833 ( 
.A(n_783),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_SL g834 ( 
.A1(n_778),
.A2(n_607),
.B(n_515),
.C(n_532),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_789),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_771),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_794),
.A2(n_721),
.B(n_641),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_796),
.A2(n_763),
.B1(n_798),
.B2(n_795),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_807),
.B(n_578),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_802),
.A2(n_721),
.B(n_641),
.Y(n_840)
);

OAI21xp33_ASAP7_75t_L g841 ( 
.A1(n_768),
.A2(n_770),
.B(n_781),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_769),
.A2(n_654),
.B(n_632),
.Y(n_842)
);

BUFx12f_ASAP7_75t_L g843 ( 
.A(n_797),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_816),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_777),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_759),
.B(n_635),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_780),
.B(n_800),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_757),
.A2(n_671),
.B(n_654),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_814),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_785),
.B(n_646),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_789),
.Y(n_851)
);

AOI22x1_ASAP7_75t_L g852 ( 
.A1(n_801),
.A2(n_455),
.B1(n_472),
.B2(n_457),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_769),
.A2(n_810),
.B(n_808),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_807),
.B(n_524),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_810),
.A2(n_560),
.B(n_547),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_806),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_763),
.A2(n_650),
.B(n_651),
.C(n_647),
.Y(n_857)
);

INVx3_ASAP7_75t_SL g858 ( 
.A(n_800),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_772),
.B(n_557),
.Y(n_859)
);

BUFx12f_ASAP7_75t_L g860 ( 
.A(n_788),
.Y(n_860)
);

BUFx12f_ASAP7_75t_L g861 ( 
.A(n_788),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_772),
.B(n_570),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_822),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_SL g864 ( 
.A1(n_812),
.A2(n_564),
.B(n_569),
.C(n_565),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_774),
.A2(n_653),
.B1(n_678),
.B2(n_666),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_780),
.B(n_687),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_762),
.A2(n_572),
.B(n_571),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_766),
.A2(n_577),
.B(n_574),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_788),
.B(n_679),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_813),
.A2(n_584),
.B(n_579),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_765),
.B(n_809),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_767),
.B(n_582),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_813),
.A2(n_589),
.B(n_587),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_793),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_784),
.B(n_436),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_764),
.Y(n_876)
);

AO32x2_ASAP7_75t_L g877 ( 
.A1(n_756),
.A2(n_522),
.A3(n_680),
.B1(n_754),
.B2(n_749),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_764),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_776),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_817),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_818),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_760),
.B(n_437),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_784),
.B(n_776),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_791),
.B(n_441),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_824),
.B(n_590),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_803),
.A2(n_599),
.B(n_598),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_758),
.B(n_443),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_803),
.A2(n_605),
.B(n_601),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_779),
.A2(n_773),
.B1(n_761),
.B2(n_823),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_SL g890 ( 
.A1(n_799),
.A2(n_609),
.B(n_610),
.C(n_608),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_779),
.A2(n_444),
.B1(n_451),
.B2(n_450),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_819),
.A2(n_511),
.B(n_516),
.C(n_435),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_799),
.A2(n_550),
.B(n_519),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_775),
.B(n_459),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_820),
.B(n_28),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_804),
.A2(n_465),
.B1(n_466),
.B2(n_461),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_825),
.A2(n_477),
.B1(n_478),
.B2(n_473),
.Y(n_897)
);

NOR3xp33_ASAP7_75t_L g898 ( 
.A(n_815),
.B(n_481),
.C(n_480),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_811),
.Y(n_899)
);

BUFx4f_ASAP7_75t_L g900 ( 
.A(n_775),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_811),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_775),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_775),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_821),
.A2(n_487),
.B(n_484),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_SL g905 ( 
.A(n_805),
.B(n_492),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_782),
.A2(n_501),
.B(n_493),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_782),
.A2(n_506),
.B(n_503),
.Y(n_907)
);

AOI32xp33_ASAP7_75t_L g908 ( 
.A1(n_796),
.A2(n_542),
.A3(n_543),
.B1(n_533),
.B2(n_508),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_789),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_782),
.A2(n_552),
.B(n_544),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_795),
.B(n_562),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_814),
.Y(n_912)
);

NOR2x1_ASAP7_75t_L g913 ( 
.A(n_805),
.B(n_580),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_790),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_795),
.B(n_575),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_790),
.A2(n_593),
.B1(n_591),
.B2(n_586),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_786),
.B(n_33),
.Y(n_917)
);

OR2x6_ASAP7_75t_SL g918 ( 
.A(n_796),
.B(n_33),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_805),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_790),
.A2(n_36),
.B(n_34),
.C(n_35),
.Y(n_920)
);

INVxp67_ASAP7_75t_SL g921 ( 
.A(n_789),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_790),
.A2(n_37),
.B(n_34),
.C(n_35),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_786),
.A2(n_538),
.B1(n_586),
.B2(n_580),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_787),
.B(n_626),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_763),
.A2(n_586),
.B1(n_631),
.B2(n_626),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_786),
.B(n_38),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_786),
.A2(n_538),
.B1(n_631),
.B2(n_626),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_804),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_763),
.A2(n_631),
.B1(n_663),
.B2(n_660),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_814),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_805),
.B(n_38),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_769),
.A2(n_660),
.B(n_663),
.C(n_631),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_782),
.A2(n_663),
.B(n_660),
.Y(n_933)
);

INVx8_ASAP7_75t_L g934 ( 
.A(n_843),
.Y(n_934)
);

CKINVDCx8_ASAP7_75t_R g935 ( 
.A(n_903),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_853),
.A2(n_674),
.B(n_667),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_826),
.A2(n_538),
.B(n_142),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_839),
.B(n_39),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_SL g939 ( 
.A1(n_828),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_939)
);

INVxp67_ASAP7_75t_SL g940 ( 
.A(n_919),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_859),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_841),
.A2(n_674),
.B(n_667),
.Y(n_942)
);

OA21x2_ASAP7_75t_L g943 ( 
.A1(n_842),
.A2(n_538),
.B(n_667),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_845),
.Y(n_944)
);

OAI21xp33_ASAP7_75t_SL g945 ( 
.A1(n_917),
.A2(n_42),
.B(n_43),
.Y(n_945)
);

BUFx2_ASAP7_75t_SL g946 ( 
.A(n_847),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_833),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_932),
.A2(n_145),
.B(n_143),
.Y(n_948)
);

AO32x2_ASAP7_75t_L g949 ( 
.A1(n_889),
.A2(n_46),
.A3(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_926),
.A2(n_695),
.B1(n_698),
.B2(n_676),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_856),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_833),
.Y(n_952)
);

AO31x2_ASAP7_75t_L g953 ( 
.A1(n_848),
.A2(n_695),
.A3(n_698),
.B(n_676),
.Y(n_953)
);

AO31x2_ASAP7_75t_L g954 ( 
.A1(n_886),
.A2(n_698),
.A3(n_695),
.B(n_49),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_831),
.A2(n_49),
.B(n_45),
.C(n_47),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_888),
.A2(n_830),
.B(n_908),
.C(n_923),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_878),
.B(n_50),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_862),
.A2(n_854),
.B(n_900),
.C(n_868),
.Y(n_958)
);

BUFx12f_ASAP7_75t_L g959 ( 
.A(n_860),
.Y(n_959)
);

OAI21x1_ASAP7_75t_L g960 ( 
.A1(n_837),
.A2(n_148),
.B(n_146),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_911),
.A2(n_152),
.B(n_150),
.Y(n_961)
);

OAI22xp33_ASAP7_75t_L g962 ( 
.A1(n_918),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_905),
.B(n_51),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_858),
.Y(n_964)
);

AOI31xp67_ASAP7_75t_L g965 ( 
.A1(n_927),
.A2(n_158),
.A3(n_159),
.B(n_154),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_846),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_857),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_915),
.A2(n_166),
.B(n_160),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_840),
.A2(n_169),
.B(n_168),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_861),
.B(n_53),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_844),
.B(n_54),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_900),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_885),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_849),
.B(n_59),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_880),
.B(n_60),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_876),
.B(n_61),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_881),
.Y(n_977)
);

CKINVDCx9p33_ASAP7_75t_R g978 ( 
.A(n_894),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_863),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_846),
.Y(n_980)
);

OA21x2_ASAP7_75t_L g981 ( 
.A1(n_933),
.A2(n_174),
.B(n_172),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_912),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_924),
.A2(n_176),
.B(n_175),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_930),
.B(n_61),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_893),
.A2(n_179),
.B(n_178),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_871),
.B(n_62),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_866),
.B(n_62),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_827),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_899),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_879),
.B(n_63),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_870),
.A2(n_183),
.B(n_181),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_895),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_829),
.A2(n_185),
.B(n_184),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_SL g994 ( 
.A1(n_885),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_850),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_906),
.A2(n_187),
.B(n_186),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_907),
.A2(n_189),
.B(n_188),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_873),
.A2(n_193),
.B(n_192),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_867),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_850),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_827),
.Y(n_1001)
);

OAI22x1_ASAP7_75t_L g1002 ( 
.A1(n_931),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_SL g1003 ( 
.A1(n_902),
.A2(n_200),
.B(n_197),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_827),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_874),
.B(n_883),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_835),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_832),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_SL g1008 ( 
.A1(n_890),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_872),
.B(n_74),
.Y(n_1009)
);

OAI21x1_ASAP7_75t_L g1010 ( 
.A1(n_929),
.A2(n_207),
.B(n_206),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_851),
.B(n_75),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_910),
.A2(n_209),
.B(n_208),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_869),
.B(n_75),
.Y(n_1013)
);

AO31x2_ASAP7_75t_L g1014 ( 
.A1(n_892),
.A2(n_79),
.A3(n_76),
.B(n_77),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_855),
.A2(n_213),
.B(n_212),
.Y(n_1015)
);

OA21x2_ASAP7_75t_L g1016 ( 
.A1(n_925),
.A2(n_215),
.B(n_214),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_851),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_928),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_875),
.A2(n_218),
.B(n_216),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_SL g1020 ( 
.A1(n_882),
.A2(n_81),
.B(n_77),
.C(n_80),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_909),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_1021)
);

OAI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_869),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1022)
);

OAI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_891),
.A2(n_86),
.B1(n_83),
.B2(n_84),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_887),
.A2(n_221),
.B(n_220),
.Y(n_1024)
);

CKINVDCx8_ASAP7_75t_R g1025 ( 
.A(n_928),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_852),
.A2(n_89),
.B1(n_86),
.B2(n_88),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_901),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_921),
.A2(n_228),
.B(n_224),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_884),
.A2(n_230),
.B(n_229),
.Y(n_1029)
);

AOI221x1_ASAP7_75t_L g1030 ( 
.A1(n_916),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.C(n_92),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_901),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_877),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_865),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_913),
.Y(n_1034)
);

NOR2x1_ASAP7_75t_SL g1035 ( 
.A(n_896),
.B(n_233),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_904),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_834),
.B(n_90),
.Y(n_1037)
);

AOI211x1_ASAP7_75t_L g1038 ( 
.A1(n_897),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_864),
.A2(n_239),
.B(n_238),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_914),
.B(n_93),
.Y(n_1040)
);

AO32x2_ASAP7_75t_L g1041 ( 
.A1(n_877),
.A2(n_94),
.A3(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_898),
.B(n_96),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_877),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_920),
.A2(n_97),
.B(n_98),
.C(n_99),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_922),
.A2(n_243),
.B(n_241),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_853),
.A2(n_245),
.B(n_244),
.Y(n_1046)
);

OA21x2_ASAP7_75t_L g1047 ( 
.A1(n_842),
.A2(n_248),
.B(n_247),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_839),
.B(n_98),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_847),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_SL g1050 ( 
.A1(n_828),
.A2(n_99),
.B(n_100),
.C(n_101),
.Y(n_1050)
);

AO21x2_ASAP7_75t_L g1051 ( 
.A1(n_888),
.A2(n_250),
.B(n_249),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_847),
.Y(n_1052)
);

BUFx8_ASAP7_75t_L g1053 ( 
.A(n_843),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_826),
.A2(n_254),
.B(n_252),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_853),
.A2(n_256),
.B(n_255),
.Y(n_1055)
);

AOI21x1_ASAP7_75t_L g1056 ( 
.A1(n_848),
.A2(n_259),
.B(n_258),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_831),
.A2(n_100),
.B(n_102),
.C(n_103),
.Y(n_1057)
);

AOI21xp33_ASAP7_75t_L g1058 ( 
.A1(n_908),
.A2(n_103),
.B(n_104),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_853),
.A2(n_261),
.B(n_260),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_826),
.A2(n_263),
.B(n_262),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_853),
.A2(n_266),
.B(n_264),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_831),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_917),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_838),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_860),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_847),
.Y(n_1066)
);

NAND2x1_ASAP7_75t_L g1067 ( 
.A(n_835),
.B(n_276),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_919),
.B(n_108),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_917),
.A2(n_109),
.B(n_110),
.C(n_111),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_853),
.A2(n_279),
.B(n_278),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_838),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_839),
.B(n_112),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_839),
.B(n_115),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_919),
.B(n_116),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_919),
.Y(n_1075)
);

INVx1_ASAP7_75t_SL g1076 ( 
.A(n_919),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_836),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_853),
.A2(n_281),
.B(n_280),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_839),
.B(n_117),
.Y(n_1079)
);

INVx5_ASAP7_75t_L g1080 ( 
.A(n_860),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_853),
.A2(n_284),
.B(n_283),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_831),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_919),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_853),
.A2(n_286),
.B(n_285),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_826),
.A2(n_344),
.B(n_421),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_838),
.B(n_118),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_847),
.B(n_120),
.Y(n_1087)
);

INVx3_ASAP7_75t_SL g1088 ( 
.A(n_858),
.Y(n_1088)
);

BUFx10_ASAP7_75t_L g1089 ( 
.A(n_846),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_SL g1090 ( 
.A1(n_888),
.A2(n_346),
.B(n_420),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_1075),
.Y(n_1091)
);

INVx5_ASAP7_75t_L g1092 ( 
.A(n_964),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_977),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_1083),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1049),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_1095)
);

BUFx8_ASAP7_75t_L g1096 ( 
.A(n_964),
.Y(n_1096)
);

AOI221xp5_ASAP7_75t_L g1097 ( 
.A1(n_1058),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.C(n_125),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_982),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_L g1099 ( 
.A1(n_942),
.A2(n_347),
.B(n_419),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_934),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_959),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_944),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_956),
.A2(n_958),
.B(n_938),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1048),
.A2(n_124),
.B(n_126),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_1088),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1066),
.B(n_126),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_967),
.A2(n_349),
.B(n_418),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_1076),
.B(n_287),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_946),
.B(n_127),
.Y(n_1109)
);

AOI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1056),
.A2(n_350),
.B(n_416),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1052),
.B(n_128),
.Y(n_1111)
);

OA21x2_ASAP7_75t_L g1112 ( 
.A1(n_948),
.A2(n_341),
.B(n_413),
.Y(n_1112)
);

INVx3_ASAP7_75t_SL g1113 ( 
.A(n_934),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_963),
.A2(n_128),
.B(n_129),
.C(n_130),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_986),
.B(n_131),
.Y(n_1115)
);

BUFx8_ASAP7_75t_L g1116 ( 
.A(n_1074),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_1061),
.A2(n_340),
.B(n_411),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_SL g1118 ( 
.A1(n_1070),
.A2(n_131),
.B(n_132),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_951),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_966),
.B(n_133),
.Y(n_1120)
);

AO21x2_ASAP7_75t_L g1121 ( 
.A1(n_1084),
.A2(n_338),
.B(n_409),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1025),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_SL g1123 ( 
.A1(n_1035),
.A2(n_133),
.B(n_134),
.Y(n_1123)
);

AO21x1_ASAP7_75t_SL g1124 ( 
.A1(n_1071),
.A2(n_134),
.B(n_135),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1053),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1074),
.B(n_135),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_SL g1127 ( 
.A1(n_1024),
.A2(n_288),
.B(n_290),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1072),
.A2(n_1079),
.B(n_1073),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1000),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_1129)
);

INVx4_ASAP7_75t_L g1130 ( 
.A(n_947),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1036),
.A2(n_1055),
.B(n_1046),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1077),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_980),
.B(n_296),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_1043),
.A2(n_297),
.A3(n_300),
.B(n_302),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1059),
.A2(n_304),
.B(n_305),
.Y(n_1135)
);

OA21x2_ASAP7_75t_L g1136 ( 
.A1(n_1085),
.A2(n_306),
.B(n_307),
.Y(n_1136)
);

NAND3xp33_ASAP7_75t_L g1137 ( 
.A(n_1063),
.B(n_308),
.C(n_311),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_952),
.Y(n_1138)
);

OA21x2_ASAP7_75t_L g1139 ( 
.A1(n_960),
.A2(n_312),
.B(n_318),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_988),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1086),
.A2(n_320),
.B1(n_323),
.B2(n_324),
.Y(n_1141)
);

BUFx10_ASAP7_75t_L g1142 ( 
.A(n_1042),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1078),
.A2(n_325),
.B(n_326),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1081),
.A2(n_328),
.B(n_330),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_995),
.B(n_333),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_979),
.A2(n_335),
.B1(n_336),
.B2(n_353),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_1065),
.B(n_355),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_976),
.B(n_357),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1087),
.B(n_1005),
.Y(n_1149)
);

OR2x6_ASAP7_75t_L g1150 ( 
.A(n_1068),
.B(n_358),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_940),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_989),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_SL g1153 ( 
.A1(n_974),
.A2(n_984),
.B(n_975),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_987),
.Y(n_1154)
);

OR2x2_ASAP7_75t_L g1155 ( 
.A(n_992),
.B(n_360),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1011),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_988),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1068),
.B(n_423),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_985),
.A2(n_361),
.B(n_362),
.Y(n_1159)
);

NAND2x1p5_ASAP7_75t_L g1160 ( 
.A(n_1080),
.B(n_363),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_957),
.B(n_366),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1031),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1009),
.B(n_368),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1006),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_943),
.A2(n_1010),
.B(n_1015),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_971),
.B(n_369),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_990),
.Y(n_1167)
);

AOI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_962),
.A2(n_373),
.B1(n_374),
.B2(n_378),
.C(n_379),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_1045),
.A2(n_380),
.A3(n_384),
.B(n_385),
.Y(n_1169)
);

BUFx8_ASAP7_75t_SL g1170 ( 
.A(n_970),
.Y(n_1170)
);

INVx2_ASAP7_75t_SL g1171 ( 
.A(n_1080),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1017),
.A2(n_395),
.B1(n_396),
.B2(n_399),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1080),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1018),
.B(n_401),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_996),
.A2(n_405),
.B(n_406),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1033),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1027),
.B(n_407),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_997),
.A2(n_1012),
.B(n_1090),
.Y(n_1178)
);

OR2x6_ASAP7_75t_L g1179 ( 
.A(n_970),
.B(n_1001),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_978),
.Y(n_1180)
);

OR3x4_ASAP7_75t_SL g1181 ( 
.A(n_1022),
.B(n_1002),
.C(n_1013),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1089),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1040),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_SL g1184 ( 
.A1(n_961),
.A2(n_968),
.B(n_1019),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1004),
.B(n_935),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_991),
.A2(n_998),
.B(n_1067),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1027),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1037),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1064),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_SL g1190 ( 
.A1(n_1029),
.A2(n_1082),
.B(n_1057),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_953),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_983),
.A2(n_1028),
.B(n_993),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1027),
.B(n_994),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_973),
.B(n_1034),
.Y(n_1194)
);

OAI21xp33_ASAP7_75t_L g1195 ( 
.A1(n_945),
.A2(n_1069),
.B(n_1026),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1047),
.A2(n_981),
.B(n_1039),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_941),
.Y(n_1197)
);

BUFx2_ASAP7_75t_R g1198 ( 
.A(n_1051),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1021),
.Y(n_1199)
);

OA21x2_ASAP7_75t_L g1200 ( 
.A1(n_950),
.A2(n_1030),
.B(n_1007),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_999),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_SL g1202 ( 
.A1(n_955),
.A2(n_1062),
.B(n_1044),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1014),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1032),
.B(n_1023),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_939),
.A2(n_1050),
.B(n_1008),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_972),
.A2(n_1038),
.B1(n_1032),
.B2(n_1016),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1014),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1020),
.B(n_954),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_953),
.A2(n_954),
.A3(n_965),
.B(n_1041),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1016),
.A2(n_981),
.B(n_1003),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1014),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_954),
.B(n_953),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1041),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_949),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_949),
.B(n_1041),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_949),
.B(n_919),
.Y(n_1216)
);

BUFx8_ASAP7_75t_L g1217 ( 
.A(n_964),
.Y(n_1217)
);

NOR2x1_ASAP7_75t_R g1218 ( 
.A(n_947),
.B(n_783),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1083),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_977),
.B(n_838),
.Y(n_1220)
);

OA21x2_ASAP7_75t_L g1221 ( 
.A1(n_937),
.A2(n_936),
.B(n_942),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_958),
.A2(n_782),
.B(n_828),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_977),
.B(n_838),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_937),
.A2(n_1060),
.B(n_1054),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_1083),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1035),
.A2(n_1084),
.B(n_1070),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1075),
.B(n_847),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_964),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_1066),
.Y(n_1229)
);

OR2x2_ASAP7_75t_L g1230 ( 
.A(n_1049),
.B(n_805),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_937),
.A2(n_1060),
.B(n_1054),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_977),
.B(n_838),
.Y(n_1232)
);

AO21x2_ASAP7_75t_L g1233 ( 
.A1(n_942),
.A2(n_888),
.B(n_969),
.Y(n_1233)
);

AO222x2_ASAP7_75t_L g1234 ( 
.A1(n_1013),
.A2(n_615),
.B1(n_617),
.B2(n_627),
.C1(n_677),
.C2(n_668),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1049),
.B(n_847),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_937),
.A2(n_1060),
.B(n_1054),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_977),
.B(n_838),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_956),
.A2(n_926),
.B(n_917),
.C(n_838),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1238),
.B(n_1220),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1093),
.Y(n_1240)
);

OA21x2_ASAP7_75t_L g1241 ( 
.A1(n_1196),
.A2(n_1212),
.B(n_1103),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1189),
.A2(n_1195),
.B1(n_1197),
.B2(n_1115),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1161),
.A2(n_1097),
.B1(n_1199),
.B2(n_1202),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1223),
.B(n_1232),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1211),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1098),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1208),
.A2(n_1207),
.B(n_1191),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1226),
.A2(n_1153),
.B(n_1128),
.Y(n_1248)
);

INVxp67_ASAP7_75t_L g1249 ( 
.A(n_1230),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1102),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1216),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1132),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1096),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1216),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1119),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1152),
.Y(n_1256)
);

AO21x2_ASAP7_75t_L g1257 ( 
.A1(n_1153),
.A2(n_1165),
.B(n_1233),
.Y(n_1257)
);

AO21x2_ASAP7_75t_L g1258 ( 
.A1(n_1127),
.A2(n_1131),
.B(n_1118),
.Y(n_1258)
);

OA21x2_ASAP7_75t_L g1259 ( 
.A1(n_1224),
.A2(n_1236),
.B(n_1231),
.Y(n_1259)
);

AO21x2_ASAP7_75t_L g1260 ( 
.A1(n_1127),
.A2(n_1118),
.B(n_1184),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1234),
.B(n_1149),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_1122),
.B(n_1179),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1235),
.B(n_1229),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1126),
.B(n_1111),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1176),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1164),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1237),
.B(n_1183),
.Y(n_1267)
);

INVx8_ASAP7_75t_L g1268 ( 
.A(n_1092),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1203),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1142),
.B(n_1150),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1162),
.Y(n_1271)
);

OAI21xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1104),
.A2(n_1215),
.B(n_1166),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1225),
.B(n_1094),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1096),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1106),
.B(n_1151),
.Y(n_1275)
);

AO21x2_ASAP7_75t_L g1276 ( 
.A1(n_1184),
.A2(n_1178),
.B(n_1205),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1194),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1206),
.A2(n_1190),
.B(n_1188),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1142),
.B(n_1150),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1222),
.A2(n_1192),
.B(n_1186),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1155),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1154),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1219),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1092),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1116),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1217),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1120),
.Y(n_1287)
);

INVx3_ASAP7_75t_SL g1288 ( 
.A(n_1113),
.Y(n_1288)
);

OR2x6_ASAP7_75t_L g1289 ( 
.A(n_1177),
.B(n_1193),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1163),
.B(n_1227),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1133),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1109),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1140),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1145),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1201),
.A2(n_1137),
.B(n_1156),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1204),
.B(n_1202),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1140),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1157),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1187),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1147),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1217),
.Y(n_1301)
);

AO21x2_ASAP7_75t_L g1302 ( 
.A1(n_1121),
.A2(n_1175),
.B(n_1099),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1091),
.B(n_1167),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1147),
.Y(n_1304)
);

INVx2_ASAP7_75t_SL g1305 ( 
.A(n_1105),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1138),
.B(n_1185),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1174),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1182),
.B(n_1130),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1125),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1167),
.B(n_1158),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1108),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1180),
.B(n_1228),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1160),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1148),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1116),
.Y(n_1315)
);

BUFx8_ASAP7_75t_SL g1316 ( 
.A(n_1170),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1100),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1095),
.B(n_1124),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1200),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1114),
.B(n_1101),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1214),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1213),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1200),
.B(n_1168),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1123),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1218),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1171),
.B(n_1173),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1209),
.B(n_1181),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1123),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1141),
.A2(n_1143),
.B(n_1144),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1112),
.B(n_1117),
.Y(n_1330)
);

NAND4xp25_ASAP7_75t_L g1331 ( 
.A(n_1146),
.B(n_1129),
.C(n_1135),
.D(n_1172),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1198),
.A2(n_1136),
.B1(n_1139),
.B2(n_1107),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1110),
.B(n_1159),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1221),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1134),
.B(n_1169),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1235),
.B(n_1230),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1212),
.A2(n_1210),
.B(n_1196),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1212),
.A2(n_1210),
.B(n_1196),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1211),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1235),
.B(n_847),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1240),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1340),
.B(n_1263),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1246),
.Y(n_1343)
);

INVxp67_ASAP7_75t_SL g1344 ( 
.A(n_1245),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1264),
.B(n_1261),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1261),
.B(n_1336),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1296),
.B(n_1275),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1268),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1244),
.B(n_1267),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1296),
.B(n_1249),
.Y(n_1350)
);

OAI221xp5_ASAP7_75t_L g1351 ( 
.A1(n_1243),
.A2(n_1242),
.B1(n_1272),
.B2(n_1331),
.C(n_1292),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1244),
.B(n_1267),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1322),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1249),
.B(n_1327),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1310),
.B(n_1320),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1242),
.A2(n_1243),
.B1(n_1318),
.B2(n_1304),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1278),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1265),
.B(n_1252),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1247),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1256),
.B(n_1266),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1271),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1273),
.B(n_1282),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1303),
.B(n_1270),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1262),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1279),
.B(n_1287),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1281),
.B(n_1283),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1245),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1239),
.A2(n_1294),
.B1(n_1277),
.B2(n_1331),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1285),
.B(n_1315),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1239),
.B(n_1300),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1277),
.B(n_1251),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1250),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1339),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1339),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1316),
.Y(n_1375)
);

NAND2x1_ASAP7_75t_L g1376 ( 
.A(n_1313),
.B(n_1295),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1255),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1319),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1278),
.Y(n_1379)
);

OR2x2_ASAP7_75t_L g1380 ( 
.A(n_1251),
.B(n_1254),
.Y(n_1380)
);

OR2x6_ASAP7_75t_L g1381 ( 
.A(n_1289),
.B(n_1268),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1284),
.B(n_1293),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1306),
.B(n_1291),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1268),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1293),
.B(n_1297),
.Y(n_1385)
);

AOI222xp33_ASAP7_75t_L g1386 ( 
.A1(n_1272),
.A2(n_1323),
.B1(n_1314),
.B2(n_1295),
.C1(n_1254),
.C2(n_1325),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1306),
.B(n_1290),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1297),
.B(n_1299),
.Y(n_1388)
);

BUFx3_ASAP7_75t_L g1389 ( 
.A(n_1308),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1311),
.A2(n_1329),
.B(n_1307),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1298),
.B(n_1305),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1248),
.B(n_1328),
.Y(n_1392)
);

OR2x6_ASAP7_75t_L g1393 ( 
.A(n_1269),
.B(n_1286),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1321),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1319),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1308),
.B(n_1317),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1253),
.B(n_1274),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1241),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1312),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1248),
.B(n_1324),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1301),
.B(n_1288),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1326),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1288),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1257),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1325),
.B(n_1309),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1335),
.B(n_1323),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1332),
.B(n_1257),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1406),
.B(n_1334),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1342),
.B(n_1334),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1367),
.B(n_1338),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1349),
.B(n_1276),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1367),
.Y(n_1412)
);

INVxp67_ASAP7_75t_SL g1413 ( 
.A(n_1344),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1373),
.B(n_1374),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1359),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1392),
.B(n_1260),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1352),
.B(n_1276),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1373),
.B(n_1337),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1394),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1353),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1347),
.B(n_1350),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1362),
.B(n_1260),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1370),
.B(n_1332),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1341),
.B(n_1258),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1343),
.B(n_1258),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1353),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1354),
.B(n_1330),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1395),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1400),
.B(n_1330),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1400),
.B(n_1280),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1400),
.B(n_1355),
.Y(n_1431)
);

BUFx2_ASAP7_75t_SL g1432 ( 
.A(n_1389),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1393),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1378),
.B(n_1259),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1399),
.Y(n_1435)
);

OR2x2_ASAP7_75t_L g1436 ( 
.A(n_1380),
.B(n_1302),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1396),
.B(n_1316),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1412),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1416),
.B(n_1393),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1409),
.B(n_1407),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1414),
.B(n_1371),
.Y(n_1441)
);

NAND2x1p5_ASAP7_75t_L g1442 ( 
.A(n_1410),
.B(n_1376),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1414),
.B(n_1398),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1409),
.B(n_1368),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1408),
.B(n_1407),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1419),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_SL g1447 ( 
.A(n_1432),
.B(n_1381),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1415),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1408),
.B(n_1357),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1435),
.B(n_1368),
.Y(n_1450)
);

NAND2x1_ASAP7_75t_L g1451 ( 
.A(n_1416),
.B(n_1390),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1431),
.B(n_1357),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1431),
.B(n_1379),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1421),
.B(n_1370),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1424),
.B(n_1379),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1433),
.Y(n_1456)
);

CKINVDCx16_ASAP7_75t_R g1457 ( 
.A(n_1437),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1413),
.B(n_1366),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1424),
.B(n_1404),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1419),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1427),
.B(n_1358),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1427),
.B(n_1410),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1425),
.B(n_1404),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1420),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1425),
.B(n_1363),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1411),
.B(n_1360),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1417),
.B(n_1386),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1420),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1426),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1433),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1422),
.B(n_1402),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1428),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1465),
.B(n_1430),
.Y(n_1473)
);

NOR2xp67_ASAP7_75t_L g1474 ( 
.A(n_1438),
.B(n_1403),
.Y(n_1474)
);

NOR2x1_ASAP7_75t_L g1475 ( 
.A(n_1450),
.B(n_1403),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1446),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1460),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1472),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1472),
.Y(n_1479)
);

INVx2_ASAP7_75t_SL g1480 ( 
.A(n_1456),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1448),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1441),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1465),
.B(n_1430),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1462),
.B(n_1436),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1441),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1464),
.Y(n_1486)
);

AO22x1_ASAP7_75t_L g1487 ( 
.A1(n_1439),
.A2(n_1423),
.B1(n_1365),
.B2(n_1369),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1468),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1469),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1467),
.A2(n_1351),
.B(n_1356),
.C(n_1345),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1461),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1461),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1443),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1443),
.Y(n_1494)
);

OAI211xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1458),
.A2(n_1387),
.B(n_1329),
.C(n_1383),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1492),
.B(n_1440),
.Y(n_1496)
);

OAI31xp33_ASAP7_75t_L g1497 ( 
.A1(n_1490),
.A2(n_1346),
.A3(n_1444),
.B(n_1471),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1494),
.B(n_1440),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_SL g1499 ( 
.A(n_1475),
.B(n_1457),
.Y(n_1499)
);

NAND2xp33_ASAP7_75t_SL g1500 ( 
.A(n_1480),
.B(n_1375),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1494),
.B(n_1445),
.Y(n_1501)
);

OAI221xp5_ASAP7_75t_L g1502 ( 
.A1(n_1490),
.A2(n_1466),
.B1(n_1454),
.B2(n_1462),
.C(n_1470),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_L g1503 ( 
.A(n_1495),
.B(n_1493),
.C(n_1474),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1481),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1478),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1480),
.B(n_1401),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1482),
.B(n_1445),
.Y(n_1507)
);

AOI32xp33_ASAP7_75t_L g1508 ( 
.A1(n_1473),
.A2(n_1449),
.A3(n_1452),
.B1(n_1453),
.B2(n_1455),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1487),
.A2(n_1455),
.B1(n_1459),
.B2(n_1463),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1479),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1476),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1477),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1473),
.B(n_1449),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1500),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1505),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1502),
.A2(n_1491),
.B1(n_1485),
.B2(n_1486),
.C(n_1488),
.Y(n_1516)
);

AOI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1497),
.A2(n_1489),
.B1(n_1483),
.B2(n_1452),
.C(n_1453),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1503),
.A2(n_1483),
.B1(n_1484),
.B2(n_1459),
.C(n_1463),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1499),
.A2(n_1439),
.B1(n_1451),
.B2(n_1429),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1500),
.A2(n_1447),
.B(n_1451),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1517),
.A2(n_1509),
.B(n_1506),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1516),
.A2(n_1518),
.B1(n_1519),
.B2(n_1439),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1514),
.B(n_1513),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1520),
.A2(n_1508),
.B(n_1506),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1515),
.B(n_1375),
.Y(n_1525)
);

NOR2x1_ASAP7_75t_L g1526 ( 
.A(n_1524),
.B(n_1405),
.Y(n_1526)
);

NOR3xp33_ASAP7_75t_L g1527 ( 
.A(n_1521),
.B(n_1391),
.C(n_1397),
.Y(n_1527)
);

AOI211xp5_ASAP7_75t_L g1528 ( 
.A1(n_1522),
.A2(n_1501),
.B(n_1498),
.C(n_1512),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_L g1529 ( 
.A(n_1525),
.B(n_1389),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1523),
.A2(n_1511),
.B(n_1496),
.Y(n_1530)
);

NAND3xp33_ASAP7_75t_SL g1531 ( 
.A(n_1524),
.B(n_1442),
.C(n_1507),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1527),
.B(n_1510),
.Y(n_1532)
);

NOR3xp33_ASAP7_75t_L g1533 ( 
.A(n_1531),
.B(n_1382),
.C(n_1384),
.Y(n_1533)
);

NOR3xp33_ASAP7_75t_L g1534 ( 
.A(n_1526),
.B(n_1384),
.C(n_1388),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1532),
.B(n_1530),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1534),
.B(n_1528),
.Y(n_1536)
);

NOR2xp67_ASAP7_75t_SL g1537 ( 
.A(n_1535),
.B(n_1348),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1537),
.B(n_1536),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1538),
.Y(n_1539)
);

NAND3xp33_ASAP7_75t_L g1540 ( 
.A(n_1538),
.B(n_1533),
.C(n_1529),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_SL g1541 ( 
.A1(n_1539),
.A2(n_1348),
.B1(n_1393),
.B2(n_1381),
.Y(n_1541)
);

NAND2xp33_ASAP7_75t_SL g1542 ( 
.A(n_1540),
.B(n_1434),
.Y(n_1542)
);

OAI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1542),
.A2(n_1385),
.B(n_1418),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1541),
.B(n_1361),
.C(n_1364),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1543),
.A2(n_1333),
.B(n_1504),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1545),
.A2(n_1544),
.B1(n_1372),
.B2(n_1377),
.Y(n_1546)
);


endmodule