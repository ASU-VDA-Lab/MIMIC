module fake_jpeg_3435_n_442 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_442);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_442;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_44),
.B(n_71),
.Y(n_91)
);

INVx2_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_45),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_9),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_72),
.Y(n_117)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_16),
.B(n_9),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_7),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_85),
.Y(n_93)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_19),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_45),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_18),
.B1(n_20),
.B2(n_36),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_115),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_29),
.B1(n_20),
.B2(n_22),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_61),
.A2(n_27),
.B1(n_19),
.B2(n_20),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_47),
.A2(n_27),
.B1(n_19),
.B2(n_20),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_58),
.A2(n_29),
.B1(n_27),
.B2(n_21),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_133),
.B1(n_39),
.B2(n_24),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_22),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_27),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_46),
.A2(n_21),
.B1(n_37),
.B2(n_36),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_131),
.A2(n_39),
.B(n_33),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_48),
.A2(n_17),
.B1(n_28),
.B2(n_35),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_143),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_82),
.B1(n_59),
.B2(n_69),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_145),
.B1(n_148),
.B2(n_152),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_17),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_149),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_76),
.B1(n_62),
.B2(n_60),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_172),
.B1(n_115),
.B2(n_92),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_142),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_37),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_35),
.B1(n_28),
.B2(n_27),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_100),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_146),
.B(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_28),
.B1(n_27),
.B2(n_68),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_97),
.B(n_0),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_110),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_126),
.A2(n_51),
.B1(n_57),
.B2(n_39),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_153),
.B(n_155),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_39),
.B(n_24),
.C(n_2),
.Y(n_154)
);

AO22x1_ASAP7_75t_L g212 ( 
.A1(n_154),
.A2(n_92),
.B1(n_98),
.B2(n_106),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_93),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_88),
.B(n_0),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_1),
.Y(n_195)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_167),
.Y(n_198)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_87),
.B(n_0),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_164),
.Y(n_191)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_29),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_174),
.Y(n_185)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_94),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_87),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_0),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_24),
.Y(n_211)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_176),
.Y(n_210)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_177),
.B(n_179),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_132),
.A2(n_39),
.B1(n_24),
.B2(n_3),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_134),
.B1(n_101),
.B2(n_113),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_182),
.A2(n_192),
.B1(n_194),
.B2(n_214),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_137),
.A2(n_99),
.B1(n_132),
.B2(n_118),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_99),
.B1(n_118),
.B2(n_120),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_195),
.B(n_1),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_109),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_215),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_175),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_150),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_146),
.B(n_121),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_223),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_157),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_233),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_237),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_202),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_228),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_144),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_245),
.C(n_209),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_139),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_183),
.A2(n_153),
.B(n_144),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_241),
.B(n_212),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_175),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_140),
.B1(n_154),
.B2(n_162),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_236),
.B1(n_240),
.B2(n_204),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_182),
.A2(n_162),
.B1(n_177),
.B2(n_174),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_163),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

OA22x2_ASAP7_75t_L g239 ( 
.A1(n_194),
.A2(n_178),
.B1(n_151),
.B2(n_171),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_239),
.A2(n_242),
.B1(n_142),
.B2(n_188),
.Y(n_280)
);

A2O1A1O1Ixp25_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_147),
.B(n_166),
.C(n_169),
.D(n_161),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_156),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_244),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_167),
.C(n_158),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_176),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_150),
.Y(n_247)
);

OAI32xp33_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_249),
.A3(n_181),
.B1(n_188),
.B2(n_199),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_248),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_210),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_187),
.B1(n_212),
.B2(n_201),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_250),
.A2(n_252),
.B1(n_259),
.B2(n_262),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_253),
.A2(n_263),
.B(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_245),
.C(n_243),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_210),
.B1(n_206),
.B2(n_205),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_249),
.Y(n_260)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_260),
.B(n_261),
.C(n_251),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_217),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_206),
.B1(n_205),
.B2(n_191),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_232),
.A2(n_198),
.B(n_204),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_242),
.A2(n_186),
.B(n_213),
.Y(n_268)
);

OAI22x1_ASAP7_75t_SL g270 ( 
.A1(n_231),
.A2(n_242),
.B1(n_239),
.B2(n_246),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g298 ( 
.A1(n_270),
.A2(n_239),
.B(n_241),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_253),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_191),
.B(n_202),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_280),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_225),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_281),
.B(n_292),
.C(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_224),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_284),
.B(n_288),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_227),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_285),
.B(n_256),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_266),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_221),
.B1(n_218),
.B2(n_237),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_289),
.A2(n_295),
.B1(n_309),
.B2(n_276),
.Y(n_335)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_291),
.Y(n_324)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_250),
.A2(n_221),
.B1(n_233),
.B2(n_239),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_278),
.B(n_220),
.Y(n_296)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_296),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_219),
.Y(n_297)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_257),
.C(n_263),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_304),
.C(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_223),
.B1(n_222),
.B2(n_230),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_301),
.A2(n_306),
.B1(n_272),
.B2(n_269),
.Y(n_316)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_302),
.Y(n_330)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_305),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_209),
.C(n_199),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

AOI21x1_ASAP7_75t_SL g334 ( 
.A1(n_307),
.A2(n_196),
.B(n_208),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_238),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_272),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_277),
.A2(n_229),
.B1(n_248),
.B2(n_160),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_308),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_325),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_281),
.B(n_271),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_321),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_318),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_280),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_319),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_323),
.B(n_329),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_287),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_289),
.B(n_251),
.Y(n_328)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_328),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_285),
.B(n_256),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_262),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_331),
.B(n_332),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_299),
.B(n_268),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_307),
.B(n_279),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_334),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_335),
.A2(n_294),
.B1(n_287),
.B2(n_309),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_337),
.B(n_314),
.Y(n_368)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_324),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_338),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_339),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_341),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_330),
.B(n_291),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_343),
.B(n_348),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_317),
.B(n_290),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_283),
.C(n_286),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_353),
.Y(n_361)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_315),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_351),
.A2(n_352),
.B1(n_355),
.B2(n_356),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_335),
.A2(n_295),
.B1(n_294),
.B2(n_298),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_283),
.C(n_298),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_305),
.C(n_303),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_329),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_326),
.A2(n_300),
.B1(n_293),
.B2(n_275),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_315),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_279),
.Y(n_357)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_357),
.B(n_323),
.C(n_333),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_318),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_313),
.B1(n_334),
.B2(n_311),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_332),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_368),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_363),
.B(n_336),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_370),
.Y(n_378)
);

BUFx24_ASAP7_75t_SL g365 ( 
.A(n_337),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_367),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_352),
.A2(n_320),
.B1(n_326),
.B2(n_327),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_371),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_344),
.A2(n_345),
.B1(n_340),
.B2(n_342),
.Y(n_372)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_372),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_324),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_373),
.B(n_375),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_311),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_276),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_377),
.C(n_350),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_273),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_SL g402 ( 
.A(n_379),
.B(n_388),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_360),
.A2(n_355),
.B1(n_353),
.B2(n_350),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_380),
.A2(n_382),
.B1(n_387),
.B2(n_134),
.Y(n_398)
);

OAI221xp5_ASAP7_75t_L g382 ( 
.A1(n_374),
.A2(n_339),
.B1(n_336),
.B2(n_357),
.C(n_338),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_7),
.Y(n_404)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_369),
.Y(n_386)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

OAI221xp5_ASAP7_75t_L g387 ( 
.A1(n_366),
.A2(n_341),
.B1(n_275),
.B2(n_273),
.C(n_196),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_377),
.B(n_208),
.C(n_141),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_375),
.A2(n_173),
.B(n_170),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_391),
.B(n_165),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_159),
.C(n_120),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_393),
.C(n_10),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_359),
.C(n_368),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_381),
.A2(n_360),
.B1(n_362),
.B2(n_369),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_401),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_383),
.A2(n_363),
.B1(n_121),
.B2(n_113),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_395),
.B(n_379),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g396 ( 
.A(n_388),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_397),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_398),
.A2(n_403),
.B1(n_11),
.B2(n_14),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_101),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_400),
.Y(n_413)
);

NOR2x1_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_39),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_378),
.A2(n_10),
.B(n_14),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_404),
.B(n_389),
.Y(n_410)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_392),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_407),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_7),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_394),
.Y(n_408)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_408),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_410),
.B(n_411),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_389),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_415),
.B(n_417),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_393),
.C(n_390),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_SL g425 ( 
.A(n_416),
.B(n_397),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_11),
.Y(n_418)
);

AOI21xp33_ASAP7_75t_L g423 ( 
.A1(n_418),
.A2(n_6),
.B(n_15),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_404),
.B(n_11),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_12),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_420),
.A2(n_422),
.B(n_423),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_416),
.A2(n_400),
.B(n_401),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_425),
.A2(n_426),
.B(n_427),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_SL g426 ( 
.A(n_409),
.B(n_6),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_408),
.A2(n_6),
.B1(n_14),
.B2(n_3),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_428),
.A2(n_412),
.B(n_414),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_429),
.A2(n_431),
.B(n_4),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_424),
.A2(n_409),
.B(n_410),
.Y(n_431)
);

O2A1O1Ixp33_ASAP7_75t_SL g432 ( 
.A1(n_421),
.A2(n_413),
.B(n_6),
.C(n_3),
.Y(n_432)
);

O2A1O1Ixp33_ASAP7_75t_SL g436 ( 
.A1(n_432),
.A2(n_4),
.B(n_13),
.C(n_15),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_421),
.Y(n_434)
);

AOI21xp33_ASAP7_75t_L g438 ( 
.A1(n_434),
.A2(n_435),
.B(n_436),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_430),
.C(n_13),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_437),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_439),
.A2(n_438),
.B(n_15),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_1),
.C(n_2),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_441),
.B(n_1),
.Y(n_442)
);


endmodule