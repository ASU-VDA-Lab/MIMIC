module real_aes_534_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_379;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_546;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
AOI222xp33_ASAP7_75t_L g152 ( .A1(n_0), .A2(n_38), .B1(n_49), .B2(n_153), .C1(n_156), .C2(n_159), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_1), .A2(n_33), .B1(n_143), .B2(n_148), .Y(n_142) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_2), .A2(n_54), .B1(n_89), .B2(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g531 ( .A1(n_3), .A2(n_17), .B1(n_532), .B2(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g533 ( .A(n_3), .Y(n_533) );
INVx1_ASAP7_75t_L g166 ( .A(n_4), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_5), .B(n_209), .Y(n_305) );
INVx1_ASAP7_75t_L g218 ( .A(n_6), .Y(n_218) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_7), .A2(n_19), .B1(n_89), .B2(n_99), .Y(n_98) );
AOI22xp33_ASAP7_75t_L g127 ( .A1(n_8), .A2(n_69), .B1(n_128), .B2(n_130), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_9), .Y(n_235) );
INVx2_ASAP7_75t_L g182 ( .A(n_10), .Y(n_182) );
INVx1_ASAP7_75t_L g314 ( .A(n_11), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g83 ( .A1(n_12), .A2(n_57), .B1(n_84), .B2(n_103), .Y(n_83) );
INVx1_ASAP7_75t_L g311 ( .A(n_13), .Y(n_311) );
INVx1_ASAP7_75t_SL g276 ( .A(n_14), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_15), .B(n_197), .Y(n_297) );
AOI33xp33_ASAP7_75t_L g247 ( .A1(n_16), .A2(n_41), .A3(n_187), .B1(n_195), .B2(n_248), .B3(n_249), .Y(n_247) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_16), .Y(n_557) );
INVx1_ASAP7_75t_L g532 ( .A(n_17), .Y(n_532) );
INVx1_ASAP7_75t_L g227 ( .A(n_18), .Y(n_227) );
OAI221xp5_ASAP7_75t_L g538 ( .A1(n_19), .A2(n_54), .B1(n_58), .B2(n_539), .C(n_541), .Y(n_538) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_20), .A2(n_71), .B(n_182), .Y(n_181) );
OR2x2_ASAP7_75t_L g210 ( .A(n_20), .B(n_71), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_21), .B(n_205), .Y(n_273) );
INVx3_ASAP7_75t_L g89 ( .A(n_22), .Y(n_89) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_23), .A2(n_32), .B1(n_136), .B2(n_139), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_24), .A2(n_520), .B1(n_521), .B2(n_522), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_24), .Y(n_520) );
INVx1_ASAP7_75t_SL g94 ( .A(n_25), .Y(n_94) );
INVx1_ASAP7_75t_L g168 ( .A(n_26), .Y(n_168) );
AND2x2_ASAP7_75t_L g203 ( .A(n_26), .B(n_166), .Y(n_203) );
AND2x2_ASAP7_75t_L g208 ( .A(n_26), .B(n_189), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_27), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_28), .B(n_205), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_29), .A2(n_180), .B1(n_209), .B2(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_30), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_31), .B(n_197), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_34), .B(n_215), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_35), .B(n_197), .Y(n_219) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_36), .A2(n_58), .B1(n_89), .B2(n_90), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_37), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g108 ( .A1(n_39), .A2(n_60), .B1(n_109), .B2(n_113), .Y(n_108) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_40), .A2(n_72), .B1(n_529), .B2(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_40), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_42), .B(n_197), .Y(n_259) );
INVx1_ASAP7_75t_L g191 ( .A(n_43), .Y(n_191) );
INVx1_ASAP7_75t_L g199 ( .A(n_43), .Y(n_199) );
AND2x2_ASAP7_75t_L g260 ( .A(n_44), .B(n_261), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g216 ( .A1(n_45), .A2(n_61), .B1(n_185), .B2(n_205), .C(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_46), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g95 ( .A(n_47), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_48), .B(n_180), .Y(n_237) );
AOI21xp5_ASAP7_75t_SL g184 ( .A1(n_50), .A2(n_185), .B(n_192), .Y(n_184) );
INVx1_ASAP7_75t_L g308 ( .A(n_51), .Y(n_308) );
INVx1_ASAP7_75t_L g258 ( .A(n_52), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_53), .A2(n_185), .B(n_257), .Y(n_256) );
INVxp33_ASAP7_75t_L g543 ( .A(n_54), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g117 ( .A1(n_55), .A2(n_66), .B1(n_118), .B2(n_122), .Y(n_117) );
INVx1_ASAP7_75t_L g189 ( .A(n_56), .Y(n_189) );
INVx1_ASAP7_75t_L g201 ( .A(n_56), .Y(n_201) );
INVxp67_ASAP7_75t_L g542 ( .A(n_58), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_59), .B(n_205), .Y(n_250) );
INVx1_ASAP7_75t_L g524 ( .A(n_61), .Y(n_524) );
AND2x2_ASAP7_75t_L g278 ( .A(n_62), .B(n_179), .Y(n_278) );
INVx1_ASAP7_75t_L g309 ( .A(n_63), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_64), .A2(n_185), .B(n_275), .Y(n_274) );
OAI22x1_ASAP7_75t_R g522 ( .A1(n_64), .A2(n_523), .B1(n_524), .B2(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g525 ( .A(n_64), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_65), .A2(n_185), .B(n_242), .C(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_67), .B(n_179), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_68), .A2(n_185), .B1(n_245), .B2(n_246), .Y(n_244) );
INVx1_ASAP7_75t_L g545 ( .A(n_68), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_68), .A2(n_537), .B1(n_546), .B2(n_552), .Y(n_551) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_70), .B(n_80), .Y(n_79) );
INVx1_ASAP7_75t_L g530 ( .A(n_72), .Y(n_530) );
INVx1_ASAP7_75t_L g193 ( .A(n_73), .Y(n_193) );
AND2x2_ASAP7_75t_L g251 ( .A(n_74), .B(n_179), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_75), .A2(n_225), .B(n_226), .C(n_229), .Y(n_224) );
BUFx2_ASAP7_75t_SL g540 ( .A(n_76), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_77), .B(n_197), .Y(n_196) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_163), .B1(n_169), .B2(n_511), .C(n_515), .Y(n_78) );
OAI222xp33_ASAP7_75t_L g515 ( .A1(n_80), .A2(n_516), .B1(n_517), .B2(n_551), .C1(n_553), .C2(n_556), .Y(n_515) );
CKINVDCx14_ASAP7_75t_R g516 ( .A(n_80), .Y(n_516) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND4xp75_ASAP7_75t_L g81 ( .A(n_82), .B(n_116), .C(n_134), .D(n_152), .Y(n_81) );
AND2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_108), .Y(n_82) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx3_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_96), .Y(n_86) );
AND2x4_ASAP7_75t_L g129 ( .A(n_87), .B(n_105), .Y(n_129) );
AND2x2_ASAP7_75t_L g147 ( .A(n_87), .B(n_120), .Y(n_147) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_91), .Y(n_87) );
INVx2_ASAP7_75t_L g107 ( .A(n_88), .Y(n_107) );
AND2x2_ASAP7_75t_L g124 ( .A(n_88), .B(n_92), .Y(n_124) );
BUFx2_ASAP7_75t_L g151 ( .A(n_88), .Y(n_151) );
INVx1_ASAP7_75t_L g90 ( .A(n_89), .Y(n_90) );
OAI22x1_ASAP7_75t_L g92 ( .A1(n_89), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_89), .Y(n_93) );
INVx2_ASAP7_75t_L g99 ( .A(n_89), .Y(n_99) );
INVx1_ASAP7_75t_L g102 ( .A(n_89), .Y(n_102) );
AND2x4_ASAP7_75t_L g106 ( .A(n_91), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g112 ( .A(n_92), .B(n_107), .Y(n_112) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_92), .Y(n_162) );
AND2x4_ASAP7_75t_L g111 ( .A(n_96), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g138 ( .A(n_96), .B(n_106), .Y(n_138) );
AND2x2_ASAP7_75t_L g155 ( .A(n_96), .B(n_124), .Y(n_155) );
AND2x4_ASAP7_75t_L g96 ( .A(n_97), .B(n_100), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x4_ASAP7_75t_L g105 ( .A(n_98), .B(n_100), .Y(n_105) );
AND2x2_ASAP7_75t_L g115 ( .A(n_98), .B(n_101), .Y(n_115) );
INVx1_ASAP7_75t_L g121 ( .A(n_98), .Y(n_121) );
INVxp67_ASAP7_75t_L g133 ( .A(n_100), .Y(n_133) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g120 ( .A(n_101), .B(n_121), .Y(n_120) );
BUFx3_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g158 ( .A(n_105), .B(n_112), .Y(n_158) );
AND2x4_ASAP7_75t_L g114 ( .A(n_106), .B(n_115), .Y(n_114) );
AND2x4_ASAP7_75t_L g141 ( .A(n_106), .B(n_120), .Y(n_141) );
INVx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx6_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x2_ASAP7_75t_L g119 ( .A(n_112), .B(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g150 ( .A(n_115), .B(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g161 ( .A(n_115), .B(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_127), .Y(n_116) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_121), .Y(n_126) );
BUFx6f_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x4_ASAP7_75t_L g132 ( .A(n_124), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx6_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_142), .Y(n_134) );
INVx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
INVx8_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx8_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx5_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx6_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx12f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OR2x2_ASAP7_75t_SL g164 ( .A(n_165), .B(n_167), .Y(n_164) );
AND2x2_ASAP7_75t_L g206 ( .A(n_165), .B(n_195), .Y(n_206) );
INVx1_ASAP7_75t_L g544 ( .A(n_165), .Y(n_544) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g190 ( .A(n_166), .B(n_191), .Y(n_190) );
AND3x1_ASAP7_75t_SL g537 ( .A(n_167), .B(n_538), .C(n_544), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_167), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2x1p5_ASAP7_75t_L g186 ( .A(n_168), .B(n_187), .Y(n_186) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND3x1_ASAP7_75t_L g171 ( .A(n_172), .B(n_401), .C(n_466), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_355), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_300), .B(n_328), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_263), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_211), .Y(n_175) );
AOI21xp33_ASAP7_75t_L g402 ( .A1(n_176), .A2(n_403), .B(n_414), .Y(n_402) );
AND2x2_ASAP7_75t_SL g437 ( .A(n_176), .B(n_344), .Y(n_437) );
AND2x2_ASAP7_75t_L g452 ( .A(n_176), .B(n_453), .Y(n_452) );
OR2x6_ASAP7_75t_L g462 ( .A(n_176), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g464 ( .A(n_176), .B(n_454), .Y(n_464) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g338 ( .A(n_177), .Y(n_338) );
AND2x2_ASAP7_75t_L g351 ( .A(n_177), .B(n_352), .Y(n_351) );
INVx4_ASAP7_75t_L g370 ( .A(n_177), .Y(n_370) );
AND2x2_ASAP7_75t_L g373 ( .A(n_177), .B(n_289), .Y(n_373) );
NOR2x1_ASAP7_75t_SL g376 ( .A(n_177), .B(n_304), .Y(n_376) );
AND2x4_ASAP7_75t_L g388 ( .A(n_177), .B(n_386), .Y(n_388) );
OR2x2_ASAP7_75t_L g398 ( .A(n_177), .B(n_270), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_177), .B(n_410), .Y(n_415) );
OR2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_183), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_179), .A2(n_224), .B1(n_230), .B2(n_231), .Y(n_223) );
INVx3_ASAP7_75t_L g231 ( .A(n_179), .Y(n_231) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_180), .B(n_234), .Y(n_233) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx4f_ASAP7_75t_L g215 ( .A(n_181), .Y(n_215) );
AND2x4_ASAP7_75t_L g209 ( .A(n_182), .B(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_SL g262 ( .A(n_182), .B(n_210), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_204), .B(n_209), .Y(n_183) );
INVxp67_ASAP7_75t_L g236 ( .A(n_185), .Y(n_236) );
AND2x4_ASAP7_75t_L g185 ( .A(n_186), .B(n_190), .Y(n_185) );
INVx1_ASAP7_75t_L g249 ( .A(n_187), .Y(n_249) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x6_ASAP7_75t_L g194 ( .A(n_188), .B(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x6_ASAP7_75t_L g313 ( .A(n_189), .B(n_198), .Y(n_313) );
AND2x6_ASAP7_75t_L g514 ( .A(n_190), .B(n_208), .Y(n_514) );
INVx2_ASAP7_75t_L g195 ( .A(n_191), .Y(n_195) );
AND2x4_ASAP7_75t_L g316 ( .A(n_191), .B(n_200), .Y(n_316) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .C(n_202), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_SL g217 ( .A1(n_194), .A2(n_202), .B(n_218), .C(n_219), .Y(n_217) );
INVxp67_ASAP7_75t_L g225 ( .A(n_194), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_194), .A2(n_202), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g275 ( .A1(n_194), .A2(n_202), .B(n_276), .C(n_277), .Y(n_275) );
INVx2_ASAP7_75t_L g299 ( .A(n_194), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_194), .A2(n_228), .B1(n_308), .B2(n_309), .Y(n_307) );
INVxp33_ASAP7_75t_L g248 ( .A(n_195), .Y(n_248) );
INVx1_ASAP7_75t_L g228 ( .A(n_197), .Y(n_228) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_200), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g245 ( .A(n_202), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_202), .A2(n_297), .B(n_298), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_202), .B(n_209), .Y(n_317) );
INVx5_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_203), .Y(n_229) );
INVx1_ASAP7_75t_L g238 ( .A(n_205), .Y(n_238) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
INVx1_ASAP7_75t_L g292 ( .A(n_206), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_207), .Y(n_293) );
BUFx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_211), .A2(n_344), .B1(n_439), .B2(n_440), .Y(n_438) );
INVx1_ASAP7_75t_SL g482 ( .A(n_211), .Y(n_482) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_239), .Y(n_211) );
INVx2_ASAP7_75t_L g413 ( .A(n_212), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_212), .B(n_359), .Y(n_485) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_221), .Y(n_212) );
BUFx3_ASAP7_75t_L g331 ( .A(n_213), .Y(n_331) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g324 ( .A(n_214), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_214), .B(n_241), .Y(n_346) );
AND2x4_ASAP7_75t_L g363 ( .A(n_214), .B(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_L g379 ( .A(n_214), .Y(n_379) );
INVx2_ASAP7_75t_L g436 ( .A(n_214), .Y(n_436) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_220), .Y(n_214) );
INVx2_ASAP7_75t_SL g242 ( .A(n_215), .Y(n_242) );
AND2x2_ASAP7_75t_L g354 ( .A(n_221), .B(n_320), .Y(n_354) );
NOR2xp67_ASAP7_75t_L g400 ( .A(n_221), .B(n_323), .Y(n_400) );
AND2x2_ASAP7_75t_L g419 ( .A(n_221), .B(n_323), .Y(n_419) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g281 ( .A(n_222), .Y(n_281) );
INVx1_ASAP7_75t_L g362 ( .A(n_222), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_222), .B(n_253), .Y(n_381) );
AND2x4_ASAP7_75t_L g435 ( .A(n_222), .B(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_232), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_231), .A2(n_254), .B(n_260), .Y(n_253) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_231), .A2(n_254), .B(n_260), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_236), .B1(n_237), .B2(n_238), .Y(n_232) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g394 ( .A(n_239), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_239), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_252), .Y(n_239) );
AND2x2_ASAP7_75t_L g378 ( .A(n_240), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g418 ( .A(n_240), .Y(n_418) );
AND2x2_ASAP7_75t_L g423 ( .A(n_240), .B(n_323), .Y(n_423) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_241), .B(n_253), .Y(n_283) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_251), .Y(n_241) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_242), .A2(n_243), .B(n_251), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_244), .B(n_250), .Y(n_243) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g359 ( .A(n_252), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_252), .B(n_331), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_252), .B(n_281), .Y(n_498) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_253), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_261), .Y(n_271) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI21xp33_ASAP7_75t_SL g263 ( .A1(n_264), .A2(n_279), .B(n_284), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_266), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g336 ( .A(n_267), .Y(n_336) );
AND2x2_ASAP7_75t_L g350 ( .A(n_267), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g384 ( .A(n_267), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g450 ( .A(n_267), .B(n_368), .Y(n_450) );
NOR3xp33_ASAP7_75t_L g496 ( .A(n_267), .B(n_497), .C(n_498), .Y(n_496) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_268), .Y(n_327) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g343 ( .A(n_270), .Y(n_343) );
AND2x2_ASAP7_75t_L g349 ( .A(n_270), .B(n_304), .Y(n_349) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_270), .Y(n_360) );
AND2x2_ASAP7_75t_L g405 ( .A(n_270), .B(n_303), .Y(n_405) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_270), .Y(n_428) );
INVx1_ASAP7_75t_L g445 ( .A(n_270), .Y(n_445) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B(n_278), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g487 ( .A(n_279), .Y(n_487) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_280), .B(n_358), .Y(n_459) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g321 ( .A(n_281), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI211x1_ASAP7_75t_L g355 ( .A1(n_285), .A2(n_356), .B(n_365), .C(n_382), .Y(n_355) );
INVx2_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_286), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g408 ( .A(n_286), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g344 ( .A(n_288), .B(n_303), .Y(n_344) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g302 ( .A(n_289), .B(n_303), .Y(n_302) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_289), .Y(n_369) );
INVx1_ASAP7_75t_L g386 ( .A(n_289), .Y(n_386) );
AND2x2_ASAP7_75t_L g454 ( .A(n_289), .B(n_304), .Y(n_454) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_295), .Y(n_289) );
NOR3xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .C(n_294), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_292), .A2(n_544), .B(n_555), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_293), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_318), .B(n_325), .Y(n_300) );
NOR2x1_ASAP7_75t_L g473 ( .A(n_301), .B(n_370), .Y(n_473) );
INVx2_ASAP7_75t_L g505 ( .A(n_301), .Y(n_505) );
INVx4_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g337 ( .A(n_302), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g410 ( .A(n_303), .Y(n_410) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g352 ( .A(n_304), .Y(n_352) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_310), .B(n_317), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B1(n_314), .B2(n_315), .Y(n_310) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
OR2x2_ASAP7_75t_L g412 ( .A(n_319), .B(n_413), .Y(n_412) );
NAND2x1_ASAP7_75t_SL g434 ( .A(n_319), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g334 ( .A(n_320), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g364 ( .A(n_320), .Y(n_364) );
INVx1_ASAP7_75t_L g488 ( .A(n_321), .Y(n_488) );
AND2x2_ASAP7_75t_L g353 ( .A(n_322), .B(n_354), .Y(n_353) );
NOR2x1_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g335 ( .A(n_323), .Y(n_335) );
INVxp33_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g392 ( .A(n_327), .B(n_385), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B(n_339), .C(n_347), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g416 ( .A(n_330), .B(n_417), .Y(n_416) );
NOR2xp67_ASAP7_75t_SL g421 ( .A(n_330), .B(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_331), .B(n_418), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_333), .B(n_337), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
AND2x2_ASAP7_75t_L g465 ( .A(n_334), .B(n_435), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g483 ( .A1(n_337), .A2(n_484), .B1(n_486), .B2(n_489), .C1(n_490), .C2(n_493), .Y(n_483) );
INVx1_ASAP7_75t_L g447 ( .A(n_338), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_345), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_343), .Y(n_374) );
AND2x4_ASAP7_75t_SL g409 ( .A(n_343), .B(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g463 ( .A(n_344), .Y(n_463) );
AND2x2_ASAP7_75t_L g508 ( .A(n_344), .B(n_360), .Y(n_508) );
AND2x2_ASAP7_75t_L g389 ( .A(n_345), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g502 ( .A(n_346), .B(n_381), .Y(n_502) );
OAI21xp33_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_350), .B(n_353), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_348), .A2(n_368), .B(n_409), .Y(n_469) );
AND2x2_ASAP7_75t_L g493 ( .A(n_349), .B(n_370), .Y(n_493) );
NOR2xp33_ASAP7_75t_SL g503 ( .A(n_349), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g441 ( .A(n_352), .Y(n_441) );
NOR2x1_ASAP7_75t_L g446 ( .A(n_352), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g476 ( .A(n_354), .Y(n_476) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_361), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x2_ASAP7_75t_L g479 ( .A(n_359), .B(n_363), .Y(n_479) );
BUFx2_ASAP7_75t_L g367 ( .A(n_360), .Y(n_367) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g390 ( .A(n_362), .Y(n_390) );
INVx2_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
AND2x2_ASAP7_75t_L g432 ( .A(n_362), .B(n_423), .Y(n_432) );
AND2x4_ASAP7_75t_L g399 ( .A(n_363), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g439 ( .A(n_363), .B(n_396), .Y(n_439) );
AND2x2_ASAP7_75t_L g490 ( .A(n_363), .B(n_491), .Y(n_490) );
AOI31xp33_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_371), .A3(n_375), .B(n_377), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
AND2x2_ASAP7_75t_L g387 ( .A(n_367), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_SL g368 ( .A(n_369), .B(n_370), .Y(n_368) );
AND2x4_ASAP7_75t_L g385 ( .A(n_370), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_373), .A2(n_425), .B1(n_456), .B2(n_459), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_373), .B(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g510 ( .A(n_373), .B(n_426), .Y(n_510) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g425 ( .A(n_376), .B(n_426), .Y(n_425) );
NAND2x1p5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
AND2x2_ASAP7_75t_L g448 ( .A(n_378), .B(n_419), .Y(n_448) );
INVx1_ASAP7_75t_L g458 ( .A(n_380), .Y(n_458) );
INVx2_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_391), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B(n_389), .Y(n_383) );
INVx1_ASAP7_75t_L g481 ( .A(n_384), .Y(n_481) );
AND2x2_ASAP7_75t_L g489 ( .A(n_385), .B(n_441), .Y(n_489) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_385), .Y(n_495) );
AND2x2_ASAP7_75t_L g440 ( .A(n_388), .B(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_393), .B1(n_397), .B2(n_399), .Y(n_391) );
NOR2xp33_ASAP7_75t_SL g393 ( .A(n_394), .B(n_395), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_394), .A2(n_413), .B1(n_507), .B2(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g406 ( .A(n_399), .Y(n_406) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_429), .Y(n_401) );
OAI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B(n_407), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
OAI21xp33_ASAP7_75t_L g407 ( .A1(n_405), .A2(n_408), .B(n_411), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_408), .A2(n_432), .B1(n_433), .B2(n_437), .Y(n_431) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_420), .B2(n_424), .Y(n_414) );
INVx1_ASAP7_75t_L g449 ( .A(n_417), .Y(n_449) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NOR2xp67_ASAP7_75t_L g429 ( .A(n_430), .B(n_442), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_438), .Y(n_430) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
NAND2xp33_ASAP7_75t_SL g484 ( .A(n_434), .B(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g457 ( .A(n_435), .Y(n_457) );
INVx3_ASAP7_75t_L g471 ( .A(n_439), .Y(n_471) );
INVxp67_ASAP7_75t_L g500 ( .A(n_440), .Y(n_500) );
NAND4xp25_ASAP7_75t_L g442 ( .A(n_443), .B(n_451), .C(n_455), .D(n_460), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_448), .B1(n_449), .B2(n_450), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
AND2x2_ASAP7_75t_L g453 ( .A(n_445), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g501 ( .A(n_449), .Y(n_501) );
NAND2xp33_ASAP7_75t_SL g456 ( .A(n_457), .B(n_458), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_464), .B(n_465), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND3x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_483), .C(n_494), .Y(n_466) );
AOI221x1_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B1(n_472), .B2(n_474), .C(n_480), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp33_ASAP7_75t_SL g474 ( .A(n_475), .B(n_478), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
NAND2xp33_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI211xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_499), .C(n_506), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_499) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_535), .B1(n_545), .B2(n_546), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_518), .Y(n_552) );
XOR2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_526), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B1(n_531), .B2(n_534), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_531), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
INVxp67_ASAP7_75t_L g550 ( .A(n_538), .Y(n_550) );
CKINVDCx8_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g548 ( .A(n_544), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_554), .Y(n_553) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
endmodule