module fake_jpeg_10728_n_169 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_9),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_0),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_2),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_3),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_81),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_3),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_64),
.Y(n_96)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

BUFx24_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_71),
.B1(n_53),
.B2(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_61),
.B1(n_7),
.B2(n_8),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_71),
.B1(n_67),
.B2(n_63),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_88),
.B1(n_97),
.B2(n_70),
.Y(n_104)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_73),
.B1(n_55),
.B2(n_68),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g91 ( 
.A(n_80),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_80),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_96),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_53),
.B1(n_70),
.B2(n_67),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_100),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_80),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_102),
.B(n_105),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_106),
.B1(n_109),
.B2(n_114),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_69),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_50),
.B1(n_59),
.B2(n_73),
.Y(n_106)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_73),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_117),
.B(n_10),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_60),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_110),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_72),
.B1(n_66),
.B2(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_4),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_4),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_5),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_61),
.B1(n_7),
.B2(n_9),
.Y(n_116)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_10),
.B(n_11),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_6),
.Y(n_117)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_27),
.A3(n_48),
.B1(n_46),
.B2(n_44),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_35),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_136),
.Y(n_148)
);

OAI22x1_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_94),
.B1(n_22),
.B2(n_26),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_124),
.B1(n_126),
.B2(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_6),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_128),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_114),
.B1(n_116),
.B2(n_101),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_121),
.B(n_137),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_100),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_134),
.C(n_127),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_13),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_135),
.Y(n_146)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_31),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_14),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_133),
.B(n_130),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_14),
.B(n_15),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_141),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_138),
.A2(n_36),
.B(n_16),
.C(n_17),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_15),
.B1(n_19),
.B2(n_28),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_145),
.B1(n_147),
.B2(n_151),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_49),
.B1(n_123),
.B2(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_149),
.B(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_134),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_157),
.A2(n_148),
.B(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_153),
.B1(n_152),
.B2(n_147),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_161),
.B1(n_156),
.B2(n_155),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_141),
.B1(n_145),
.B2(n_151),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_163),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_156),
.B(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_142),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_142),
.Y(n_169)
);


endmodule