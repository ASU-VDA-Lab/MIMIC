module fake_aes_6721_n_27 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_27);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_27;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_2), .Y(n_10) );
NAND2xp5_ASAP7_75t_SL g11 ( .A(n_7), .B(n_0), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_5), .Y(n_13) );
AOI21x1_ASAP7_75t_L g14 ( .A1(n_2), .A2(n_1), .B(n_8), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_5), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_3), .B(n_9), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_10), .B(n_0), .Y(n_17) );
A2O1A1Ixp33_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_11), .B(n_15), .C(n_13), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AOI222xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_11), .B1(n_18), .B2(n_12), .C1(n_19), .C2(n_14), .Y(n_22) );
AOI211xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_19), .B(n_16), .C(n_14), .Y(n_23) );
BUFx12f_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
BUFx2_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_24), .B(n_19), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_25), .B1(n_4), .B2(n_6), .Y(n_27) );
endmodule