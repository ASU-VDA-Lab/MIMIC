module real_aes_2512_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_753, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_754, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_753;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_754;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_404;
wire n_288;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_717;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g153 ( .A(n_0), .B(n_127), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_1), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_2), .B(n_111), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_3), .B(n_129), .Y(n_446) );
INVx1_ASAP7_75t_L g118 ( .A(n_4), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_5), .B(n_111), .Y(n_180) );
NAND2xp33_ASAP7_75t_SL g223 ( .A(n_6), .B(n_117), .Y(n_223) );
INVx1_ASAP7_75t_L g215 ( .A(n_7), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g748 ( .A(n_8), .Y(n_748) );
AND2x2_ASAP7_75t_L g178 ( .A(n_9), .B(n_135), .Y(n_178) );
AND2x2_ASAP7_75t_L g448 ( .A(n_10), .B(n_131), .Y(n_448) );
AND2x2_ASAP7_75t_L g458 ( .A(n_11), .B(n_221), .Y(n_458) );
INVx2_ASAP7_75t_L g133 ( .A(n_12), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_13), .B(n_129), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_14), .Y(n_418) );
AOI221x1_ASAP7_75t_L g218 ( .A1(n_15), .A2(n_120), .B1(n_219), .B2(n_221), .C(n_222), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g110 ( .A(n_16), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_17), .B(n_111), .Y(n_503) );
INVx1_ASAP7_75t_L g421 ( .A(n_18), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_19), .A2(n_88), .B1(n_111), .B2(n_164), .Y(n_462) );
AOI221xp5_ASAP7_75t_SL g142 ( .A1(n_20), .A2(n_36), .B1(n_111), .B2(n_120), .C(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_21), .A2(n_120), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_22), .B(n_127), .Y(n_183) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_23), .A2(n_87), .B(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g136 ( .A(n_23), .B(n_87), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_24), .B(n_129), .Y(n_128) );
INVxp67_ASAP7_75t_L g217 ( .A(n_25), .Y(n_217) );
AND2x2_ASAP7_75t_L g204 ( .A(n_26), .B(n_141), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_27), .A2(n_120), .B(n_152), .Y(n_151) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_28), .A2(n_221), .B(n_494), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_29), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_30), .B(n_129), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_31), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_31), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_32), .A2(n_120), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_33), .B(n_129), .Y(n_518) );
AND2x2_ASAP7_75t_L g117 ( .A(n_34), .B(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g121 ( .A(n_34), .B(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g172 ( .A(n_34), .Y(n_172) );
OR2x6_ASAP7_75t_L g419 ( .A(n_35), .B(n_420), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g746 ( .A(n_35), .B(n_747), .C(n_749), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_37), .B(n_111), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_38), .A2(n_79), .B1(n_120), .B2(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_39), .B(n_129), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_40), .B(n_111), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_41), .B(n_127), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_42), .A2(n_120), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g156 ( .A(n_43), .B(n_141), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_44), .B(n_127), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_45), .B(n_141), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_46), .B(n_111), .Y(n_495) );
INVx1_ASAP7_75t_L g114 ( .A(n_47), .Y(n_114) );
INVx1_ASAP7_75t_L g124 ( .A(n_47), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_48), .B(n_129), .Y(n_456) );
AND2x2_ASAP7_75t_L g485 ( .A(n_49), .B(n_141), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_50), .B(n_111), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_51), .B(n_127), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_52), .B(n_127), .Y(n_517) );
AND2x2_ASAP7_75t_L g195 ( .A(n_53), .B(n_141), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_54), .B(n_111), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_55), .B(n_129), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_56), .B(n_111), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_57), .A2(n_120), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_SL g134 ( .A(n_58), .B(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_59), .B(n_127), .Y(n_192) );
AND2x2_ASAP7_75t_L g509 ( .A(n_60), .B(n_135), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_61), .A2(n_120), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_62), .B(n_129), .Y(n_184) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_63), .B(n_131), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_64), .B(n_127), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_65), .B(n_127), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_66), .A2(n_90), .B1(n_120), .B2(n_170), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_67), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_68), .B(n_129), .Y(n_506) );
INVx1_ASAP7_75t_L g116 ( .A(n_69), .Y(n_116) );
INVx1_ASAP7_75t_L g122 ( .A(n_69), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_70), .B(n_127), .Y(n_445) );
OAI222xp33_ASAP7_75t_L g101 ( .A1(n_71), .A2(n_102), .B1(n_710), .B2(n_711), .C1(n_717), .C2(n_720), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_71), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_72), .A2(n_120), .B(n_489), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g435 ( .A1(n_73), .A2(n_120), .B(n_436), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_74), .A2(n_120), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g520 ( .A(n_75), .B(n_135), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_76), .B(n_141), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_77), .A2(n_81), .B1(n_111), .B2(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_78), .B(n_111), .Y(n_193) );
INVx1_ASAP7_75t_L g422 ( .A(n_80), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_82), .B(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_83), .B(n_127), .Y(n_145) );
AND2x2_ASAP7_75t_L g439 ( .A(n_84), .B(n_131), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_85), .Y(n_731) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_86), .A2(n_120), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_89), .B(n_129), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_91), .A2(n_120), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_92), .B(n_129), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_93), .B(n_111), .Y(n_155) );
INVxp67_ASAP7_75t_L g220 ( .A(n_94), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_95), .B(n_129), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_96), .A2(n_120), .B(n_125), .Y(n_119) );
BUFx2_ASAP7_75t_L g508 ( .A(n_97), .Y(n_508) );
BUFx2_ASAP7_75t_L g725 ( .A(n_98), .Y(n_725) );
BUFx2_ASAP7_75t_SL g734 ( .A(n_98), .Y(n_734) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_742), .B(n_750), .Y(n_99) );
OA21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_721), .B(n_732), .Y(n_100) );
AOI22xp5_ASAP7_75t_SL g102 ( .A1(n_103), .A2(n_417), .B1(n_423), .B2(n_707), .Y(n_102) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_103), .A2(n_423), .B1(n_713), .B2(n_716), .Y(n_712) );
INVx3_ASAP7_75t_SL g738 ( .A(n_103), .Y(n_738) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_103), .Y(n_739) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_309), .Y(n_103) );
NOR3xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_237), .C(n_287), .Y(n_104) );
OAI211xp5_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_157), .B(n_205), .C(n_226), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_137), .Y(n_106) );
AND2x2_ASAP7_75t_L g236 ( .A(n_107), .B(n_138), .Y(n_236) );
INVx1_ASAP7_75t_L g367 ( .A(n_107), .Y(n_367) );
NOR2x1p5_ASAP7_75t_L g399 ( .A(n_107), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g210 ( .A(n_108), .B(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g258 ( .A(n_108), .Y(n_258) );
OR2x2_ASAP7_75t_L g262 ( .A(n_108), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_108), .B(n_140), .Y(n_274) );
OR2x2_ASAP7_75t_L g296 ( .A(n_108), .B(n_140), .Y(n_296) );
AND2x4_ASAP7_75t_L g302 ( .A(n_108), .B(n_266), .Y(n_302) );
OR2x2_ASAP7_75t_L g319 ( .A(n_108), .B(n_212), .Y(n_319) );
INVx1_ASAP7_75t_L g354 ( .A(n_108), .Y(n_354) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_108), .Y(n_376) );
OR2x2_ASAP7_75t_L g390 ( .A(n_108), .B(n_323), .Y(n_390) );
AND2x4_ASAP7_75t_SL g394 ( .A(n_108), .B(n_212), .Y(n_394) );
OR2x6_ASAP7_75t_L g108 ( .A(n_109), .B(n_134), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_119), .B(n_131), .Y(n_109) );
AND2x4_ASAP7_75t_L g111 ( .A(n_112), .B(n_117), .Y(n_111) );
INVx1_ASAP7_75t_L g224 ( .A(n_112), .Y(n_224) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
AND2x6_ASAP7_75t_L g127 ( .A(n_113), .B(n_122), .Y(n_127) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g129 ( .A(n_115), .B(n_124), .Y(n_129) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx5_ASAP7_75t_L g130 ( .A(n_117), .Y(n_130) );
AND2x2_ASAP7_75t_L g123 ( .A(n_118), .B(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_118), .Y(n_167) );
AND2x6_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
BUFx3_ASAP7_75t_L g168 ( .A(n_121), .Y(n_168) );
INVx2_ASAP7_75t_L g174 ( .A(n_122), .Y(n_174) );
AND2x4_ASAP7_75t_L g170 ( .A(n_123), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_128), .B(n_130), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_127), .B(n_508), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_130), .A2(n_144), .B(n_145), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_130), .A2(n_153), .B(n_154), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_130), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_130), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_130), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_130), .A2(n_437), .B(n_438), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_130), .A2(n_445), .B(n_446), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_130), .A2(n_455), .B(n_456), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_130), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_130), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_130), .A2(n_506), .B(n_507), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_130), .A2(n_517), .B(n_518), .Y(n_516) );
INVx2_ASAP7_75t_SL g161 ( .A(n_131), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_131), .A2(n_503), .B(n_504), .Y(n_502) );
BUFx4f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx3_ASAP7_75t_L g149 ( .A(n_132), .Y(n_149) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_133), .B(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g185 ( .A(n_133), .B(n_136), .Y(n_185) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g346 ( .A(n_138), .B(n_302), .Y(n_346) );
AND2x2_ASAP7_75t_L g393 ( .A(n_138), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_147), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
AND2x2_ASAP7_75t_L g256 ( .A(n_140), .B(n_147), .Y(n_256) );
INVx2_ASAP7_75t_L g263 ( .A(n_140), .Y(n_263) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_140), .Y(n_384) );
BUFx3_ASAP7_75t_L g400 ( .A(n_140), .Y(n_400) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_146), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_141), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_141), .A2(n_434), .B(n_435), .Y(n_433) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_141), .A2(n_462), .B(n_463), .Y(n_461) );
INVx2_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_147), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g323 ( .A(n_147), .B(n_263), .Y(n_323) );
INVx1_ASAP7_75t_L g341 ( .A(n_147), .Y(n_341) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_147), .Y(n_357) );
INVx1_ASAP7_75t_L g379 ( .A(n_147), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_147), .B(n_258), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_147), .B(n_212), .Y(n_416) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21x1_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_156), .Y(n_148) );
INVx4_ASAP7_75t_L g221 ( .A(n_149), .Y(n_221) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_149), .A2(n_452), .B(n_458), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
INVx1_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_176), .Y(n_158) );
AND2x4_ASAP7_75t_L g230 ( .A(n_159), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g241 ( .A(n_159), .Y(n_241) );
AND2x2_ASAP7_75t_L g246 ( .A(n_159), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g281 ( .A(n_159), .B(n_186), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_159), .B(n_187), .Y(n_291) );
OR2x2_ASAP7_75t_L g371 ( .A(n_159), .B(n_286), .Y(n_371) );
OAI322xp33_ASAP7_75t_L g401 ( .A1(n_159), .A2(n_314), .A3(n_353), .B1(n_386), .B2(n_402), .C1(n_403), .C2(n_404), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_159), .B(n_384), .Y(n_402) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g235 ( .A(n_160), .Y(n_235) );
AOI21x1_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_175), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_169), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_164), .A2(n_170), .B1(n_214), .B2(n_216), .Y(n_213) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_168), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
NOR2x1p5_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_176), .A2(n_348), .B1(n_352), .B2(n_355), .Y(n_347) );
AOI211xp5_ASAP7_75t_L g407 ( .A1(n_176), .A2(n_408), .B(n_409), .C(n_412), .Y(n_407) );
AND2x4_ASAP7_75t_SL g176 ( .A(n_177), .B(n_186), .Y(n_176) );
AND2x4_ASAP7_75t_L g229 ( .A(n_177), .B(n_197), .Y(n_229) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_177), .Y(n_233) );
INVx5_ASAP7_75t_L g245 ( .A(n_177), .Y(n_245) );
INVx2_ASAP7_75t_L g254 ( .A(n_177), .Y(n_254) );
AND2x2_ASAP7_75t_L g277 ( .A(n_177), .B(n_187), .Y(n_277) );
AND2x2_ASAP7_75t_L g306 ( .A(n_177), .B(n_196), .Y(n_306) );
OR2x2_ASAP7_75t_L g315 ( .A(n_177), .B(n_235), .Y(n_315) );
OR2x2_ASAP7_75t_L g330 ( .A(n_177), .B(n_244), .Y(n_330) );
OR2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_185), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_185), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_185), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_185), .B(n_220), .Y(n_219) );
NOR3xp33_ASAP7_75t_L g222 ( .A(n_185), .B(n_223), .C(n_224), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_185), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_185), .A2(n_495), .B(n_496), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_186), .B(n_206), .Y(n_205) );
INVx3_ASAP7_75t_SL g314 ( .A(n_186), .Y(n_314) );
AND2x2_ASAP7_75t_L g337 ( .A(n_186), .B(n_245), .Y(n_337) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_196), .Y(n_186) );
INVx2_ASAP7_75t_L g231 ( .A(n_187), .Y(n_231) );
AND2x2_ASAP7_75t_L g234 ( .A(n_187), .B(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g248 ( .A(n_187), .B(n_197), .Y(n_248) );
INVx1_ASAP7_75t_L g252 ( .A(n_187), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_187), .B(n_197), .Y(n_286) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_187), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_187), .B(n_245), .Y(n_361) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_194), .B(n_195), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_193), .Y(n_188) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_194), .A2(n_198), .B(n_204), .Y(n_197) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_194), .A2(n_198), .B(n_204), .Y(n_244) );
AOI21x1_ASAP7_75t_L g441 ( .A1(n_194), .A2(n_442), .B(n_448), .Y(n_441) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
AND2x2_ASAP7_75t_L g351 ( .A(n_197), .B(n_235), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_199), .B(n_203), .Y(n_198) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_210), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_207), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OR2x6_ASAP7_75t_SL g415 ( .A(n_208), .B(n_416), .Y(n_415) );
INVxp67_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_209), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_209), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g363 ( .A(n_209), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_210), .A2(n_272), .B1(n_275), .B2(n_282), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_211), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g307 ( .A(n_211), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_211), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_211), .B(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_225), .Y(n_211) );
AND2x2_ASAP7_75t_L g257 ( .A(n_212), .B(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g266 ( .A(n_212), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_212), .A2(n_273), .B1(n_325), .B2(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g332 ( .A(n_212), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_212), .B(n_326), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_212), .B(n_256), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_212), .B(n_263), .Y(n_405) );
AND2x4_ASAP7_75t_L g212 ( .A(n_213), .B(n_218), .Y(n_212) );
INVx3_ASAP7_75t_L g513 ( .A(n_221), .Y(n_513) );
OAI21xp33_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_232), .B(n_236), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_230), .Y(n_227) );
NAND4xp25_ASAP7_75t_SL g275 ( .A(n_228), .B(n_276), .C(n_278), .D(n_280), .Y(n_275) );
INVx2_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_229), .B(n_336), .Y(n_365) );
AND2x2_ASAP7_75t_L g392 ( .A(n_229), .B(n_230), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_229), .B(n_252), .Y(n_403) );
INVx1_ASAP7_75t_L g268 ( .A(n_230), .Y(n_268) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_230), .A2(n_293), .B1(n_304), .B2(n_307), .Y(n_303) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_230), .B(n_243), .C(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_230), .B(n_245), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_230), .B(n_253), .Y(n_396) );
AND2x2_ASAP7_75t_L g328 ( .A(n_231), .B(n_235), .Y(n_328) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_231), .Y(n_389) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g284 ( .A(n_233), .Y(n_284) );
INVx1_ASAP7_75t_L g374 ( .A(n_234), .Y(n_374) );
AND2x2_ASAP7_75t_L g381 ( .A(n_234), .B(n_245), .Y(n_381) );
BUFx2_ASAP7_75t_L g336 ( .A(n_235), .Y(n_336) );
NAND3xp33_ASAP7_75t_SL g237 ( .A(n_238), .B(n_259), .C(n_271), .Y(n_237) );
OAI31xp33_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_246), .A3(n_249), .B(n_255), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_239), .A2(n_293), .B1(n_297), .B2(n_298), .Y(n_292) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
OR2x2_ASAP7_75t_L g278 ( .A(n_241), .B(n_279), .Y(n_278) );
NOR2x1_ASAP7_75t_L g304 ( .A(n_241), .B(n_305), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g373 ( .A1(n_242), .A2(n_344), .B(n_374), .C(n_375), .Y(n_373) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_243), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_244), .B(n_252), .Y(n_279) );
AND2x2_ASAP7_75t_L g297 ( .A(n_244), .B(n_277), .Y(n_297) );
AND2x2_ASAP7_75t_L g414 ( .A(n_247), .B(n_336), .Y(n_414) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g270 ( .A(n_248), .B(n_254), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_253), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g345 ( .A(n_253), .B(n_328), .Y(n_345) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_254), .B(n_328), .Y(n_334) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g326 ( .A(n_256), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_257), .B(n_357), .Y(n_356) );
AOI32xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_267), .A3(n_268), .B1(n_269), .B2(n_753), .Y(n_259) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_260), .A2(n_345), .B1(n_381), .B2(n_382), .C(n_385), .Y(n_380) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_263), .Y(n_308) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g273 ( .A(n_265), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g378 ( .A(n_266), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_267), .B(n_289), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g311 ( .A1(n_269), .A2(n_312), .B1(n_316), .B2(n_320), .C(n_324), .Y(n_311) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OAI211xp5_ASAP7_75t_L g287 ( .A1(n_274), .A2(n_288), .B(n_292), .C(n_303), .Y(n_287) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OAI322xp33_ASAP7_75t_L g385 ( .A1(n_280), .A2(n_290), .A3(n_339), .B1(n_386), .B2(n_387), .C1(n_388), .C2(n_390), .Y(n_385) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI21xp33_ASAP7_75t_L g412 ( .A1(n_283), .A2(n_413), .B(n_415), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_289), .A2(n_370), .B(n_372), .C(n_373), .Y(n_369) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g411 ( .A(n_296), .B(n_377), .Y(n_411) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_302), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g386 ( .A(n_302), .Y(n_386) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI31xp33_ASAP7_75t_L g342 ( .A1(n_306), .A2(n_343), .A3(n_345), .B(n_346), .Y(n_342) );
NOR2x1_ASAP7_75t_L g309 ( .A(n_310), .B(n_368), .Y(n_309) );
NAND5xp2_ASAP7_75t_L g310 ( .A(n_311), .B(n_331), .C(n_342), .D(n_347), .E(n_358), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AOI21xp33_ASAP7_75t_L g409 ( .A1(n_314), .A2(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g382 ( .A(n_318), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B(n_335), .C(n_338), .Y(n_331) );
INVxp33_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
OR2x2_ASAP7_75t_L g360 ( .A(n_336), .B(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_339), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g410 ( .A(n_351), .Y(n_410) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_362), .B(n_364), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI21xp33_ASAP7_75t_L g364 ( .A1(n_360), .A2(n_365), .B(n_366), .Y(n_364) );
NAND4xp25_ASAP7_75t_L g368 ( .A(n_369), .B(n_380), .C(n_391), .D(n_407), .Y(n_368) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_378), .B(n_399), .Y(n_398) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g408 ( .A(n_390), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_395), .B2(n_397), .C(n_401), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_417), .Y(n_715) );
AND2x6_ASAP7_75t_SL g417 ( .A(n_418), .B(n_419), .Y(n_417) );
OR2x6_ASAP7_75t_SL g708 ( .A(n_418), .B(n_709), .Y(n_708) );
OR2x2_ASAP7_75t_L g719 ( .A(n_418), .B(n_419), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_418), .B(n_709), .Y(n_730) );
CKINVDCx16_ASAP7_75t_R g749 ( .A(n_418), .Y(n_749) );
CKINVDCx5p33_ASAP7_75t_R g709 ( .A(n_419), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_421), .B(n_422), .Y(n_745) );
AND2x4_ASAP7_75t_L g423 ( .A(n_424), .B(n_620), .Y(n_423) );
NOR4xp75_ASAP7_75t_L g424 ( .A(n_425), .B(n_543), .C(n_568), .D(n_595), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_480), .B(n_521), .Y(n_425) );
NOR4xp25_ASAP7_75t_L g426 ( .A(n_427), .B(n_464), .C(n_471), .D(n_475), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_449), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_440), .Y(n_430) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_431), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_431), .B(n_468), .Y(n_614) );
AND2x2_ASAP7_75t_L g639 ( .A(n_431), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g664 ( .A(n_431), .B(n_459), .Y(n_664) );
AND2x2_ASAP7_75t_L g705 ( .A(n_431), .B(n_473), .Y(n_705) );
INVx4_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_SL g477 ( .A(n_432), .B(n_470), .Y(n_477) );
AND2x2_ASAP7_75t_L g479 ( .A(n_432), .B(n_451), .Y(n_479) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_432), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g540 ( .A(n_432), .Y(n_540) );
AND2x2_ASAP7_75t_L g546 ( .A(n_432), .B(n_473), .Y(n_546) );
BUFx2_ASAP7_75t_L g559 ( .A(n_432), .Y(n_559) );
AND2x4_ASAP7_75t_L g590 ( .A(n_432), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g637 ( .A(n_432), .B(n_638), .Y(n_637) );
OR2x6_ASAP7_75t_L g432 ( .A(n_433), .B(n_439), .Y(n_432) );
INVx1_ASAP7_75t_L g631 ( .A(n_440), .Y(n_631) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g470 ( .A(n_441), .Y(n_470) );
AND2x2_ASAP7_75t_L g473 ( .A(n_441), .B(n_451), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_447), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_449), .B(n_649), .Y(n_702) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g539 ( .A(n_450), .B(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_459), .Y(n_450) );
INVx2_ASAP7_75t_L g469 ( .A(n_451), .Y(n_469) );
INVx2_ASAP7_75t_L g530 ( .A(n_451), .Y(n_530) );
AND2x2_ASAP7_75t_L g640 ( .A(n_451), .B(n_470), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .Y(n_452) );
INVx2_ASAP7_75t_L g528 ( .A(n_459), .Y(n_528) );
BUFx3_ASAP7_75t_L g545 ( .A(n_459), .Y(n_545) );
AND2x2_ASAP7_75t_L g572 ( .A(n_459), .B(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
AND2x4_ASAP7_75t_L g466 ( .A(n_460), .B(n_461), .Y(n_466) );
NOR2x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
INVx2_ASAP7_75t_L g474 ( .A(n_465), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_465), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g643 ( .A(n_465), .B(n_583), .Y(n_643) );
AND2x2_ASAP7_75t_L g667 ( .A(n_465), .B(n_477), .Y(n_667) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g563 ( .A(n_466), .B(n_469), .Y(n_563) );
AND2x2_ASAP7_75t_L g645 ( .A(n_466), .B(n_638), .Y(n_645) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g688 ( .A(n_468), .Y(n_688) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g573 ( .A(n_469), .Y(n_573) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_470), .Y(n_577) );
INVx2_ASAP7_75t_L g585 ( .A(n_470), .Y(n_585) );
INVx1_ASAP7_75t_L g591 ( .A(n_470), .Y(n_591) );
AOI222xp33_ASAP7_75t_SL g521 ( .A1(n_471), .A2(n_522), .B1(n_526), .B2(n_531), .C1(n_538), .C2(n_541), .Y(n_521) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g598 ( .A(n_473), .Y(n_598) );
BUFx2_ASAP7_75t_L g627 ( .A(n_473), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g621 ( .A1(n_474), .A2(n_622), .B(n_626), .C(n_634), .Y(n_621) );
OR2x2_ASAP7_75t_L g692 ( .A(n_474), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g700 ( .A(n_474), .B(n_605), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_477), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g675 ( .A(n_477), .B(n_563), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_477), .B(n_655), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_478), .B(n_545), .Y(n_683) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g605 ( .A(n_479), .B(n_577), .Y(n_605) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_500), .Y(n_481) );
INVx1_ASAP7_75t_L g699 ( .A(n_482), .Y(n_699) );
NOR2xp67_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
AND2x2_ASAP7_75t_L g542 ( .A(n_483), .B(n_501), .Y(n_542) );
INVx1_ASAP7_75t_L g619 ( .A(n_483), .Y(n_619) );
OR2x2_ASAP7_75t_L g678 ( .A(n_483), .B(n_501), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_483), .B(n_550), .Y(n_684) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g525 ( .A(n_484), .Y(n_525) );
OR2x2_ASAP7_75t_L g557 ( .A(n_484), .B(n_511), .Y(n_557) );
AND2x2_ASAP7_75t_L g566 ( .A(n_484), .B(n_493), .Y(n_566) );
NAND2x1_ASAP7_75t_L g594 ( .A(n_484), .B(n_501), .Y(n_594) );
AND2x2_ASAP7_75t_L g641 ( .A(n_484), .B(n_536), .Y(n_641) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g524 ( .A(n_493), .Y(n_524) );
INVx1_ASAP7_75t_L g534 ( .A(n_493), .Y(n_534) );
AND2x2_ASAP7_75t_L g550 ( .A(n_493), .B(n_537), .Y(n_550) );
INVx2_ASAP7_75t_L g555 ( .A(n_493), .Y(n_555) );
OR2x2_ASAP7_75t_L g651 ( .A(n_493), .B(n_501), .Y(n_651) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
NOR2x1_ASAP7_75t_SL g536 ( .A(n_501), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g554 ( .A(n_501), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g567 ( .A(n_501), .B(n_511), .Y(n_567) );
BUFx2_ASAP7_75t_L g586 ( .A(n_501), .Y(n_586) );
INVx2_ASAP7_75t_SL g613 ( .A(n_501), .Y(n_613) );
OR2x6_ASAP7_75t_L g501 ( .A(n_502), .B(n_509), .Y(n_501) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g523 ( .A(n_511), .B(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g669 ( .A(n_511), .B(n_611), .Y(n_669) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_520), .Y(n_512) );
AO21x1_ASAP7_75t_SL g537 ( .A1(n_513), .A2(n_514), .B(n_520), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_519), .Y(n_514) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_522), .A2(n_546), .B(n_686), .C(n_690), .Y(n_685) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_523), .B(n_601), .Y(n_636) );
BUFx2_ASAP7_75t_L g600 ( .A(n_524), .Y(n_600) );
OR2x2_ASAP7_75t_L g548 ( .A(n_525), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g633 ( .A(n_525), .B(n_567), .Y(n_633) );
AND2x2_ASAP7_75t_L g654 ( .A(n_525), .B(n_610), .Y(n_654) );
INVx2_ASAP7_75t_L g661 ( .A(n_525), .Y(n_661) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_526), .A2(n_667), .B(n_668), .Y(n_666) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
AND2x2_ASAP7_75t_L g608 ( .A(n_527), .B(n_590), .Y(n_608) );
OR2x2_ASAP7_75t_L g687 ( .A(n_527), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_528), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_530), .Y(n_561) );
AND2x2_ASAP7_75t_L g638 ( .A(n_530), .B(n_585), .Y(n_638) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g623 ( .A(n_533), .B(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_SL g632 ( .A(n_533), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_533), .B(n_542), .Y(n_665) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g541 ( .A(n_534), .B(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g660 ( .A(n_535), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g610 ( .A(n_536), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g580 ( .A(n_537), .B(n_555), .Y(n_580) );
OAI31xp33_ASAP7_75t_L g587 ( .A1(n_538), .A2(n_588), .A3(n_590), .B(n_592), .Y(n_587) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_540), .B(n_563), .Y(n_589) );
AO21x1_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_547), .B(n_551), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
OR2x2_ASAP7_75t_L g599 ( .A(n_545), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g704 ( .A(n_545), .Y(n_704) );
INVx2_ASAP7_75t_SL g689 ( .A(n_546), .Y(n_689) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g593 ( .A(n_549), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g677 ( .A(n_549), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_550), .B(n_613), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_558), .B1(n_562), .B2(n_564), .Y(n_551) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_552), .A2(n_671), .B(n_672), .Y(n_670) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
INVx1_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g625 ( .A(n_557), .B(n_586), .Y(n_625) );
OR2x2_ASAP7_75t_L g650 ( .A(n_557), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_559), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_559), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g649 ( .A(n_559), .Y(n_649) );
INVx2_ASAP7_75t_L g578 ( .A(n_560), .Y(n_578) );
INVx1_ASAP7_75t_L g658 ( .A(n_561), .Y(n_658) );
AND2x2_ASAP7_75t_L g581 ( .A(n_563), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g655 ( .A(n_563), .Y(n_655) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_569), .B(n_587), .Y(n_568) );
OAI321xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_574), .A3(n_579), .B1(n_580), .B2(n_581), .C(n_586), .Y(n_569) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_570), .A2(n_601), .A3(n_696), .B1(n_698), .B2(n_700), .C1(n_701), .C2(n_706), .Y(n_695) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx2_ASAP7_75t_L g648 ( .A(n_573), .Y(n_648) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_575), .B(n_655), .Y(n_672) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g680 ( .A(n_578), .Y(n_680) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp33_ASAP7_75t_SL g612 ( .A(n_580), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI21xp33_ASAP7_75t_SL g679 ( .A1(n_583), .A2(n_589), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx3_ASAP7_75t_L g601 ( .A(n_594), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_615), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_601), .B1(n_602), .B2(n_603), .C(n_606), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_598), .Y(n_617) );
AND2x2_ASAP7_75t_L g602 ( .A(n_600), .B(n_601), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OAI22xp33_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_609), .B1(n_612), .B2(n_614), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g618 ( .A(n_610), .B(n_619), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_613), .A2(n_702), .B(n_703), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR3xp33_ASAP7_75t_SL g620 ( .A(n_621), .B(n_652), .C(n_673), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_625), .A2(n_660), .B1(n_687), .B2(n_689), .Y(n_686) );
OAI21xp33_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_628), .B(n_632), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_627), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_633), .A2(n_675), .B1(n_676), .B2(n_679), .C(n_681), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .B1(n_639), .B2(n_641), .C(n_642), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g671 ( .A(n_637), .Y(n_671) );
INVx1_ASAP7_75t_L g693 ( .A(n_638), .Y(n_693) );
INVx1_ASAP7_75t_SL g691 ( .A(n_639), .Y(n_691) );
AOI31xp33_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .A3(n_646), .B(n_650), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_643), .A2(n_653), .B1(n_655), .B2(n_656), .C(n_754), .Y(n_652) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B(n_662), .C(n_670), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g668 ( .A(n_661), .B(n_669), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_665), .B(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g697 ( .A(n_669), .Y(n_697) );
BUFx2_ASAP7_75t_SL g706 ( .A(n_669), .Y(n_706) );
NAND3xp33_ASAP7_75t_SL g673 ( .A(n_674), .B(n_685), .C(n_695), .Y(n_673) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B(n_684), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B(n_694), .Y(n_690) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_SL g716 ( .A(n_707), .Y(n_716) );
CKINVDCx11_ASAP7_75t_R g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx4_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx3_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx3_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_726), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_727), .A2(n_736), .B(n_740), .Y(n_735) );
NOR2xp33_ASAP7_75t_SL g727 ( .A(n_728), .B(n_731), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
BUFx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
BUFx2_ASAP7_75t_L g741 ( .A(n_730), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
CKINVDCx5p33_ASAP7_75t_R g733 ( .A(n_734), .Y(n_733) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_744), .B(n_751), .Y(n_750) );
AND2x4_ASAP7_75t_SL g744 ( .A(n_745), .B(n_746), .Y(n_744) );
endmodule