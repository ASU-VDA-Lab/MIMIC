module fake_jpeg_5594_n_174 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_174);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_3),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_41),
.Y(n_58)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_27),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_53),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_19),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_31),
.B1(n_28),
.B2(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_57),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_15),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_26),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_23),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_71),
.B1(n_63),
.B2(n_49),
.Y(n_92)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_61),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_17),
.B1(n_34),
.B2(n_30),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_66),
.B1(n_55),
.B2(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_17),
.B1(n_15),
.B2(n_30),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_18),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_54),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_63),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_45),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_91),
.C(n_51),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_69),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_89),
.B1(n_71),
.B2(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_49),
.B(n_58),
.C(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_92),
.A2(n_93),
.B1(n_69),
.B2(n_42),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_51),
.B1(n_58),
.B2(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_93),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_89),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_42),
.B(n_70),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_107),
.B(n_86),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_83),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_70),
.B(n_56),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_101),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_56),
.C(n_43),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_111),
.C(n_112),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_43),
.C(n_64),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_64),
.C(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_97),
.B(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_120),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_119),
.B1(n_125),
.B2(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_76),
.B(n_18),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_126),
.C(n_105),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_94),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_61),
.C(n_76),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_18),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_98),
.B1(n_101),
.B2(n_99),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_3),
.B(n_4),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_136),
.C(n_113),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_108),
.C(n_103),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_1),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_25),
.B(n_22),
.C(n_16),
.D(n_23),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_16),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_149),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_116),
.B1(n_120),
.B2(n_16),
.Y(n_141)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_147),
.C(n_13),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_0),
.B(n_1),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_145),
.B(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_3),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_10),
.C(n_12),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_11),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_7),
.C(n_8),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_154),
.B(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_139),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_134),
.B(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_140),
.C(n_149),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_4),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_162),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_157),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_132),
.C(n_143),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_153),
.B(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_148),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_167),
.B(n_160),
.C(n_4),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_166),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_6),
.B(n_170),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_168),
.C(n_6),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);


endmodule