module fake_jpeg_3839_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_35),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_17),
.C(n_29),
.Y(n_52)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_44),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_54),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_16),
.B1(n_19),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_47),
.B1(n_27),
.B2(n_24),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g83 ( 
.A(n_50),
.Y(n_83)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_63),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_22),
.B1(n_25),
.B2(n_16),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_29),
.B1(n_27),
.B2(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_16),
.B1(n_19),
.B2(n_22),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_17),
.B1(n_27),
.B2(n_29),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_38),
.Y(n_102)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_82),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_60),
.Y(n_80)
);

NOR2x1_ASAP7_75t_R g101 ( 
.A(n_80),
.B(n_34),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_39),
.Y(n_95)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_44),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_102),
.B(n_28),
.Y(n_126)
);

AOI32xp33_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_51),
.A3(n_50),
.B1(n_56),
.B2(n_34),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_72),
.Y(n_112)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_108),
.Y(n_130)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_49),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_103),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_75),
.B(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_28),
.B1(n_21),
.B2(n_18),
.Y(n_127)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_107),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_35),
.C(n_49),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_78),
.C(n_65),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_17),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_20),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_111),
.C(n_114),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_113),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_65),
.C(n_80),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_127),
.B1(n_107),
.B2(n_89),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_84),
.C(n_69),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_122),
.B(n_98),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_82),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_69),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_125),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_76),
.B1(n_79),
.B2(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_128),
.B1(n_95),
.B2(n_87),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_74),
.B(n_73),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_18),
.B1(n_55),
.B2(n_39),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_108),
.B(n_87),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_64),
.C(n_34),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_30),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_21),
.B1(n_55),
.B2(n_54),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_131),
.B(n_133),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_97),
.B1(n_105),
.B2(n_103),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_139),
.B(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_97),
.B1(n_88),
.B2(n_86),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_135),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_136),
.B(n_138),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_144),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_89),
.B1(n_104),
.B2(n_90),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_31),
.B1(n_26),
.B2(n_64),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_31),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_54),
.B1(n_33),
.B2(n_59),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_116),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_59),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_157),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_125),
.C(n_119),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_158),
.C(n_30),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_139),
.A2(n_112),
.B(n_115),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_30),
.B(n_1),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_126),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_127),
.C(n_33),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_130),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_26),
.Y(n_179)
);

NAND4xp25_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_57),
.C(n_33),
.D(n_26),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_161),
.Y(n_172)
);

OA21x2_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_33),
.B(n_31),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_163),
.B(n_148),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_31),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_177),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_144),
.B(n_151),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_181),
.B(n_157),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_179),
.C(n_182),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_146),
.A3(n_136),
.B1(n_140),
.B2(n_131),
.C1(n_145),
.C2(n_141),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_147),
.B1(n_57),
.B2(n_26),
.Y(n_178)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_184),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_152),
.A2(n_30),
.B(n_26),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_170),
.A2(n_159),
.B1(n_167),
.B2(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_194),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_155),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_190),
.C(n_191),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_156),
.C(n_162),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_158),
.C(n_160),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_183),
.B(n_181),
.C(n_175),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_173),
.C(n_174),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_187),
.C(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_154),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_200),
.A2(n_203),
.B(n_205),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_172),
.B1(n_173),
.B2(n_169),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_161),
.A3(n_168),
.B1(n_187),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_188),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_190),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_206),
.B(n_210),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_212),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_191),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_203),
.Y(n_213)
);

OAI321xp33_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_6),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_218),
.C(n_8),
.Y(n_221)
);

A2O1A1O1Ixp25_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_0),
.B(n_1),
.C(n_2),
.D(n_4),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_215),
.B(n_9),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_6),
.B(n_7),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_221),
.B(n_222),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_13),
.C1(n_216),
.C2(n_213),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_9),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_224),
.Y(n_226)
);


endmodule