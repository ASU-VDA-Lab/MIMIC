module fake_jpeg_14192_n_553 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_553);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_553;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_SL g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_11),
.B(n_7),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_22),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_57),
.B(n_91),
.Y(n_126)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_64),
.B(n_106),
.Y(n_127)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g164 ( 
.A(n_68),
.B(n_50),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_69),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_70),
.Y(n_111)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_74),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_85),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_99),
.Y(n_109)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_13),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_94),
.Y(n_163)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_97),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_40),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

CKINVDCx6p67_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_19),
.B(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_53),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_113),
.B(n_133),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_38),
.B1(n_51),
.B2(n_25),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_115),
.A2(n_118),
.B1(n_128),
.B2(n_105),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_77),
.A2(n_49),
.B1(n_31),
.B2(n_17),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_66),
.A2(n_26),
.B1(n_39),
.B2(n_38),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_122),
.A2(n_129),
.B1(n_146),
.B2(n_169),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_80),
.A2(n_17),
.B1(n_31),
.B2(n_49),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_66),
.A2(n_26),
.B1(n_39),
.B2(n_51),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_26),
.B1(n_49),
.B2(n_31),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_130),
.A2(n_147),
.B1(n_46),
.B2(n_35),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_45),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_131),
.B(n_141),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_68),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_135),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_70),
.B(n_45),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_48),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_46),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_70),
.A2(n_39),
.B1(n_17),
.B2(n_25),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_81),
.A2(n_20),
.B1(n_42),
.B2(n_37),
.Y(n_147)
);

INVx6_ASAP7_75t_SL g151 ( 
.A(n_84),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_151),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_103),
.A2(n_18),
.B(n_32),
.Y(n_158)
);

OAI32xp33_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_3),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_164),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_85),
.B(n_41),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_40),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_86),
.A2(n_18),
.B1(n_48),
.B2(n_47),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_173),
.Y(n_176)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_178),
.Y(n_251)
);

AND2x2_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_59),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_179),
.B(n_219),
.C(n_119),
.Y(n_252)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_180),
.Y(n_253)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_139),
.A2(n_37),
.B1(n_42),
.B2(n_30),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_139),
.A2(n_30),
.B1(n_50),
.B2(n_47),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_183),
.Y(n_264)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_186),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_189),
.B(n_199),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_227),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_115),
.A2(n_92),
.B1(n_98),
.B2(n_96),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_120),
.A2(n_93),
.B1(n_88),
.B2(n_87),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_194),
.Y(n_272)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_196),
.Y(n_274)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_197),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_146),
.A2(n_74),
.B1(n_62),
.B2(n_55),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_198),
.A2(n_201),
.B1(n_203),
.B2(n_212),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_126),
.B(n_41),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_200),
.B(n_208),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_129),
.A2(n_35),
.B1(n_32),
.B2(n_4),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_205),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_163),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_206)
);

AOI32xp33_ASAP7_75t_L g281 ( 
.A1(n_206),
.A2(n_207),
.A3(n_160),
.B1(n_202),
.B2(n_199),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_127),
.B(n_132),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_156),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_224),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_152),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_122),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_213),
.B(n_221),
.Y(n_282)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_214),
.Y(n_292)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_136),
.Y(n_215)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_117),
.Y(n_216)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_216),
.Y(n_279)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_121),
.B(n_8),
.Y(n_219)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_123),
.B(n_9),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_222),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_172),
.Y(n_223)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_156),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_124),
.B(n_12),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_225),
.B(n_221),
.Y(n_286)
);

AO22x1_ASAP7_75t_SL g226 ( 
.A1(n_137),
.A2(n_12),
.B1(n_13),
.B2(n_142),
.Y(n_226)
);

AO22x1_ASAP7_75t_SL g269 ( 
.A1(n_226),
.A2(n_229),
.B1(n_145),
.B2(n_170),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_112),
.A2(n_13),
.B1(n_162),
.B2(n_165),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_140),
.A2(n_13),
.B1(n_149),
.B2(n_138),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_152),
.A2(n_111),
.B1(n_161),
.B2(n_167),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_231),
.Y(n_288)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_155),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_234),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_125),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_108),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_108),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_235),
.B(n_236),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_125),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_110),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_238),
.Y(n_285)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_138),
.A2(n_149),
.B1(n_162),
.B2(n_112),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_239),
.A2(n_160),
.B1(n_190),
.B2(n_240),
.Y(n_277)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_140),
.Y(n_240)
);

NAND2x1_ASAP7_75t_SL g295 ( 
.A(n_240),
.B(n_235),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_111),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_243),
.B(n_256),
.C(n_293),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_200),
.B(n_119),
.CI(n_167),
.CON(n_244),
.SN(n_244)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_244),
.B(n_246),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_188),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_210),
.B(n_172),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_249),
.B(n_273),
.Y(n_348)
);

XNOR2x1_ASAP7_75t_L g317 ( 
.A(n_252),
.B(n_204),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_205),
.B(n_110),
.C(n_145),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_176),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_265),
.B(n_267),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_176),
.Y(n_267)
);

NOR2x1p5_ASAP7_75t_L g268 ( 
.A(n_210),
.B(n_119),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_290),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_269),
.A2(n_281),
.B1(n_252),
.B2(n_264),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_217),
.B(n_170),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_271),
.B(n_289),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_179),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_276),
.B(n_291),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_277),
.A2(n_247),
.B1(n_253),
.B2(n_294),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_286),
.B(n_298),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_187),
.B(n_225),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_219),
.B(n_207),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_179),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_219),
.B(n_184),
.C(n_180),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_238),
.B(n_195),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_250),
.A2(n_201),
.B1(n_198),
.B2(n_229),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_299),
.A2(n_318),
.B1(n_343),
.B2(n_275),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_282),
.A2(n_206),
.B(n_213),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_300),
.A2(n_333),
.B(n_275),
.Y(n_359)
);

OAI22x1_ASAP7_75t_SL g301 ( 
.A1(n_250),
.A2(n_229),
.B1(n_226),
.B2(n_216),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_301),
.B(n_315),
.Y(n_358)
);

O2A1O1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_264),
.A2(n_229),
.B(n_226),
.C(n_233),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_302),
.B(n_305),
.Y(n_366)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_304),
.Y(n_350)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_266),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_312),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_255),
.A2(n_277),
.B1(n_257),
.B2(n_283),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_284),
.Y(n_312)
);

NAND2x1_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_177),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g379 ( 
.A1(n_313),
.A2(n_348),
.B(n_309),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_243),
.B(n_254),
.C(n_293),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_314),
.B(n_338),
.C(n_344),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_181),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_255),
.A2(n_214),
.B(n_178),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_316),
.A2(n_335),
.B(n_309),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_322),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_290),
.A2(n_218),
.B1(n_220),
.B2(n_209),
.Y(n_318)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_258),
.Y(n_320)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_321),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_254),
.B(n_237),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_257),
.A2(n_223),
.B1(n_237),
.B2(n_288),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_330),
.Y(n_363)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_242),
.Y(n_326)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_326),
.Y(n_371)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_297),
.Y(n_327)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_328),
.Y(n_378)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_329),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_244),
.B(n_241),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_339),
.Y(n_361)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_297),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_332),
.B(n_334),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_249),
.A2(n_244),
.B1(n_269),
.B2(n_256),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_262),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_249),
.A2(n_269),
.B(n_278),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_336),
.A2(n_258),
.B1(n_294),
.B2(n_270),
.Y(n_349)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_251),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_337),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_259),
.B(n_263),
.Y(n_338)
);

NOR2x1p5_ASAP7_75t_SL g339 ( 
.A(n_295),
.B(n_274),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_262),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_341),
.Y(n_360)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_261),
.A2(n_260),
.B1(n_287),
.B2(n_272),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_285),
.C(n_253),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_247),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_345),
.Y(n_353)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_261),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_367),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_315),
.B(n_270),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_369),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_324),
.B(n_273),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_313),
.B(n_292),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_374),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_338),
.B(n_279),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_325),
.A2(n_279),
.B(n_330),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_379),
.A2(n_381),
.B(n_320),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_331),
.B(n_313),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_389),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_335),
.B(n_322),
.Y(n_382)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_314),
.B(n_317),
.C(n_303),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_344),
.C(n_334),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_316),
.A2(n_311),
.B(n_333),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_385),
.A2(n_327),
.B(n_332),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_299),
.A2(n_318),
.B1(n_302),
.B2(n_301),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_386),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_311),
.A2(n_300),
.B1(n_347),
.B2(n_303),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_388),
.A2(n_348),
.B1(n_340),
.B2(n_339),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_346),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_391),
.B(n_374),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_357),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_407),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_348),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_399),
.C(n_401),
.Y(n_436)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_350),
.Y(n_396)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_396),
.Y(n_428)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_352),
.Y(n_398)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_398),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_304),
.C(n_306),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_358),
.A2(n_337),
.B1(n_329),
.B2(n_328),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_403),
.A2(n_418),
.B1(n_422),
.B2(n_355),
.Y(n_425)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_352),
.Y(n_408)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_408),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_321),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_412),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_419),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_375),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_413),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_366),
.A2(n_343),
.B1(n_358),
.B2(n_388),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_414),
.A2(n_421),
.B1(n_423),
.B2(n_353),
.Y(n_449)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_357),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_417),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_385),
.A2(n_359),
.B1(n_382),
.B2(n_351),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_375),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_368),
.Y(n_420)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_420),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_366),
.A2(n_370),
.B1(n_377),
.B2(n_364),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_366),
.A2(n_361),
.B1(n_380),
.B2(n_363),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_354),
.A2(n_379),
.B1(n_361),
.B2(n_365),
.Y(n_423)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_356),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_431),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_393),
.B(n_365),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_427),
.B(n_432),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g431 ( 
.A(n_404),
.Y(n_431)
);

XNOR2x1_ASAP7_75t_SL g433 ( 
.A(n_422),
.B(n_363),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_433),
.B(n_445),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_362),
.C(n_360),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_437),
.B(n_442),
.C(n_447),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_395),
.Y(n_438)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_438),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_405),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_439),
.B(n_451),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_406),
.A2(n_353),
.B1(n_349),
.B2(n_362),
.Y(n_441)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_375),
.C(n_387),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_443),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_391),
.B(n_383),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_394),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_390),
.Y(n_448)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_449),
.A2(n_409),
.B1(n_418),
.B2(n_400),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_394),
.B(n_383),
.C(n_372),
.Y(n_451)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_454),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_414),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_476),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_454),
.Y(n_460)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_460),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_420),
.Y(n_461)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_407),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_463),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_464),
.A2(n_467),
.B1(n_421),
.B2(n_435),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_402),
.C(n_416),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_427),
.C(n_432),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_446),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_466),
.B(n_437),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_449),
.A2(n_409),
.B1(n_400),
.B2(n_453),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_405),
.Y(n_470)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_470),
.Y(n_495)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_428),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_473),
.Y(n_483)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_430),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_434),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_475),
.Y(n_489)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_440),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_416),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_444),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_452),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_429),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_480),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_482),
.A2(n_496),
.B(n_479),
.Y(n_501)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g485 ( 
.A(n_460),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_485),
.A2(n_488),
.B1(n_490),
.B2(n_493),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_457),
.A2(n_441),
.B1(n_425),
.B2(n_426),
.Y(n_490)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_491),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_442),
.C(n_445),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_492),
.B(n_497),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_457),
.A2(n_390),
.B1(n_435),
.B2(n_411),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_419),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_458),
.B(n_398),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_470),
.B(n_413),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_467),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_433),
.C(n_419),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_456),
.C(n_477),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_501),
.A2(n_486),
.B(n_455),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_487),
.B(n_456),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_502),
.B(n_508),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_465),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_503),
.B(n_507),
.Y(n_520)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_504),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_506),
.B(n_511),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_492),
.B(n_464),
.C(n_477),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_499),
.B(n_476),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_469),
.Y(n_511)
);

OAI22x1_ASAP7_75t_L g512 ( 
.A1(n_481),
.A2(n_472),
.B1(n_463),
.B2(n_462),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_512),
.A2(n_403),
.B1(n_408),
.B2(n_376),
.Y(n_527)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_495),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_491),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_482),
.B(n_472),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_495),
.C(n_481),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_516),
.B(n_524),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_517),
.B(n_521),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_500),
.A2(n_486),
.B1(n_494),
.B2(n_461),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_518),
.B(n_513),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_494),
.C(n_480),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_480),
.C(n_496),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_512),
.C(n_507),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_489),
.Y(n_523)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_523),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_510),
.A2(n_483),
.B1(n_397),
.B2(n_396),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_526),
.A2(n_372),
.B1(n_376),
.B2(n_378),
.Y(n_535)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_527),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_530),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_525),
.A2(n_505),
.B1(n_506),
.B2(n_415),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_532),
.B(n_536),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_535),
.B(n_526),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_527),
.A2(n_503),
.B1(n_378),
.B2(n_502),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_538),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_531),
.B(n_528),
.C(n_520),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_540),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_533),
.B(n_516),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_541),
.A2(n_542),
.B(n_530),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_537),
.B(n_522),
.Y(n_542)
);

O2A1O1Ixp33_ASAP7_75t_SL g547 ( 
.A1(n_544),
.A2(n_543),
.B(n_539),
.C(n_537),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_547),
.B(n_548),
.Y(n_549)
);

OAI21xp33_ASAP7_75t_L g548 ( 
.A1(n_546),
.A2(n_534),
.B(n_529),
.Y(n_548)
);

OAI211xp5_ASAP7_75t_L g550 ( 
.A1(n_549),
.A2(n_545),
.B(n_535),
.C(n_521),
.Y(n_550)
);

OAI21x1_ASAP7_75t_SL g551 ( 
.A1(n_550),
.A2(n_519),
.B(n_373),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_519),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_373),
.Y(n_553)
);


endmodule