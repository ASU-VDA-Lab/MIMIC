module fake_jpeg_19518_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_4),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_11),
.B(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_0),
.B(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_32),
.Y(n_52)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_22),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_15),
.B1(n_26),
.B2(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_43),
.B1(n_49),
.B2(n_60),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_15),
.B1(n_26),
.B2(n_19),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_32),
.C(n_33),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_48),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_25),
.C(n_20),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_49)
);

AO22x1_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_22),
.B1(n_23),
.B2(n_13),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_28),
.B(n_29),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_10),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_13),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_17),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_34),
.A2(n_23),
.B1(n_20),
.B2(n_17),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_71),
.B(n_76),
.Y(n_85)
);

AOI32xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_44),
.A3(n_28),
.B1(n_48),
.B2(n_46),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_73),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_57),
.B(n_50),
.C(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_33),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_78),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_35),
.B(n_29),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_52),
.B(n_51),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_72),
.B1(n_74),
.B2(n_64),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_52),
.C(n_47),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_89),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_67),
.B(n_76),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_52),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_5),
.C(n_6),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_71),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_64),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_103),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_100),
.B(n_101),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_12),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_98),
.A2(n_99),
.B(n_11),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_9),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_70),
.B1(n_71),
.B2(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_107),
.B1(n_92),
.B2(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_81),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_111),
.C(n_113),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_82),
.C(n_85),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_91),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_85),
.C(n_88),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_71),
.B1(n_86),
.B2(n_78),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_104),
.C(n_96),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_119),
.C(n_122),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_104),
.C(n_103),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_121),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_108),
.C(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_126),
.Y(n_130)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_100),
.B1(n_108),
.B2(n_86),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_79),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_131),
.B(n_123),
.Y(n_132)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_8),
.B(n_77),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_7),
.A3(n_8),
.B1(n_58),
.B2(n_66),
.C1(n_77),
.C2(n_123),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.C(n_130),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_128),
.B(n_129),
.Y(n_135)
);

BUFx24_ASAP7_75t_SL g136 ( 
.A(n_135),
.Y(n_136)
);


endmodule