module fake_ariane_1147_n_1131 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_262, n_20, n_174, n_275, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_122, n_268, n_257, n_266, n_198, n_148, n_232, n_164, n_52, n_277, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_276, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1131);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_262;
input n_20;
input n_174;
input n_275;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_277;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_276;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1131;

wire n_295;
wire n_556;
wire n_356;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_515;
wire n_445;
wire n_807;
wire n_765;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_926;
wire n_813;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1068;
wire n_1052;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_557;
wire n_405;
wire n_1107;
wire n_989;
wire n_645;
wire n_858;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_600;
wire n_433;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_821;
wire n_770;
wire n_839;
wire n_928;
wire n_1099;
wire n_507;
wire n_465;
wire n_486;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_604;
wire n_439;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_1080;
wire n_576;
wire n_843;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_654;
wire n_455;
wire n_429;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_612;
wire n_333;
wire n_449;
wire n_388;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_658;
wire n_630;
wire n_570;
wire n_1055;
wire n_543;
wire n_362;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_939;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_571;
wire n_680;
wire n_414;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_1108;
wire n_355;
wire n_609;
wire n_444;
wire n_851;
wire n_278;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_664;
wire n_629;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_626;
wire n_430;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_697;
wire n_622;
wire n_437;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_1027;
wire n_615;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_108),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_82),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_136),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_174),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_144),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_13),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_143),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_215),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_45),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_102),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_129),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_128),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_35),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_169),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_92),
.B(n_277),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_25),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_27),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_161),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_53),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_29),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_197),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_85),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_262),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_109),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_135),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_31),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_140),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_198),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_255),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_97),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_110),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_167),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_17),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_176),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_162),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_100),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_242),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_192),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_84),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_63),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_166),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_12),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_260),
.B(n_137),
.Y(n_322)
);

BUFx10_ASAP7_75t_L g323 ( 
.A(n_22),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_257),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_42),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_51),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_4),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_23),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_175),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_152),
.B(n_25),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_32),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_43),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_210),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_274),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_105),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_12),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_74),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_91),
.Y(n_338)
);

INVx4_ASAP7_75t_R g339 ( 
.A(n_68),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_39),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_111),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_79),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_44),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_267),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_142),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_122),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_229),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_119),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_15),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_203),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_173),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_146),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_171),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_40),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_187),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_177),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_107),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_150),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_132),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_88),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_251),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_259),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_275),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_185),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_241),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_49),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_148),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_249),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_205),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_253),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_248),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_223),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_52),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_121),
.Y(n_374)
);

BUFx2_ASAP7_75t_SL g375 ( 
.A(n_264),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_254),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_28),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_96),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_120),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_258),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_151),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_59),
.Y(n_382)
);

INVx4_ASAP7_75t_R g383 ( 
.A(n_200),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_95),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_41),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_89),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_80),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_245),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_33),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_207),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_70),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_190),
.Y(n_392)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_2),
.B(n_58),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_117),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_99),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_47),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_219),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_38),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_228),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_32),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_23),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_62),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_73),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_60),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_67),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_116),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_178),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_123),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_226),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_103),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_17),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_34),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_46),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_240),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_125),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_147),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_16),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_21),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_118),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_61),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_75),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_26),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_165),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_57),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_256),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_208),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_16),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_6),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_182),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_261),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_37),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_236),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_188),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_48),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_170),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_71),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_101),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_217),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_83),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_195),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_232),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_276),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_272),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_141),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_154),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_263),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_196),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_26),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g449 ( 
.A(n_193),
.B(n_124),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_186),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_55),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_72),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_145),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_246),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_153),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_421),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_347),
.B(n_0),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_421),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_286),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_279),
.A2(n_0),
.B(n_1),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_336),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_347),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_284),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_328),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_302),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_398),
.B(n_5),
.Y(n_466)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_297),
.A2(n_163),
.B(n_270),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_328),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_303),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_398),
.B(n_7),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_407),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_421),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_393),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_323),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_328),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_317),
.B(n_10),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_338),
.A2(n_168),
.B(n_269),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_323),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_295),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_328),
.Y(n_480)
);

INVx6_ASAP7_75t_L g481 ( 
.A(n_411),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_331),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_335),
.B(n_11),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_294),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_428),
.B(n_11),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_411),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_299),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_337),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_421),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_331),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_321),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_327),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_352),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_377),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_352),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_331),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_282),
.B(n_13),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_401),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_308),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_331),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_287),
.B(n_14),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_340),
.B(n_18),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_417),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_349),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_296),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_289),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_349),
.Y(n_508)
);

OA21x2_ASAP7_75t_L g509 ( 
.A1(n_290),
.A2(n_19),
.B(n_20),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_418),
.B(n_422),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_291),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_349),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_427),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_379),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

INVx6_ASAP7_75t_L g516 ( 
.A(n_447),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_363),
.B(n_19),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_305),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_395),
.B(n_20),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_300),
.B(n_21),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_352),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_301),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_402),
.B(n_424),
.Y(n_523)
);

BUFx8_ASAP7_75t_SL g524 ( 
.A(n_313),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_332),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_443),
.B(n_24),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_446),
.B(n_28),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_306),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_307),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_359),
.A2(n_184),
.B(n_268),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_309),
.B(n_29),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_312),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_448),
.B(n_30),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_310),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_333),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_389),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_389),
.Y(n_537)
);

BUFx8_ASAP7_75t_L g538 ( 
.A(n_368),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_389),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_314),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_318),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_454),
.B(n_50),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_372),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_320),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_384),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_324),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_413),
.B(n_54),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_341),
.B(n_56),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_350),
.B(n_273),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_342),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_351),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_357),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_360),
.B(n_266),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_361),
.B(n_364),
.Y(n_554)
);

INVx5_ASAP7_75t_L g555 ( 
.A(n_339),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_370),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_374),
.B(n_69),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_378),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_493),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_493),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_479),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_518),
.B(n_292),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_503),
.A2(n_440),
.B1(n_453),
.B2(n_452),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_491),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_523),
.B(n_367),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_494),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_497),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_518),
.B(n_292),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_473),
.A2(n_344),
.B1(n_438),
.B2(n_450),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_517),
.B(n_345),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_482),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_482),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_456),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_504),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_456),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_508),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_519),
.B(n_345),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_488),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_L g581 ( 
.A(n_457),
.B(n_278),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_547),
.B(n_371),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_513),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_464),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_468),
.Y(n_585)
);

AND3x2_ASAP7_75t_L g586 ( 
.A(n_470),
.B(n_483),
.C(n_476),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_475),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_507),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_480),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_459),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_456),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_490),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_528),
.B(n_367),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_507),
.Y(n_594)
);

BUFx4f_ASAP7_75t_L g595 ( 
.A(n_543),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_R g596 ( 
.A(n_459),
.B(n_471),
.Y(n_596)
);

INVx8_ASAP7_75t_L g597 ( 
.A(n_555),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_471),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_488),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_466),
.B(n_397),
.C(n_371),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_547),
.B(n_462),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_532),
.B(n_280),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_496),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_511),
.Y(n_604)
);

AO21x2_ASAP7_75t_L g605 ( 
.A1(n_548),
.A2(n_330),
.B(n_380),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_511),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_481),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_516),
.B(n_281),
.Y(n_608)
);

AND2x6_ASAP7_75t_L g609 ( 
.A(n_476),
.B(n_381),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_501),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_522),
.Y(n_611)
);

NAND3xp33_ASAP7_75t_L g612 ( 
.A(n_466),
.B(n_406),
.C(n_397),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_514),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_495),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_483),
.B(n_386),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_544),
.B(n_391),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_516),
.A2(n_355),
.B1(n_387),
.B2(n_420),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_495),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_495),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_515),
.B(n_557),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_495),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_522),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_536),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_551),
.B(n_392),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_554),
.B(n_406),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_541),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_543),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_536),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_536),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_536),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_541),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_556),
.B(n_394),
.Y(n_632)
);

AOI21x1_ASAP7_75t_L g633 ( 
.A1(n_548),
.A2(n_403),
.B(n_396),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_546),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_516),
.B(n_348),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_558),
.B(n_405),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_481),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_546),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_543),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_527),
.B(n_285),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_L g641 ( 
.A(n_526),
.B(n_288),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_543),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_542),
.B(n_408),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_637),
.B(n_538),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_627),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_627),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_590),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_643),
.B(n_555),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_643),
.B(n_555),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_609),
.B(n_555),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_609),
.B(n_552),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_561),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_637),
.B(n_538),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_564),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_609),
.B(n_552),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_600),
.A2(n_485),
.B1(n_527),
.B2(n_533),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_566),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_567),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_600),
.A2(n_485),
.B1(n_529),
.B2(n_534),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_570),
.A2(n_473),
.B1(n_469),
.B2(n_465),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_568),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_562),
.B(n_545),
.Y(n_662)
);

A2O1A1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_582),
.A2(n_553),
.B(n_498),
.C(n_520),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_573),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_573),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_562),
.B(n_569),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_559),
.B(n_481),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_572),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_559),
.B(n_484),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_569),
.B(n_560),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_602),
.B(n_506),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_597),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_560),
.B(n_545),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_609),
.B(n_545),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_584),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_585),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_565),
.B(n_545),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_575),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_598),
.B(n_532),
.Y(n_679)
);

O2A1O1Ixp5_ASAP7_75t_L g680 ( 
.A1(n_633),
.A2(n_502),
.B(n_498),
.C(n_520),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_615),
.B(n_540),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_596),
.Y(n_682)
);

INVx8_ASAP7_75t_L g683 ( 
.A(n_597),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_565),
.B(n_608),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_587),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_615),
.B(n_549),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_615),
.B(n_549),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_583),
.Y(n_688)
);

A2O1A1Ixp33_ASAP7_75t_L g689 ( 
.A1(n_582),
.A2(n_553),
.B(n_531),
.C(n_502),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_635),
.B(n_486),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_625),
.B(n_521),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_599),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_640),
.B(n_474),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_613),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_589),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_592),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_625),
.B(n_521),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_620),
.B(n_615),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_620),
.B(n_521),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_603),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_612),
.A2(n_477),
.B(n_467),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_615),
.B(n_521),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_610),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_588),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_577),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_599),
.B(n_537),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_578),
.Y(n_707)
);

OR2x6_ASAP7_75t_L g708 ( 
.A(n_570),
.B(n_525),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_640),
.B(n_531),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_601),
.B(n_537),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_594),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_604),
.Y(n_712)
);

NOR3xp33_ASAP7_75t_L g713 ( 
.A(n_612),
.B(n_525),
.C(n_461),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_639),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_606),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_601),
.B(n_537),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_607),
.B(n_550),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_611),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_622),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_596),
.B(n_535),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_571),
.A2(n_500),
.B1(n_463),
.B2(n_499),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_626),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_571),
.B(n_579),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_631),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_605),
.B(n_409),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_634),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_579),
.A2(n_510),
.B1(n_460),
.B2(n_509),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_586),
.B(n_510),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_581),
.A2(n_463),
.B1(n_487),
.B2(n_499),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_SL g730 ( 
.A(n_586),
.B(n_358),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_652),
.Y(n_731)
);

O2A1O1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_666),
.A2(n_593),
.B(n_624),
.C(n_636),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_670),
.B(n_593),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_654),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_691),
.A2(n_641),
.B(n_597),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_709),
.B(n_605),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_728),
.B(n_617),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_671),
.B(n_563),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_657),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_SL g740 ( 
.A1(n_663),
.A2(n_616),
.B(n_624),
.C(n_636),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_697),
.A2(n_632),
.B(n_616),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_723),
.A2(n_632),
.B(n_530),
.C(n_638),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_686),
.A2(n_595),
.B(n_642),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_705),
.Y(n_744)
);

O2A1O1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_689),
.A2(n_487),
.B(n_512),
.C(n_505),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_698),
.A2(n_375),
.B1(n_444),
.B2(n_416),
.Y(n_746)
);

OAI21xp5_ASAP7_75t_L g747 ( 
.A1(n_701),
.A2(n_509),
.B(n_460),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_707),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_728),
.B(n_580),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_669),
.B(n_365),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_692),
.B(n_595),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_664),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_647),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_684),
.B(n_478),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_692),
.B(n_667),
.Y(n_755)
);

CKINVDCx10_ASAP7_75t_R g756 ( 
.A(n_708),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_658),
.A2(n_433),
.B(n_451),
.C(n_426),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_679),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_730),
.B(n_693),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_648),
.B(n_298),
.Y(n_760)
);

NAND2x1p5_ASAP7_75t_L g761 ( 
.A(n_672),
.B(n_430),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_661),
.A2(n_434),
.B(n_441),
.C(n_431),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_682),
.Y(n_763)
);

AOI22x1_ASAP7_75t_L g764 ( 
.A1(n_701),
.A2(n_455),
.B1(n_435),
.B2(n_432),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_686),
.A2(n_293),
.B(n_283),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_680),
.A2(n_283),
.B(n_293),
.C(n_322),
.Y(n_766)
);

AO21x1_ASAP7_75t_L g767 ( 
.A1(n_725),
.A2(n_618),
.B(n_614),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_687),
.A2(n_621),
.B(n_619),
.Y(n_768)
);

AO21x2_ASAP7_75t_L g769 ( 
.A1(n_725),
.A2(n_449),
.B(n_630),
.Y(n_769)
);

AO22x1_ASAP7_75t_L g770 ( 
.A1(n_713),
.A2(n_524),
.B1(n_478),
.B2(n_304),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_687),
.A2(n_629),
.B(n_628),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_SL g772 ( 
.A(n_730),
.B(n_524),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_727),
.A2(n_623),
.B(n_315),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_708),
.A2(n_404),
.B1(n_316),
.B2(n_319),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_656),
.A2(n_410),
.B1(n_325),
.B2(n_326),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_729),
.B(n_537),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_690),
.B(n_311),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_681),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_672),
.B(n_329),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_694),
.Y(n_780)
);

OAI21x1_ASAP7_75t_L g781 ( 
.A1(n_702),
.A2(n_383),
.B(n_576),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_660),
.B(n_415),
.C(n_343),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_648),
.B(n_334),
.Y(n_783)
);

O2A1O1Ixp5_ASAP7_75t_L g784 ( 
.A1(n_651),
.A2(n_655),
.B(n_688),
.C(n_678),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_662),
.A2(n_419),
.B(n_353),
.Y(n_785)
);

BUFx4f_ASAP7_75t_L g786 ( 
.A(n_683),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_649),
.B(n_346),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_704),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_649),
.A2(n_425),
.B(n_356),
.Y(n_789)
);

OAI21xp33_ASAP7_75t_L g790 ( 
.A1(n_721),
.A2(n_659),
.B(n_664),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_717),
.B(n_354),
.Y(n_791)
);

BUFx4f_ASAP7_75t_L g792 ( 
.A(n_683),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_651),
.B(n_362),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_711),
.B(n_366),
.Y(n_794)
);

AOI21x1_ASAP7_75t_L g795 ( 
.A1(n_681),
.A2(n_489),
.B(n_458),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_710),
.A2(n_436),
.B(n_373),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_668),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_655),
.A2(n_423),
.B(n_376),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_716),
.A2(n_439),
.B(n_385),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_720),
.B(n_369),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_660),
.A2(n_445),
.B(n_390),
.C(n_399),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_665),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_708),
.B(n_388),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_712),
.A2(n_412),
.B(n_414),
.C(n_429),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_706),
.A2(n_591),
.B(n_576),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_715),
.B(n_437),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_644),
.B(n_442),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_699),
.A2(n_591),
.B(n_576),
.Y(n_808)
);

NAND2x1p5_ASAP7_75t_L g809 ( 
.A(n_718),
.B(n_539),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_675),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_759),
.B(n_653),
.Y(n_811)
);

NOR2xp67_ASAP7_75t_L g812 ( 
.A(n_763),
.B(n_677),
.Y(n_812)
);

OAI21x1_ASAP7_75t_SL g813 ( 
.A1(n_745),
.A2(n_645),
.B(n_646),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_733),
.B(n_719),
.Y(n_814)
);

O2A1O1Ixp33_ASAP7_75t_SL g815 ( 
.A1(n_766),
.A2(n_650),
.B(n_674),
.C(n_673),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_750),
.B(n_722),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_784),
.A2(n_726),
.B(n_724),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_731),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_734),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_732),
.B(n_676),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_747),
.A2(n_714),
.B(n_650),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_790),
.B(n_685),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_736),
.B(n_695),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_753),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_758),
.B(n_696),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_800),
.A2(n_703),
.B(n_700),
.C(n_683),
.Y(n_826)
);

AO31x2_ASAP7_75t_L g827 ( 
.A1(n_767),
.A2(n_539),
.A3(n_489),
.B(n_472),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_786),
.Y(n_828)
);

INVx5_ASAP7_75t_L g829 ( 
.A(n_752),
.Y(n_829)
);

AOI21xp33_ASAP7_75t_L g830 ( 
.A1(n_791),
.A2(n_591),
.B(n_574),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_741),
.A2(n_574),
.B(n_489),
.Y(n_831)
);

OA21x2_ASAP7_75t_L g832 ( 
.A1(n_747),
.A2(n_742),
.B(n_771),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_739),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_805),
.A2(n_76),
.B(n_77),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_801),
.A2(n_489),
.B(n_472),
.C(n_458),
.Y(n_835)
);

INVx5_ASAP7_75t_L g836 ( 
.A(n_752),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_738),
.B(n_539),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_788),
.B(n_776),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_755),
.B(n_539),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_756),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_751),
.A2(n_574),
.B(n_472),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_740),
.A2(n_472),
.B(n_458),
.Y(n_842)
);

AOI21x1_ASAP7_75t_L g843 ( 
.A1(n_795),
.A2(n_458),
.B(n_456),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_754),
.B(n_265),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_803),
.B(n_772),
.Y(n_845)
);

AOI21x1_ASAP7_75t_L g846 ( 
.A1(n_743),
.A2(n_78),
.B(n_81),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_760),
.A2(n_86),
.B(n_87),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_778),
.B(n_90),
.Y(n_848)
);

OAI21x1_ASAP7_75t_L g849 ( 
.A1(n_768),
.A2(n_93),
.B(n_94),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_781),
.A2(n_98),
.B(n_104),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_786),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_765),
.A2(n_106),
.B(n_112),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_782),
.A2(n_113),
.B(n_114),
.C(n_115),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_774),
.B(n_126),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_792),
.B(n_127),
.Y(n_855)
);

OA21x2_ASAP7_75t_L g856 ( 
.A1(n_773),
.A2(n_130),
.B(n_131),
.Y(n_856)
);

AO31x2_ASAP7_75t_L g857 ( 
.A1(n_783),
.A2(n_133),
.A3(n_134),
.B(n_138),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_808),
.A2(n_139),
.B(n_149),
.Y(n_858)
);

AOI21x1_ASAP7_75t_L g859 ( 
.A1(n_793),
.A2(n_155),
.B(n_156),
.Y(n_859)
);

AOI21x1_ASAP7_75t_L g860 ( 
.A1(n_787),
.A2(n_157),
.B(n_158),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_764),
.A2(n_159),
.B(n_160),
.Y(n_861)
);

NAND2x1p5_ASAP7_75t_L g862 ( 
.A(n_792),
.B(n_164),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_798),
.A2(n_172),
.B(n_179),
.C(n_180),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_821),
.A2(n_773),
.B(n_809),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_828),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_828),
.B(n_780),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_811),
.B(n_807),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_814),
.B(n_737),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_820),
.A2(n_798),
.B(n_789),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_848),
.A2(n_735),
.B(n_779),
.Y(n_870)
);

NAND2x1p5_ASAP7_75t_L g871 ( 
.A(n_829),
.B(n_749),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_842),
.A2(n_802),
.B(n_785),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_815),
.A2(n_799),
.B(n_796),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_851),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_827),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_834),
.A2(n_809),
.B(n_761),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_817),
.A2(n_774),
.B(n_746),
.Y(n_877)
);

AO21x2_ASAP7_75t_L g878 ( 
.A1(n_822),
.A2(n_769),
.B(n_804),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_851),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_851),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_838),
.B(n_761),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_818),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_850),
.A2(n_757),
.B(n_762),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_824),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_827),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_819),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_816),
.B(n_744),
.Y(n_887)
);

OAI21x1_ASAP7_75t_L g888 ( 
.A1(n_849),
.A2(n_748),
.B(n_797),
.Y(n_888)
);

OAI21x1_ASAP7_75t_SL g889 ( 
.A1(n_852),
.A2(n_806),
.B(n_794),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_854),
.B(n_775),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_827),
.Y(n_891)
);

CKINVDCx16_ASAP7_75t_R g892 ( 
.A(n_845),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_831),
.A2(n_810),
.B(n_777),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_833),
.Y(n_894)
);

AND2x4_ASAP7_75t_SL g895 ( 
.A(n_844),
.B(n_772),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_861),
.A2(n_769),
.B(n_183),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_825),
.Y(n_897)
);

OAI21x1_ASAP7_75t_L g898 ( 
.A1(n_846),
.A2(n_181),
.B(n_189),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_894),
.B(n_829),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_L g900 ( 
.A(n_876),
.B(n_894),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_897),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_875),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_886),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_866),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_884),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_886),
.Y(n_906)
);

OA21x2_ASAP7_75t_L g907 ( 
.A1(n_875),
.A2(n_839),
.B(n_823),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_868),
.B(n_837),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_885),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_865),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_885),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_891),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_865),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_882),
.B(n_829),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_877),
.A2(n_863),
.B(n_812),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_L g916 ( 
.A(n_890),
.B(n_853),
.C(n_770),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_888),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_891),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_878),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_878),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_895),
.B(n_836),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_878),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_874),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_866),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_888),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_896),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_887),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_866),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_903),
.B(n_892),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_915),
.A2(n_890),
.B(n_889),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_902),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_903),
.B(n_867),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_905),
.B(n_840),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_902),
.Y(n_934)
);

NAND2x1p5_ASAP7_75t_SL g935 ( 
.A(n_926),
.B(n_889),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_901),
.B(n_879),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_902),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_910),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_904),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_918),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_910),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_928),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_906),
.B(n_881),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_906),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_914),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_904),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_927),
.B(n_857),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_914),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_927),
.B(n_895),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_909),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_900),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_908),
.B(n_857),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_918),
.B(n_832),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_SL g954 ( 
.A1(n_921),
.A2(n_879),
.B1(n_880),
.B2(n_856),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_908),
.B(n_879),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_900),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_904),
.B(n_880),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_924),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_900),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_924),
.B(n_857),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_924),
.B(n_899),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_909),
.B(n_832),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_942),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_933),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_944),
.B(n_909),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_940),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_940),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_947),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_931),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_952),
.B(n_911),
.Y(n_970)
);

NAND4xp25_ASAP7_75t_L g971 ( 
.A(n_930),
.B(n_916),
.C(n_869),
.D(n_873),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_929),
.B(n_932),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_936),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_952),
.B(n_911),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_945),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_949),
.A2(n_921),
.B1(n_899),
.B2(n_871),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_947),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_929),
.B(n_911),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_932),
.B(n_899),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_931),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_953),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_960),
.B(n_912),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_946),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_960),
.B(n_912),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_955),
.B(n_899),
.Y(n_985)
);

INVxp33_ASAP7_75t_L g986 ( 
.A(n_948),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_953),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_934),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_961),
.B(n_912),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_951),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_934),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_937),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_961),
.B(n_951),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_937),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_962),
.B(n_919),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_943),
.B(n_962),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_943),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_950),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_958),
.B(n_939),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_997),
.B(n_996),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_967),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_967),
.Y(n_1002)
);

OR2x2_ASAP7_75t_L g1003 ( 
.A(n_975),
.B(n_956),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_975),
.B(n_993),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_996),
.B(n_956),
.Y(n_1005)
);

INVx3_ASAP7_75t_SL g1006 ( 
.A(n_964),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_966),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_969),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_963),
.Y(n_1009)
);

NAND4xp25_ASAP7_75t_L g1010 ( 
.A(n_971),
.B(n_938),
.C(n_941),
.D(n_870),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_965),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_993),
.B(n_939),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_981),
.B(n_959),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_973),
.B(n_972),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_990),
.B(n_959),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_965),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_973),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_968),
.B(n_950),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_968),
.B(n_935),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_989),
.B(n_941),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_969),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_986),
.B(n_938),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_999),
.Y(n_1023)
);

INVx1_ASAP7_75t_SL g1024 ( 
.A(n_983),
.Y(n_1024)
);

AND2x4_ASAP7_75t_L g1025 ( 
.A(n_989),
.B(n_941),
.Y(n_1025)
);

AND2x4_ASAP7_75t_SL g1026 ( 
.A(n_989),
.B(n_874),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_978),
.B(n_938),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_977),
.B(n_978),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_999),
.B(n_957),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1000),
.B(n_981),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_1000),
.B(n_977),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_1009),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_1028),
.B(n_987),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_1024),
.A2(n_856),
.B1(n_979),
.B2(n_985),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1014),
.B(n_990),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1004),
.B(n_987),
.Y(n_1036)
);

NAND2x1p5_ASAP7_75t_L g1037 ( 
.A(n_1024),
.B(n_954),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1004),
.B(n_982),
.Y(n_1038)
);

NAND2x1_ASAP7_75t_L g1039 ( 
.A(n_1015),
.B(n_976),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_1006),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1023),
.B(n_982),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1007),
.Y(n_1042)
);

NAND4xp25_ASAP7_75t_L g1043 ( 
.A(n_1019),
.B(n_835),
.C(n_872),
.D(n_893),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1001),
.Y(n_1044)
);

AOI32xp33_ASAP7_75t_SL g1045 ( 
.A1(n_1027),
.A2(n_935),
.A3(n_925),
.B1(n_919),
.B2(n_922),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1002),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1013),
.B(n_995),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1011),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1016),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1013),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1037),
.A2(n_1005),
.B1(n_1029),
.B2(n_1017),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_1032),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_1040),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1032),
.Y(n_1054)
);

OR2x6_ASAP7_75t_L g1055 ( 
.A(n_1039),
.B(n_1015),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_1035),
.B(n_1023),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1031),
.B(n_1005),
.Y(n_1057)
);

INVxp33_ASAP7_75t_L g1058 ( 
.A(n_1038),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_1030),
.B(n_1003),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_1030),
.B(n_1012),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1041),
.B(n_1022),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_1050),
.Y(n_1062)
);

AO22x1_ASAP7_75t_L g1063 ( 
.A1(n_1042),
.A2(n_1025),
.B1(n_1020),
.B2(n_984),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1037),
.A2(n_1015),
.B1(n_1025),
.B2(n_1020),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1036),
.B(n_984),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1044),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_1033),
.B(n_1018),
.Y(n_1067)
);

OAI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_1047),
.A2(n_1010),
.B(n_995),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1034),
.A2(n_1026),
.B1(n_910),
.B2(n_913),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1051),
.A2(n_1068),
.B1(n_1064),
.B2(n_1069),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1066),
.Y(n_1071)
);

OAI221xp5_ASAP7_75t_L g1072 ( 
.A1(n_1055),
.A2(n_1034),
.B1(n_1062),
.B2(n_1047),
.C(n_1066),
.Y(n_1072)
);

AOI211xp5_ASAP7_75t_SL g1073 ( 
.A1(n_1052),
.A2(n_1054),
.B(n_1056),
.C(n_1045),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_1063),
.A2(n_1049),
.B(n_1048),
.C(n_1046),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1059),
.B(n_1043),
.Y(n_1075)
);

AOI221xp5_ASAP7_75t_L g1076 ( 
.A1(n_1067),
.A2(n_1010),
.B1(n_847),
.B2(n_970),
.C(n_974),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1060),
.B(n_970),
.Y(n_1077)
);

O2A1O1Ixp5_ASAP7_75t_L g1078 ( 
.A1(n_1058),
.A2(n_1057),
.B(n_1061),
.C(n_1065),
.Y(n_1078)
);

AOI311xp33_ASAP7_75t_L g1079 ( 
.A1(n_1053),
.A2(n_925),
.A3(n_830),
.B(n_841),
.C(n_826),
.Y(n_1079)
);

AOI211xp5_ASAP7_75t_L g1080 ( 
.A1(n_1055),
.A2(n_923),
.B(n_883),
.C(n_898),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1066),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1061),
.B(n_974),
.Y(n_1082)
);

AOI221xp5_ASAP7_75t_L g1083 ( 
.A1(n_1068),
.A2(n_1021),
.B1(n_1008),
.B2(n_813),
.C(n_920),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1051),
.A2(n_923),
.B1(n_994),
.B2(n_992),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1066),
.Y(n_1085)
);

AOI21xp33_ASAP7_75t_SL g1086 ( 
.A1(n_1053),
.A2(n_913),
.B(n_910),
.Y(n_1086)
);

AOI221xp5_ASAP7_75t_L g1087 ( 
.A1(n_1068),
.A2(n_920),
.B1(n_922),
.B2(n_926),
.C(n_991),
.Y(n_1087)
);

OAI21xp33_ASAP7_75t_L g1088 ( 
.A1(n_1073),
.A2(n_860),
.B(n_913),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1075),
.B(n_980),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1070),
.A2(n_913),
.B1(n_917),
.B2(n_862),
.Y(n_1090)
);

NAND4xp25_ASAP7_75t_L g1091 ( 
.A(n_1073),
.B(n_865),
.C(n_917),
.D(n_992),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1072),
.A2(n_855),
.B(n_871),
.C(n_991),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1074),
.A2(n_883),
.B(n_994),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1084),
.A2(n_998),
.B1(n_988),
.B2(n_980),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_1077),
.B(n_874),
.Y(n_1095)
);

NAND4xp25_ASAP7_75t_L g1096 ( 
.A(n_1076),
.B(n_1078),
.C(n_1080),
.D(n_1079),
.Y(n_1096)
);

AOI222xp33_ASAP7_75t_L g1097 ( 
.A1(n_1087),
.A2(n_998),
.B1(n_988),
.B2(n_898),
.C1(n_896),
.C2(n_864),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_L g1098 ( 
.A(n_1086),
.B(n_859),
.C(n_876),
.Y(n_1098)
);

OAI221xp5_ASAP7_75t_SL g1099 ( 
.A1(n_1083),
.A2(n_871),
.B1(n_858),
.B2(n_864),
.C(n_836),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1081),
.A2(n_907),
.B(n_836),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1085),
.B(n_907),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1071),
.A2(n_907),
.B1(n_843),
.B2(n_199),
.Y(n_1102)
);

NAND4xp75_ASAP7_75t_L g1103 ( 
.A(n_1082),
.B(n_907),
.C(n_194),
.D(n_201),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_1074),
.B(n_191),
.Y(n_1104)
);

AOI211xp5_ASAP7_75t_L g1105 ( 
.A1(n_1072),
.A2(n_202),
.B(n_204),
.C(n_206),
.Y(n_1105)
);

NAND5xp2_ASAP7_75t_L g1106 ( 
.A(n_1088),
.B(n_1105),
.C(n_1092),
.D(n_1096),
.E(n_1091),
.Y(n_1106)
);

NAND4xp25_ASAP7_75t_L g1107 ( 
.A(n_1090),
.B(n_209),
.C(n_211),
.D(n_212),
.Y(n_1107)
);

AOI221xp5_ASAP7_75t_L g1108 ( 
.A1(n_1104),
.A2(n_213),
.B1(n_214),
.B2(n_216),
.C(n_218),
.Y(n_1108)
);

NOR2xp67_ASAP7_75t_L g1109 ( 
.A(n_1101),
.B(n_220),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1095),
.B(n_221),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1106),
.B(n_1089),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_SL g1112 ( 
.A(n_1108),
.B(n_1097),
.C(n_1098),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1109),
.Y(n_1113)
);

NAND4xp25_ASAP7_75t_L g1114 ( 
.A(n_1110),
.B(n_1099),
.C(n_1093),
.D(n_1100),
.Y(n_1114)
);

NOR2x1_ASAP7_75t_L g1115 ( 
.A(n_1107),
.B(n_1103),
.Y(n_1115)
);

NAND4xp75_ASAP7_75t_L g1116 ( 
.A(n_1115),
.B(n_1094),
.C(n_1102),
.D(n_225),
.Y(n_1116)
);

NOR3xp33_ASAP7_75t_L g1117 ( 
.A(n_1112),
.B(n_222),
.C(n_224),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_L g1118 ( 
.A(n_1111),
.B(n_227),
.C(n_230),
.Y(n_1118)
);

NOR3x1_ASAP7_75t_L g1119 ( 
.A(n_1114),
.B(n_231),
.C(n_234),
.Y(n_1119)
);

INVxp67_ASAP7_75t_SL g1120 ( 
.A(n_1119),
.Y(n_1120)
);

XOR2xp5_ASAP7_75t_L g1121 ( 
.A(n_1116),
.B(n_1113),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1117),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1118),
.B(n_235),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1123),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1122),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1125),
.A2(n_1120),
.B1(n_1121),
.B2(n_239),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_1126),
.B(n_1124),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_1127),
.B(n_237),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1128),
.B(n_238),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_1129),
.A2(n_243),
.B(n_244),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1130),
.A2(n_247),
.B1(n_250),
.B2(n_252),
.Y(n_1131)
);


endmodule