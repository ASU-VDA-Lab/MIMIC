module fake_jpeg_27158_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_4),
.B(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_1),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g14 ( 
.A(n_3),
.B(n_5),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_15),
.A2(n_16),
.B1(n_7),
.B2(n_11),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_8),
.B1(n_7),
.B2(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_19),
.Y(n_27)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_6),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_22),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_10),
.A2(n_0),
.B(n_6),
.C(n_5),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_6),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_21),
.B(n_16),
.C(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_20),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_17),
.C(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_25),
.B(n_27),
.Y(n_36)
);

AOI21x1_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_28),
.B(n_26),
.Y(n_35)
);

OAI21x1_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_37),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_39),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_25),
.B(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_30),
.C(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_18),
.B1(n_23),
.B2(n_15),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_20),
.B(n_12),
.C(n_9),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_18),
.B1(n_40),
.B2(n_42),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_SL g47 ( 
.A1(n_46),
.A2(n_45),
.B(n_41),
.C(n_12),
.Y(n_47)
);


endmodule