module fake_netlist_1_244_n_25 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_25);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_25;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
NOR2x1p5_ASAP7_75t_L g11 ( .A(n_2), .B(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_10), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_12), .A2(n_6), .B(n_8), .Y(n_17) );
NAND3xp33_ASAP7_75t_SL g18 ( .A(n_16), .B(n_0), .C(n_1), .Y(n_18) );
NAND3xp33_ASAP7_75t_SL g19 ( .A(n_17), .B(n_13), .C(n_14), .Y(n_19) );
INVx5_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_18), .B1(n_11), .B2(n_13), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
AO22x2_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_20), .B1(n_15), .B2(n_1), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI22xp5_ASAP7_75t_SL g25 ( .A1(n_24), .A2(n_23), .B1(n_7), .B2(n_9), .Y(n_25) );
endmodule