module fake_jpeg_30255_n_104 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_32),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_30),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_19),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_32),
.B1(n_14),
.B2(n_27),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_47),
.B1(n_1),
.B2(n_3),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_53),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_15),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_30),
.A2(n_15),
.B1(n_25),
.B2(n_20),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_55),
.B1(n_1),
.B2(n_2),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_25),
.B1(n_20),
.B2(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_56),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_30),
.A2(n_19),
.B1(n_22),
.B2(n_2),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_28),
.B(n_12),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AND2x6_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_7),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_66),
.Y(n_72)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_9),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_45),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_50),
.B(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_74),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_68),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_87),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_73),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_85),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_76),
.Y(n_87)
);

MAJx2_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_74),
.C(n_79),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_94),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_82),
.B(n_92),
.C(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_94),
.A2(n_84),
.B1(n_78),
.B2(n_61),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_97),
.B1(n_43),
.B2(n_95),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_54),
.B1(n_48),
.B2(n_64),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_97),
.B1(n_96),
.B2(n_98),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_100),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_99),
.Y(n_104)
);


endmodule