module fake_jpeg_23066_n_8 (n_3, n_2, n_1, n_0, n_4, n_8);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_8;

wire n_6;
wire n_5;
wire n_7;

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_1),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

MAJIxp5_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_4),
.C(n_2),
.Y(n_7)
);

NAND4xp25_ASAP7_75t_SL g8 ( 
.A(n_6),
.B(n_0),
.C(n_5),
.D(n_7),
.Y(n_8)
);


endmodule