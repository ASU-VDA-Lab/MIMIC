module fake_jpeg_11605_n_203 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_203);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_54),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_15),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_8),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_24),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_95),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_69),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_1),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_68),
.Y(n_102)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_72),
.B1(n_62),
.B2(n_68),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_104),
.B1(n_107),
.B2(n_79),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_92),
.B(n_66),
.Y(n_116)
);

NAND2x1p5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_62),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_85),
.B1(n_79),
.B2(n_78),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_62),
.B1(n_83),
.B2(n_84),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_83),
.B1(n_60),
.B2(n_74),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_58),
.B1(n_84),
.B2(n_74),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_58),
.B1(n_60),
.B2(n_80),
.Y(n_119)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_81),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_117),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_94),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_71),
.B(n_64),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_134),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_125),
.B1(n_129),
.B2(n_26),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_5),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_70),
.B1(n_65),
.B2(n_67),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_63),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_27),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_77),
.B1(n_76),
.B2(n_85),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_79),
.B1(n_2),
.B2(n_3),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_131),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_136)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_1),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_2),
.B(n_3),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_10),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_147),
.B1(n_153),
.B2(n_43),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_9),
.CI(n_10),
.CON(n_148),
.SN(n_148)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_149),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_11),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_12),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_21),
.C(n_22),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_130),
.B1(n_31),
.B2(n_32),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_148),
.B1(n_156),
.B2(n_170),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_30),
.B(n_33),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_154),
.B(n_136),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_170),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_166),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_50),
.B(n_52),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_156),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_179),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_162),
.B1(n_174),
.B2(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_181),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_143),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_185),
.C(n_164),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_187),
.A2(n_191),
.B1(n_178),
.B2(n_172),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_188),
.A2(n_177),
.B1(n_184),
.B2(n_161),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_181),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_194),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_190),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_186),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_193),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_178),
.Y(n_203)
);


endmodule