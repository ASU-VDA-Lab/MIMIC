module real_jpeg_15709_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_12;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_2),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_2),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_3),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_88)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_93),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_3),
.A2(n_93),
.B1(n_157),
.B2(n_161),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_3),
.A2(n_93),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_4),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_5),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_5),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_5),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_6),
.Y(n_198)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_7),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_7),
.Y(n_123)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_8),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_8),
.A2(n_53),
.B1(n_99),
.B2(n_103),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_8),
.A2(n_47),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_8),
.B(n_178),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_8),
.A2(n_69),
.A3(n_227),
.B1(n_228),
.B2(n_231),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_8),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_8),
.B(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_10),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_219),
.B1(n_309),
.B2(n_310),
.Y(n_12)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_13),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_218),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_183),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_17),
.B(n_183),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.C(n_175),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_18),
.B(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_96),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_55),
.B2(n_56),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_21),
.B(n_55),
.C(n_96),
.Y(n_217)
);

AOI21x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_31),
.B(n_45),
.Y(n_21)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_22),
.Y(n_282)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2x1_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_34),
.Y(n_33)
);

AO22x2_ASAP7_75t_L g193 ( 
.A1(n_23),
.A2(n_33),
.B1(n_46),
.B2(n_194),
.Y(n_193)
);

AO22x1_ASAP7_75t_L g244 ( 
.A1(n_23),
.A2(n_33),
.B1(n_46),
.B2(n_194),
.Y(n_244)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_23)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_25),
.Y(n_155)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_26),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_29),
.Y(n_264)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_36),
.Y(n_200)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_43),
.Y(n_227)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_43),
.Y(n_233)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_48),
.B(n_52),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI32xp33_ASAP7_75t_L g250 ( 
.A1(n_52),
.A2(n_155),
.A3(n_251),
.B1(n_255),
.B2(n_259),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_53),
.B(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_55),
.A2(n_56),
.B1(n_193),
.B2(n_215),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_55),
.B(n_193),
.C(n_225),
.Y(n_302)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_67),
.B1(n_79),
.B2(n_88),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_57),
.A2(n_67),
.B1(n_79),
.B2(n_88),
.Y(n_176)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_63),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_63),
.Y(n_281)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_119),
.B1(n_121),
.B2(n_123),
.Y(n_118)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

NAND2x1p5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_79),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_79),
.Y(n_246)
);

OA22x2_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_84),
.Y(n_254)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_91),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_106),
.B1(n_118),
.B2(n_124),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_98),
.A2(n_106),
.B1(n_118),
.B2(n_124),
.Y(n_187)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21x1_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_113),
.B(n_118),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_128),
.B(n_175),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_149),
.B2(n_150),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_149),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_149),
.A2(n_150),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_150),
.B(n_243),
.C(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_150),
.B(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_150),
.B(n_280),
.Y(n_283)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_156),
.B1(n_164),
.B2(n_168),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_169),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_152),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_156),
.A2(n_180),
.B(n_182),
.Y(n_179)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_160),
.Y(n_174)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_160),
.Y(n_276)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_168),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.C(n_179),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_176),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_176),
.A2(n_186),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_177),
.A2(n_179),
.B1(n_285),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_177),
.Y(n_300)
);

NOR2x1_ASAP7_75t_L g270 ( 
.A(n_179),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_179),
.Y(n_285)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_203),
.B(n_211),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_190),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_189),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_187),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_216),
.B2(n_217),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_201),
.B1(n_202),
.B2(n_215),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_193),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_193),
.B(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_193),
.A2(n_215),
.B1(n_250),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_219),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_304),
.B(n_308),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_291),
.B(n_303),
.Y(n_221)
);

OAI21x1_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_247),
.B(n_290),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_242),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_224),
.B(n_242),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_241),
.Y(n_224)
);

XOR2x2_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_226),
.B(n_234),
.Y(n_294)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_237),
.Y(n_278)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_243),
.A2(n_244),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_243),
.B(n_294),
.C(n_296),
.Y(n_305)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_245),
.Y(n_267)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_268),
.B(n_289),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_265),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_249),
.B(n_265),
.Y(n_289)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_284),
.B(n_288),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_279),
.B(n_283),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp33_ASAP7_75t_SL g288 ( 
.A(n_285),
.B(n_286),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_302),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_302),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_296),
.B1(n_297),
.B2(n_301),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);


endmodule