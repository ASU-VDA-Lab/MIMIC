module real_jpeg_6558_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_1),
.A2(n_150),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_1),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_1),
.A2(n_124),
.B1(n_155),
.B2(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_1),
.A2(n_155),
.B1(n_182),
.B2(n_311),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_1),
.A2(n_155),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_3),
.A2(n_107),
.B1(n_117),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_3),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_3),
.A2(n_121),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g239 ( 
.A1(n_3),
.A2(n_121),
.B1(n_152),
.B2(n_240),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_3),
.A2(n_121),
.B1(n_392),
.B2(n_394),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_4),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_4),
.A2(n_36),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_5),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_5),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_5),
.A2(n_151),
.B1(n_291),
.B2(n_293),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_5),
.A2(n_34),
.B1(n_151),
.B2(n_320),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_5),
.A2(n_151),
.B1(n_378),
.B2(n_380),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_6),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_6),
.A2(n_82),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_6),
.A2(n_82),
.B1(n_218),
.B2(n_221),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_7),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_7),
.A2(n_183),
.B1(n_274),
.B2(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_7),
.B(n_80),
.C(n_282),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_7),
.B(n_108),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_7),
.B(n_326),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_7),
.B(n_90),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_7),
.B(n_387),
.Y(n_386)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_8),
.Y(n_98)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_9),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_9),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_9),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g395 ( 
.A(n_9),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_9),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_10),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_10),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_10),
.A2(n_59),
.B1(n_199),
.B2(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_10),
.A2(n_199),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_10),
.A2(n_199),
.B1(n_293),
.B2(n_416),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_11),
.A2(n_45),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_12),
.Y(n_103)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_13),
.Y(n_134)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_13),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_13),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_13),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_14),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_14),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_14),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_14),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_14),
.Y(n_198)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_14),
.Y(n_201)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_14),
.Y(n_242)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_14),
.Y(n_265)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_16),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_16),
.A2(n_58),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_16),
.A2(n_58),
.B1(n_188),
.B2(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_245),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_244),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_209),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_20),
.B(n_209),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_159),
.C(n_174),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_21),
.B(n_159),
.CI(n_174),
.CON(n_297),
.SN(n_297)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_91),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_22),
.B(n_92),
.C(n_129),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_23),
.B(n_51),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_33),
.B1(n_40),
.B2(n_44),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_24),
.A2(n_44),
.B(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_24),
.A2(n_279),
.B1(n_284),
.B2(n_287),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_24),
.A2(n_319),
.B(n_324),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_24),
.A2(n_274),
.B(n_324),
.Y(n_347)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_25),
.A2(n_187),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_25),
.B(n_327),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_25),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_25),
.A2(n_280),
.B1(n_391),
.B2(n_422),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_31),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_32),
.Y(n_283)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_33),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_43),
.Y(n_286)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_43),
.Y(n_366)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_46),
.Y(n_188)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_47),
.Y(n_329)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_48),
.Y(n_189)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_49),
.Y(n_393)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_50),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_63),
.B1(n_81),
.B2(n_90),
.Y(n_51)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_52),
.Y(n_185)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_57),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_57),
.Y(n_168)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_59),
.Y(n_380)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_65),
.B1(n_67),
.B2(n_70),
.Y(n_64)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_63),
.A2(n_81),
.B1(n_90),
.B2(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_63),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_63),
.A2(n_90),
.B1(n_162),
.B2(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_63),
.B(n_310),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_72),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_72),
.A2(n_334),
.B(n_336),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_77),
.B2(n_79),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_75),
.Y(n_330)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g355 ( 
.A(n_78),
.Y(n_355)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_89),
.Y(n_230)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_89),
.Y(n_312)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_90),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_90),
.B(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_129),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_116),
.B1(n_122),
.B2(n_123),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g204 ( 
.A(n_93),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_93),
.A2(n_122),
.B1(n_290),
.B2(n_415),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_108),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_99),
.B1(n_104),
.B2(n_106),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_102),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g397 ( 
.A(n_102),
.Y(n_397)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_103),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_103),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_SL g404 ( 
.A(n_104),
.B(n_165),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_108),
.Y(n_122)
);

AOI22x1_ASAP7_75t_L g203 ( 
.A1(n_108),
.A2(n_204),
.B1(n_205),
.B2(n_208),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_108),
.A2(n_204),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_113),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g335 ( 
.A(n_110),
.Y(n_335)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_115),
.Y(n_403)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_116),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_122),
.B(n_206),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_122),
.A2(n_415),
.B(n_418),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_123),
.Y(n_216)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_128),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_148),
.B(n_153),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_130),
.A2(n_148),
.B1(n_196),
.B2(n_202),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_131),
.B(n_154),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_131),
.A2(n_438),
.B(n_439),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_141),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_142),
.B1(n_144),
.B2(n_146),
.Y(n_141)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_139),
.Y(n_270)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_152),
.Y(n_276)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_153),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_158),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_158),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_169),
.B2(n_173),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_161),
.B(n_169),
.Y(n_234)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_SL g315 ( 
.A(n_168),
.Y(n_315)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_169),
.A2(n_173),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_194),
.C(n_203),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_175),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_186),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_176),
.B(n_186),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_184),
.B2(n_185),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_177),
.A2(n_307),
.B(n_309),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_177),
.A2(n_184),
.B1(n_334),
.B2(n_377),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_177),
.A2(n_309),
.B(n_377),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_178),
.A2(n_184),
.B(n_336),
.Y(n_442)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_187),
.Y(n_287)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_193),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_194),
.A2(n_195),
.B1(n_203),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_196),
.A2(n_202),
.B(n_243),
.Y(n_256)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g438 ( 
.A1(n_200),
.A2(n_273),
.B(n_274),
.Y(n_438)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_202),
.B(n_274),
.Y(n_420)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_204),
.A2(n_289),
.B(n_296),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_204),
.A2(n_296),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_204),
.B(n_205),
.Y(n_418)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_232),
.B2(n_233),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_222),
.B(n_231),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_223),
.Y(n_231)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g417 ( 
.A(n_220),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_228),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_230),
.Y(n_400)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_298),
.B(n_467),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_297),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_248),
.B(n_297),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.C(n_254),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_253),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_254),
.B(n_457),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.C(n_288),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_255),
.A2(n_256),
.B1(n_288),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_257),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_277),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_258),
.A2(n_277),
.B1(n_278),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_258),
.Y(n_431)
);

OAI32xp33_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_263),
.A3(n_266),
.B1(n_269),
.B2(n_273),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_262),
.Y(n_384)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_SL g383 ( 
.A1(n_274),
.A2(n_384),
.B(n_385),
.Y(n_383)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_288),
.Y(n_452)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_297),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_445),
.B(n_464),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

AOI21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_426),
.B(n_444),
.Y(n_300)
);

AO21x1_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_406),
.B(n_425),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_371),
.B(n_405),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_339),
.B(n_370),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_317),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_305),
.B(n_317),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_313),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_306),
.A2(n_313),
.B1(n_314),
.B2(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_306),
.Y(n_368)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_312),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_331),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_318),
.B(n_332),
.C(n_338),
.Y(n_372)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_322),
.Y(n_394)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_337),
.B2(n_338),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_361),
.B(n_369),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_348),
.B(n_360),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_346),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_359),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_349),
.B(n_359),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_356),
.B(n_358),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_358),
.A2(n_390),
.B(n_395),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_367),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_367),
.Y(n_369)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_373),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_388),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_381),
.B2(n_382),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_381),
.C(n_388),
.Y(n_407)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI32xp33_ASAP7_75t_L g396 ( 
.A1(n_386),
.A2(n_397),
.A3(n_398),
.B1(n_401),
.B2(n_404),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_396),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_396),
.Y(n_412)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx8_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_407),
.B(n_408),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_410),
.B1(n_413),
.B2(n_424),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_412),
.C(n_424),
.Y(n_427)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_413),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_419),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_414),
.B(n_420),
.C(n_421),
.Y(n_432)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_427),
.B(n_428),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_435),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_432),
.B1(n_433),
.B2(n_434),
.Y(n_429)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_430),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_432),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_433),
.C(n_435),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_440),
.B2(n_443),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_441),
.C(n_442),
.Y(n_455)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_440),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_459),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_465),
.B(n_466),
.Y(n_464)
);

NOR2x1_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_456),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_456),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_453),
.C(n_455),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_462),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_453),
.A2(n_454),
.B1(n_455),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_455),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_461),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);


endmodule