module real_jpeg_4539_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_1),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_121),
.B1(n_124),
.B2(n_125),
.Y(n_120)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_1),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_1),
.A2(n_125),
.B1(n_161),
.B2(n_163),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_1),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_1),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_2),
.A2(n_29),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_2),
.A2(n_50),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_50),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_2),
.A2(n_50),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_2),
.A2(n_263),
.B(n_266),
.C(n_269),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_2),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_2),
.B(n_55),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_2),
.B(n_305),
.C(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_2),
.B(n_113),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_2),
.B(n_78),
.C(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_2),
.B(n_31),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_3),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_80),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_3),
.A2(n_80),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_3),
.A2(n_80),
.B1(n_174),
.B2(n_178),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_4),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_4),
.A2(n_28),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_28),
.B1(n_75),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_4),
.A2(n_28),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_5),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_6),
.Y(n_177)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_8),
.Y(n_171)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_8),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_8),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_8),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_9),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_9),
.Y(n_268)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_12),
.Y(n_131)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_13),
.Y(n_305)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_419),
.B(n_421),
.Y(n_19)
);

AO21x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_134),
.B(n_418),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_128),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_22),
.B(n_128),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_119),
.C(n_126),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_23),
.B(n_415),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_52),
.C(n_82),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_24),
.A2(n_142),
.B1(n_143),
.B2(n_156),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_24),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_24),
.B(n_143),
.C(n_157),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_24),
.B(n_244),
.C(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_24),
.A2(n_156),
.B1(n_244),
.B2(n_343),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_24),
.A2(n_156),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_46),
.B2(n_51),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g232 ( 
.A1(n_25),
.A2(n_30),
.B1(n_46),
.B2(n_51),
.Y(n_232)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_29),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_30),
.A2(n_46),
.B1(n_51),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_30),
.A2(n_51),
.B1(n_120),
.B2(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_30),
.A2(n_46),
.B(n_51),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g420 ( 
.A1(n_30),
.A2(n_51),
.B(n_129),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_31)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_32),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_33),
.Y(n_149)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_34),
.Y(n_155)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_40),
.Y(n_123)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_41),
.Y(n_133)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g266 ( 
.A1(n_50),
.A2(n_145),
.B(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_52),
.A2(n_82),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_52),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_52),
.B(n_232),
.C(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_52),
.A2(n_393),
.B1(n_395),
.B2(n_402),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_77),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_53),
.B(n_192),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_65),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_54),
.A2(n_65),
.B1(n_186),
.B2(n_191),
.Y(n_185)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_55),
.A2(n_200),
.B(n_207),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_55),
.B(n_187),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_55),
.A2(n_66),
.B1(n_77),
.B2(n_200),
.Y(n_243)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_68),
.B1(n_71),
.B2(n_74),
.Y(n_67)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_59),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_59),
.Y(n_229)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_59),
.Y(n_276)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_62),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_66),
.B(n_192),
.Y(n_208)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_70),
.Y(n_206)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_76),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_76),
.Y(n_196)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_82),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_90),
.B1(n_113),
.B2(n_114),
.Y(n_82)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_83),
.Y(n_396)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_90),
.B(n_231),
.Y(n_397)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_105),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_91),
.A2(n_105),
.B1(n_144),
.B2(n_150),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_91),
.A2(n_105),
.B1(n_144),
.B2(n_150),
.Y(n_244)
);

NAND2x1_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_105),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_98),
.B1(n_100),
.B2(n_103),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_102),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_105),
.A2(n_396),
.B(n_397),
.Y(n_395)
);

AOI22x1_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_111),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_119),
.B(n_126),
.Y(n_415)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_127),
.B(n_231),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_128),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_128),
.B(n_420),
.Y(n_422)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_413),
.B(n_417),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_384),
.B(n_410),
.Y(n_135)
);

OAI211xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_280),
.B(n_378),
.C(n_383),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_249),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_138),
.A2(n_249),
.B(n_379),
.C(n_382),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_233),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_139),
.B(n_233),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_197),
.C(n_215),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_140),
.B(n_197),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_157),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_142),
.A2(n_143),
.B1(n_218),
.B2(n_299),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_142),
.B(n_299),
.C(n_320),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_142),
.A2(n_143),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_143),
.B(n_232),
.C(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_144),
.Y(n_231)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_155),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_184),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_158),
.A2(n_184),
.B1(n_185),
.B2(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_158),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_164),
.B1(n_172),
.B2(n_181),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_160),
.A2(n_221),
.B(n_224),
.Y(n_220)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_163),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_164),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_165),
.A2(n_226),
.B1(n_272),
.B2(n_277),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_165),
.A2(n_222),
.B1(n_226),
.B2(n_272),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_171),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_210),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_178),
.Y(n_306)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_180),
.Y(n_273)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_184),
.A2(n_185),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_184),
.A2(n_185),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_185),
.B(n_271),
.C(n_313),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_185),
.B(n_335),
.C(n_337),
.Y(n_348)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_209),
.B2(n_214),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_209),
.Y(n_240)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_206),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_209),
.A2(n_214),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_209),
.A2(n_239),
.B(n_240),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_210),
.B(n_226),
.Y(n_328)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_230),
.C(n_232),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_255),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_218),
.A2(n_299),
.B1(n_300),
.B2(n_307),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_218),
.A2(n_220),
.B1(n_299),
.B2(n_369),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_220),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_230),
.A2(n_232),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_232),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_232),
.A2(n_256),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_232),
.A2(n_256),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_232),
.A2(n_256),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_232),
.B(n_389),
.C(n_394),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_247),
.B2(n_248),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_241),
.B1(n_242),
.B2(n_246),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_241),
.B(n_246),
.C(n_248),
.Y(n_409)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_244),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_244),
.A2(n_339),
.B1(n_340),
.B2(n_343),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_244),
.Y(n_343)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_245),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_245),
.A2(n_399),
.B1(n_403),
.B2(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_250),
.B(n_252),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.C(n_260),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_253),
.A2(n_254),
.B1(n_258),
.B2(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_258),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_260),
.B(n_376),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_261),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_270),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_262),
.A2(n_270),
.B1(n_271),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_262),
.Y(n_360)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_271),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_294),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_362),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_347),
.B(n_361),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_332),
.B(n_346),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_317),
.B(n_331),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_309),
.B(n_316),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_296),
.B(n_308),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_293),
.B(n_295),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_292),
.A2(n_297),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_341),
.C(n_343),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_307),
.Y(n_315)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_304),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_315),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_315),
.Y(n_316)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_319),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_330),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_329),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_329),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_345),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_345),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_337),
.B1(n_338),
.B2(n_344),
.Y(n_333)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_349),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_355),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_357),
.C(n_358),
.Y(n_371)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NOR2x1_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_372),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_371),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_371),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_365),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_370),
.C(n_374),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_372),
.A2(n_380),
.B(n_381),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_375),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_405),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_385),
.A2(n_411),
.B(n_412),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_398),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_398),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_394),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_395),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_403),
.C(n_404),
.Y(n_398)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_399),
.Y(n_408)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_407),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_409),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_414),
.B(n_416),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_422),
.Y(n_421)
);


endmodule