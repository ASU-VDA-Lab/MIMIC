module fake_netlist_5_1222_n_1913 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1913);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1913;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_38),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_12),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_125),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_165),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_11),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_85),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_57),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_12),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_55),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_7),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_173),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_75),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_6),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_43),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_47),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_70),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_74),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_77),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_108),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_50),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_91),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_55),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_143),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_32),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_151),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_19),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_56),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_19),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_104),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_39),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_102),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_167),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_78),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_65),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_93),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_30),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_81),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_66),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_170),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_30),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_62),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_61),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_144),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_157),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_56),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_127),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_115),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_149),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_33),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_76),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_24),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_18),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_136),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_94),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_154),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_162),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_178),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_122),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_132),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_54),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_105),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_153),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_126),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_63),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_64),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_67),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_148),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_109),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_158),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_28),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_84),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_174),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_43),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_176),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_45),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_187),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_69),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_134),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_27),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_53),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_86),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_146),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_138),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_59),
.Y(n_284)
);

BUFx2_ASAP7_75t_SL g285 ( 
.A(n_18),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_61),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_79),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_99),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_92),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_161),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_180),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_111),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_49),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_42),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_26),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_66),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_90),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_3),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_37),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_40),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_11),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_128),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_68),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_103),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_37),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_23),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_44),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_181),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_101),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_47),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_40),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_89),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_123),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_57),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_72),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_155),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_141),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_175),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_35),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_112),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_50),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_188),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_21),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_1),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_10),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_20),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_95),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_140),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_51),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_29),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_82),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_80),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_58),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_60),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_135),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_17),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_15),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_1),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_4),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_87),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_117),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_147),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_9),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_35),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_25),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_177),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_33),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_124),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_16),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_150),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_14),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_114),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_45),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_8),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_27),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_83),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_113),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_2),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_32),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_34),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_133),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_88),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_159),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_156),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_106),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_63),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_121),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_0),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_6),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_26),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_24),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_15),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_168),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_3),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_8),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_25),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_120),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_228),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_259),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_259),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_191),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_189),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_191),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_315),
.B(n_0),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_298),
.B(n_2),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_261),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_259),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_259),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_194),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_250),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_259),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_305),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_203),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_204),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_221),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_209),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_289),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_298),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_217),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_225),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_198),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_300),
.B(n_4),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_201),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_227),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_297),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_305),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_305),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_198),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_199),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_199),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_202),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_315),
.B(n_5),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_192),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_193),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_202),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_237),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_197),
.B(n_5),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_195),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_268),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_196),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_212),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_238),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_256),
.B(n_7),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_212),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_239),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_213),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_213),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_263),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_272),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_256),
.B(n_9),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_298),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_214),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_205),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_274),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_278),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_214),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_206),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_300),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_245),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_275),
.B(n_10),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_284),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_305),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_208),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_305),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_293),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_211),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_296),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_245),
.Y(n_449)
);

INVxp33_ASAP7_75t_SL g450 ( 
.A(n_299),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_215),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_298),
.Y(n_452)
);

NOR2xp67_ASAP7_75t_L g453 ( 
.A(n_345),
.B(n_13),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_306),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_275),
.B(n_13),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_257),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_257),
.B(n_14),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_267),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_190),
.B(n_16),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_216),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_218),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_267),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_288),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_288),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_307),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_347),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_347),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_314),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_319),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_347),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_303),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_220),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_285),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_402),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_402),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_402),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_402),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_379),
.Y(n_478)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_402),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

CKINVDCx11_ASAP7_75t_R g481 ( 
.A(n_378),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_385),
.A2(n_353),
.B1(n_330),
.B2(n_333),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_409),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_409),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_409),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_386),
.B(n_265),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_420),
.B(n_439),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_391),
.B(n_347),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_380),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_380),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_388),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_399),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_399),
.B(n_265),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_432),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_432),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_452),
.Y(n_500)
);

CKINVDCx8_ASAP7_75t_R g501 ( 
.A(n_382),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_439),
.B(n_265),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_452),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_473),
.B(n_248),
.Y(n_505)
);

OA21x2_ASAP7_75t_L g506 ( 
.A1(n_392),
.A2(n_309),
.B(n_303),
.Y(n_506)
);

AND3x1_ASAP7_75t_L g507 ( 
.A(n_418),
.B(n_210),
.C(n_190),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_392),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_393),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_408),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_443),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_403),
.B(n_198),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_443),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_403),
.B(n_248),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_445),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_414),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_424),
.B(n_198),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_466),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_415),
.A2(n_337),
.B1(n_321),
.B2(n_374),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_466),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_396),
.B(n_301),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_467),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_450),
.B(n_413),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_467),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_470),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_470),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_381),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_384),
.B(n_302),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_411),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_412),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_422),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_431),
.B(n_285),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_425),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_427),
.B(n_302),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_433),
.B(n_301),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_437),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_440),
.B(n_291),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_SL g546 ( 
.A(n_441),
.B(n_210),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_449),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_456),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_458),
.A2(n_316),
.B(n_309),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_462),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_463),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_464),
.B(n_471),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_528),
.B(n_419),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_496),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_550),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_550),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_496),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_496),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_490),
.B(n_421),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_395),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_496),
.B(n_316),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_550),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_550),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_532),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_532),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_481),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_529),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_L g568 ( 
.A(n_522),
.B(n_198),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_501),
.B(n_434),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_534),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_524),
.B(n_382),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_526),
.B(n_390),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_489),
.B(n_438),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_522),
.B(n_262),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_507),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_534),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_533),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_535),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_522),
.A2(n_457),
.B1(n_455),
.B2(n_347),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_518),
.B(n_486),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_529),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_503),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_474),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_474),
.Y(n_584)
);

OR2x6_ASAP7_75t_L g585 ( 
.A(n_539),
.B(n_453),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_505),
.B(n_444),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_535),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_537),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_510),
.Y(n_589)
);

INVxp33_ASAP7_75t_L g590 ( 
.A(n_543),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_543),
.B(n_423),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_474),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_474),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_474),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_518),
.B(n_390),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_537),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_L g597 ( 
.A(n_522),
.B(n_262),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_518),
.B(n_394),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_540),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_552),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_491),
.Y(n_601)
);

INVx5_ASAP7_75t_L g602 ( 
.A(n_516),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_518),
.B(n_394),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_533),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_474),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_540),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_542),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_539),
.B(n_404),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_501),
.B(n_397),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_516),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_483),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_483),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_482),
.B(n_447),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_539),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_539),
.B(n_376),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_486),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_539),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_491),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_541),
.B(n_451),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_491),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_486),
.B(n_522),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_542),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_502),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_552),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_486),
.B(n_291),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_533),
.B(n_317),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_502),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_547),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_521),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_547),
.B(n_317),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

AND2x6_ASAP7_75t_L g632 ( 
.A(n_545),
.B(n_312),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_522),
.B(n_400),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_502),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_510),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_478),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_516),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_480),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_476),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_522),
.B(n_400),
.Y(n_640)
);

XOR2xp5_ASAP7_75t_L g641 ( 
.A(n_521),
.B(n_387),
.Y(n_641)
);

INVx8_ASAP7_75t_L g642 ( 
.A(n_516),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_546),
.Y(n_643)
);

AND2x6_ASAP7_75t_L g644 ( 
.A(n_545),
.B(n_312),
.Y(n_644)
);

NAND2xp33_ASAP7_75t_SL g645 ( 
.A(n_545),
.B(n_401),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_549),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_480),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_492),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_510),
.Y(n_649)
);

NOR2x1p5_ASAP7_75t_L g650 ( 
.A(n_536),
.B(n_200),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_511),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_511),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_492),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_511),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_493),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_512),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_512),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_522),
.A2(n_376),
.B1(n_459),
.B2(n_326),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_516),
.A2(n_200),
.B1(n_326),
.B2(n_383),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_512),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_493),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_536),
.B(n_426),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_545),
.B(n_544),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_544),
.B(n_548),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_494),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_494),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_499),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_548),
.B(n_499),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_548),
.B(n_454),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_549),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_549),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_508),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_508),
.Y(n_673)
);

AND3x2_ASAP7_75t_L g674 ( 
.A(n_509),
.B(n_322),
.C(n_346),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_538),
.B(n_460),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_516),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_509),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_516),
.A2(n_249),
.B1(n_323),
.B2(n_324),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_483),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_538),
.B(n_405),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_538),
.B(n_461),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_483),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_513),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_513),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_510),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_538),
.B(n_417),
.Y(n_686)
);

XOR2xp5_ASAP7_75t_L g687 ( 
.A(n_549),
.B(n_398),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_516),
.B(n_551),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_514),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_551),
.B(n_472),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_551),
.B(n_417),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_551),
.A2(n_339),
.B1(n_224),
.B2(n_344),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_483),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_514),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_483),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_551),
.B(n_429),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_551),
.B(n_429),
.Y(n_697)
);

BUFx4f_ASAP7_75t_L g698 ( 
.A(n_506),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_484),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_517),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_517),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_506),
.A2(n_469),
.B1(n_430),
.B2(n_465),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_582),
.B(n_430),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_590),
.B(n_435),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_616),
.B(n_637),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_625),
.B(n_222),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_554),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_662),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_L g709 ( 
.A(n_553),
.B(n_436),
.C(n_435),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_591),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_616),
.B(n_637),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_554),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_577),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_691),
.B(n_697),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_557),
.Y(n_715)
);

BUFx5_ASAP7_75t_L g716 ( 
.A(n_646),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_580),
.B(n_436),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_557),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_577),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_663),
.B(n_442),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_663),
.B(n_446),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_560),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_702),
.A2(n_406),
.B1(n_469),
.B2(n_446),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_560),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_604),
.B(n_564),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_637),
.B(n_262),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_608),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_558),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_573),
.B(n_465),
.C(n_448),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_600),
.A2(n_249),
.B(n_323),
.C(n_310),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_604),
.B(n_448),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_591),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_572),
.B(n_468),
.Y(n_733)
);

AO221x1_ASAP7_75t_L g734 ( 
.A1(n_575),
.A2(n_262),
.B1(n_223),
.B2(n_231),
.C(n_233),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_613),
.A2(n_271),
.B1(n_251),
.B2(n_308),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_564),
.B(n_565),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_669),
.B(n_250),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_595),
.B(n_325),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_601),
.Y(n_739)
);

AND2x2_ASAP7_75t_SL g740 ( 
.A(n_568),
.B(n_346),
.Y(n_740)
);

NOR3xp33_ASAP7_75t_L g741 ( 
.A(n_571),
.B(n_334),
.C(n_329),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_569),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_L g743 ( 
.A(n_624),
.B(n_338),
.C(n_336),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_598),
.B(n_343),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_558),
.Y(n_745)
);

OAI221xp5_ASAP7_75t_L g746 ( 
.A1(n_579),
.A2(n_576),
.B1(n_578),
.B2(n_570),
.C(n_565),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_570),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_637),
.B(n_262),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_576),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_637),
.B(n_497),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_637),
.B(n_497),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_602),
.B(n_497),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_670),
.A2(n_646),
.B1(n_671),
.B2(n_698),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_578),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_602),
.B(n_497),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_670),
.A2(n_506),
.B1(n_233),
.B2(n_354),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_602),
.B(n_497),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_587),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_587),
.B(n_519),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_588),
.B(n_519),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_588),
.B(n_520),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_614),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_596),
.Y(n_763)
);

INVxp33_ASAP7_75t_L g764 ( 
.A(n_669),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_596),
.B(n_520),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_599),
.B(n_523),
.Y(n_766)
);

AOI221xp5_ASAP7_75t_L g767 ( 
.A1(n_692),
.A2(n_280),
.B1(n_294),
.B2(n_207),
.C(n_219),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_662),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_601),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_599),
.B(n_523),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_606),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_603),
.A2(n_362),
.B1(n_356),
.B2(n_341),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_608),
.B(n_349),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_618),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_586),
.B(n_359),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_606),
.B(n_525),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_607),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_607),
.B(n_622),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_650),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_SL g780 ( 
.A(n_559),
.B(n_247),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_622),
.B(n_525),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_633),
.A2(n_362),
.B1(n_356),
.B2(n_341),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_628),
.B(n_527),
.Y(n_783)
);

NOR3xp33_ASAP7_75t_L g784 ( 
.A(n_619),
.B(n_366),
.C(n_360),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_618),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_676),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_628),
.B(n_527),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_696),
.B(n_369),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_664),
.B(n_531),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_698),
.A2(n_264),
.B(n_223),
.C(n_375),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_602),
.B(n_610),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_620),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_632),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_675),
.B(n_495),
.Y(n_794)
);

NAND3xp33_ASAP7_75t_L g795 ( 
.A(n_645),
.B(n_371),
.C(n_370),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_620),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_602),
.B(n_497),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_623),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_681),
.A2(n_260),
.B1(n_234),
.B2(n_232),
.Y(n_799)
);

OAI22xp33_ASAP7_75t_L g800 ( 
.A1(n_585),
.A2(n_264),
.B1(n_324),
.B2(n_310),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_664),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_668),
.B(n_531),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_585),
.A2(n_269),
.B1(n_351),
.B2(n_242),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_610),
.B(n_498),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_668),
.B(n_506),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_671),
.B(n_498),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_690),
.B(n_328),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_631),
.B(n_498),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_631),
.B(n_498),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_609),
.B(n_250),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_650),
.B(n_328),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_636),
.B(n_498),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_575),
.B(n_342),
.Y(n_813)
);

OAI221xp5_ASAP7_75t_L g814 ( 
.A1(n_678),
.A2(n_269),
.B1(n_242),
.B2(n_235),
.C(n_231),
.Y(n_814)
);

CKINVDCx16_ASAP7_75t_R g815 ( 
.A(n_641),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_626),
.B(n_342),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_617),
.B(n_250),
.Y(n_817)
);

AO22x1_ASAP7_75t_L g818 ( 
.A1(n_617),
.A2(n_235),
.B1(n_221),
.B2(n_286),
.Y(n_818)
);

INVxp33_ASAP7_75t_L g819 ( 
.A(n_641),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_585),
.Y(n_820)
);

BUFx6f_ASAP7_75t_SL g821 ( 
.A(n_615),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_626),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_L g823 ( 
.A(n_640),
.B(n_495),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_626),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_680),
.B(n_348),
.C(n_350),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_561),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_630),
.B(n_279),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_561),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_623),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_658),
.A2(n_348),
.B1(n_350),
.B2(n_357),
.Y(n_830)
);

NAND3xp33_ASAP7_75t_L g831 ( 
.A(n_686),
.B(n_357),
.C(n_361),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_636),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_627),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_638),
.Y(n_834)
);

INVx8_ASAP7_75t_L g835 ( 
.A(n_585),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_627),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_610),
.B(n_698),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_634),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_647),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_647),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_648),
.B(n_498),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_648),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_610),
.B(n_621),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_653),
.B(n_500),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_653),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_615),
.B(n_361),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_655),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_655),
.B(n_500),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_661),
.B(n_665),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_661),
.B(n_500),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_665),
.B(n_500),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_677),
.B(n_500),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_630),
.A2(n_561),
.B(n_295),
.C(n_351),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_677),
.B(n_500),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_634),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_689),
.Y(n_856)
);

OAI22xp33_ASAP7_75t_L g857 ( 
.A1(n_615),
.A2(n_286),
.B1(n_295),
.B2(n_354),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_689),
.B(n_504),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_555),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_555),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_687),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_556),
.B(n_562),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_556),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_651),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_687),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_676),
.B(n_504),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_562),
.B(n_504),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_563),
.B(n_504),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_615),
.B(n_355),
.Y(n_869)
);

OAI22xp33_ASAP7_75t_L g870 ( 
.A1(n_630),
.A2(n_355),
.B1(n_368),
.B2(n_372),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_716),
.B(n_676),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_713),
.Y(n_872)
);

O2A1O1Ixp5_ASAP7_75t_L g873 ( 
.A1(n_807),
.A2(n_639),
.B(n_688),
.C(n_563),
.Y(n_873)
);

AOI21x1_ASAP7_75t_L g874 ( 
.A1(n_705),
.A2(n_667),
.B(n_666),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_714),
.A2(n_805),
.B(n_753),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_SL g876 ( 
.A(n_780),
.B(n_566),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_753),
.A2(n_642),
.B(n_574),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_758),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_807),
.A2(n_659),
.B(n_377),
.C(n_700),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_768),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_764),
.B(n_629),
.Y(n_881)
);

NOR2x1_ASAP7_75t_L g882 ( 
.A(n_729),
.B(n_643),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_713),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_806),
.A2(n_725),
.B(n_843),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_758),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_779),
.B(n_674),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_790),
.A2(n_701),
.B(n_700),
.C(n_667),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_764),
.B(n_629),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_713),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_713),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_843),
.A2(n_642),
.B(n_574),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_771),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_837),
.A2(n_642),
.B(n_597),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_837),
.A2(n_642),
.B(n_597),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_815),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_788),
.B(n_666),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_703),
.B(n_566),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_866),
.A2(n_568),
.B(n_589),
.Y(n_898)
);

OAI21xp33_ASAP7_75t_L g899 ( 
.A1(n_775),
.A2(n_813),
.B(n_737),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_866),
.A2(n_635),
.B(n_589),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_869),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_821),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_719),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_821),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_788),
.B(n_775),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_786),
.A2(n_635),
.B(n_589),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_704),
.B(n_672),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_786),
.A2(n_649),
.B(n_635),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_786),
.A2(n_685),
.B(n_649),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_727),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_716),
.B(n_672),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_822),
.B(n_673),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_786),
.A2(n_685),
.B(n_649),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_771),
.B(n_673),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_859),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_801),
.B(n_683),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_860),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_794),
.A2(n_685),
.B(n_605),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_863),
.Y(n_919)
);

O2A1O1Ixp5_ASAP7_75t_L g920 ( 
.A1(n_736),
.A2(n_694),
.B(n_683),
.C(n_684),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_716),
.B(n_684),
.Y(n_921)
);

AND2x6_ASAP7_75t_L g922 ( 
.A(n_793),
.B(n_694),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_832),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_719),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_719),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_SL g926 ( 
.A1(n_790),
.A2(n_581),
.B(n_567),
.C(n_375),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_756),
.A2(n_625),
.B(n_651),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_747),
.B(n_625),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_710),
.A2(n_581),
.B(n_567),
.C(n_652),
.Y(n_929)
);

OAI22xp5_ASAP7_75t_L g930 ( 
.A1(n_756),
.A2(n_276),
.B1(n_373),
.B2(n_367),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_710),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_808),
.A2(n_652),
.B(n_654),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_722),
.B(n_724),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_739),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_809),
.A2(n_841),
.B(n_812),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_719),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_853),
.A2(n_654),
.B(n_656),
.C(n_657),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_834),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_762),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_862),
.A2(n_625),
.B(n_656),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_844),
.A2(n_657),
.B(n_660),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_749),
.B(n_754),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_738),
.A2(n_660),
.B(n_695),
.C(n_693),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_763),
.B(n_625),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_704),
.B(n_732),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_817),
.B(n_279),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_716),
.B(n_226),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_705),
.A2(n_475),
.B(n_477),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_848),
.A2(n_699),
.B(n_695),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_777),
.B(n_625),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_746),
.A2(n_625),
.B(n_632),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_711),
.A2(n_699),
.B(n_695),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_716),
.B(n_229),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_824),
.A2(n_255),
.B1(n_365),
.B2(n_364),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_745),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_769),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_716),
.B(n_230),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_835),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_762),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_839),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_745),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_R g962 ( 
.A(n_835),
.B(n_632),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_835),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_840),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_850),
.A2(n_852),
.B(n_851),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_842),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_774),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_742),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_717),
.B(n_699),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_785),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_826),
.Y(n_971)
);

AOI21xp33_ASAP7_75t_L g972 ( 
.A1(n_733),
.A2(n_254),
.B(n_236),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_791),
.A2(n_584),
.B(n_605),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_791),
.A2(n_584),
.B(n_605),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_792),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_845),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_823),
.A2(n_584),
.B(n_605),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_711),
.A2(n_802),
.B(n_789),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_828),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_720),
.Y(n_980)
);

AO21x1_ASAP7_75t_L g981 ( 
.A1(n_782),
.A2(n_372),
.B(n_475),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_707),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_718),
.A2(n_584),
.B(n_605),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_SL g984 ( 
.A(n_861),
.B(n_279),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_847),
.B(n_632),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_856),
.B(n_632),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_778),
.B(n_632),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_854),
.A2(n_693),
.B(n_682),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_738),
.A2(n_744),
.B1(n_712),
.B2(n_715),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_858),
.A2(n_693),
.B(n_682),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_728),
.A2(n_682),
.B(n_583),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_849),
.B(n_632),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_744),
.B(n_644),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_867),
.A2(n_868),
.B(n_721),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_733),
.B(n_583),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_731),
.B(n_583),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_723),
.B(n_592),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_759),
.A2(n_592),
.B(n_612),
.Y(n_998)
);

OAI21xp33_ASAP7_75t_L g999 ( 
.A1(n_813),
.A2(n_246),
.B(n_240),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_760),
.A2(n_765),
.B(n_761),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_796),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_793),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_816),
.B(n_644),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_735),
.B(n_592),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_784),
.B(n_241),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_816),
.B(n_644),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_766),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_770),
.A2(n_593),
.B(n_612),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_776),
.A2(n_593),
.B(n_612),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_853),
.A2(n_593),
.B(n_594),
.C(n_611),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_810),
.B(n_279),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_709),
.B(n_243),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_706),
.A2(n_679),
.B(n_584),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_752),
.A2(n_757),
.B(n_755),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_752),
.A2(n_679),
.B(n_611),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_781),
.A2(n_611),
.B(n_594),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_783),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_787),
.B(n_644),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_820),
.B(n_644),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_740),
.A2(n_332),
.B1(n_252),
.B2(n_253),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_755),
.A2(n_594),
.B(n_679),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_846),
.A2(n_644),
.B1(n_331),
.B2(n_327),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_757),
.A2(n_679),
.B(n_484),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_798),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_800),
.B(n_244),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_829),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_833),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_836),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_838),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_797),
.A2(n_679),
.B(n_484),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_855),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_800),
.B(n_258),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_797),
.A2(n_488),
.B(n_484),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_827),
.B(n_644),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_864),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_740),
.A2(n_475),
.B(n_477),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_804),
.A2(n_488),
.B(n_484),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_804),
.A2(n_488),
.B(n_484),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_750),
.A2(n_488),
.B(n_485),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_811),
.Y(n_1040)
);

AOI22x1_ASAP7_75t_L g1041 ( 
.A1(n_811),
.A2(n_320),
.B1(n_270),
.B2(n_273),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_750),
.A2(n_488),
.B(n_485),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_751),
.A2(n_488),
.B(n_485),
.Y(n_1043)
);

O2A1O1Ixp5_ASAP7_75t_L g1044 ( 
.A1(n_772),
.A2(n_477),
.B(n_487),
.C(n_495),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_803),
.B(n_266),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_751),
.A2(n_485),
.B(n_476),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_865),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_773),
.A2(n_335),
.B1(n_281),
.B2(n_282),
.Y(n_1048)
);

INVx4_ASAP7_75t_L g1049 ( 
.A(n_818),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_730),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_SL g1051 ( 
.A(n_819),
.B(n_311),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_846),
.A2(n_487),
.B(n_476),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_743),
.B(n_277),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_799),
.B(n_803),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_825),
.A2(n_487),
.B(n_476),
.Y(n_1055)
);

BUFx8_ASAP7_75t_L g1056 ( 
.A(n_767),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_726),
.A2(n_485),
.B(n_504),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_726),
.A2(n_485),
.B(n_504),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_831),
.B(n_495),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_870),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_961),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_905),
.B(n_857),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1007),
.B(n_857),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_899),
.B(n_741),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_R g1065 ( 
.A(n_895),
.B(n_283),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_875),
.A2(n_951),
.B(n_987),
.Y(n_1066)
);

CKINVDCx16_ASAP7_75t_R g1067 ( 
.A(n_876),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1054),
.A2(n_795),
.B1(n_830),
.B2(n_814),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_968),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_939),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_883),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_923),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_1047),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1017),
.B(n_870),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_875),
.A2(n_748),
.B(n_734),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_945),
.B(n_748),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_989),
.A2(n_877),
.B1(n_907),
.B2(n_995),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_992),
.A2(n_510),
.B(n_530),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1049),
.B(n_287),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1018),
.A2(n_530),
.B(n_515),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_883),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_980),
.B(n_942),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_919),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_1049),
.B(n_290),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_892),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1026),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_883),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_971),
.B(n_318),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_978),
.A2(n_530),
.B(n_515),
.Y(n_1089)
);

OAI21xp33_ASAP7_75t_L g1090 ( 
.A1(n_984),
.A2(n_340),
.B(n_304),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_946),
.B(n_881),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_SL g1092 ( 
.A1(n_1053),
.A2(n_292),
.B(n_363),
.C(n_352),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_SL g1093 ( 
.A(n_897),
.B(n_963),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_971),
.B(n_313),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_993),
.A2(n_1000),
.B(n_884),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_972),
.A2(n_311),
.B(n_20),
.C(n_21),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_938),
.B(n_530),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1000),
.A2(n_515),
.B(n_510),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1026),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_910),
.B(n_311),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_927),
.A2(n_530),
.B(n_515),
.Y(n_1101)
);

CKINVDCx16_ASAP7_75t_R g1102 ( 
.A(n_1051),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_971),
.B(n_311),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_960),
.B(n_530),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_888),
.B(n_17),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_964),
.B(n_515),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_896),
.A2(n_479),
.B(n_184),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_959),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_SL g1109 ( 
.A(n_963),
.B(n_479),
.Y(n_1109)
);

OAI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_933),
.A2(n_901),
.B1(n_1060),
.B2(n_1040),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_966),
.B(n_22),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_976),
.B(n_22),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_917),
.B(n_23),
.Y(n_1113)
);

INVx6_ASAP7_75t_L g1114 ( 
.A(n_958),
.Y(n_1114)
);

AOI221xp5_ASAP7_75t_L g1115 ( 
.A1(n_1050),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.C(n_34),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_SL g1116 ( 
.A(n_1011),
.B(n_31),
.C(n_36),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_931),
.B(n_36),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1056),
.A2(n_479),
.B1(n_39),
.B2(n_41),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_912),
.B(n_38),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_934),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_979),
.B(n_98),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_940),
.A2(n_479),
.B(n_97),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_997),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_979),
.B(n_1056),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_952),
.A2(n_110),
.B(n_182),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_916),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_958),
.B(n_479),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_880),
.B(n_46),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_956),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1024),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1025),
.A2(n_46),
.B(n_48),
.C(n_51),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_912),
.B(n_48),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_967),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_882),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_879),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_SL g1136 ( 
.A(n_902),
.B(n_52),
.C(n_58),
.Y(n_1136)
);

INVx3_ASAP7_75t_SL g1137 ( 
.A(n_904),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_994),
.A2(n_119),
.B(n_171),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_948),
.A2(n_118),
.B(n_169),
.Y(n_1139)
);

BUFx5_ASAP7_75t_L g1140 ( 
.A(n_922),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_874),
.A2(n_116),
.B(n_164),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1004),
.A2(n_100),
.B1(n_160),
.B2(n_142),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_958),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_994),
.A2(n_96),
.B(n_139),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_886),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_886),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_969),
.A2(n_1034),
.B(n_999),
.C(n_996),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1048),
.B(n_59),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1032),
.A2(n_60),
.B(n_62),
.C(n_64),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1002),
.A2(n_71),
.B1(n_130),
.B2(n_131),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_982),
.B(n_65),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1029),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1045),
.B(n_137),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_889),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1035),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_887),
.A2(n_172),
.B(n_944),
.C(n_928),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_982),
.B(n_1012),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_1005),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_878),
.B(n_885),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_890),
.B(n_1019),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_R g1161 ( 
.A(n_872),
.B(n_903),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1019),
.A2(n_1003),
.B1(n_1006),
.B2(n_1002),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_961),
.B(n_955),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_955),
.B(n_914),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_970),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_930),
.A2(n_1020),
.B(n_954),
.C(n_926),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_873),
.A2(n_920),
.B(n_965),
.Y(n_1167)
);

AO32x1_ASAP7_75t_L g1168 ( 
.A1(n_975),
.A2(n_1028),
.A3(n_1027),
.B1(n_1001),
.B2(n_1031),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_935),
.A2(n_965),
.B(n_1013),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_935),
.A2(n_950),
.B(n_894),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_893),
.A2(n_894),
.B(n_918),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_937),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_962),
.B(n_936),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_893),
.A2(n_891),
.B(n_986),
.Y(n_1174)
);

O2A1O1Ixp5_ASAP7_75t_L g1175 ( 
.A1(n_947),
.A2(n_957),
.B(n_953),
.C(n_943),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_872),
.Y(n_1176)
);

OR2x6_ASAP7_75t_SL g1177 ( 
.A(n_1059),
.B(n_985),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_891),
.A2(n_1010),
.B(n_929),
.C(n_898),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_903),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_924),
.B(n_936),
.Y(n_1180)
);

NAND2x1_ASAP7_75t_L g1181 ( 
.A(n_922),
.B(n_925),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_925),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1052),
.B(n_1055),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1044),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1036),
.A2(n_921),
.B(n_911),
.C(n_1008),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_922),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1041),
.B(n_1022),
.C(n_1014),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_922),
.A2(n_871),
.B1(n_981),
.B2(n_898),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_L g1189 ( 
.A(n_922),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1021),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_998),
.A2(n_1008),
.B(n_1016),
.C(n_1009),
.Y(n_1191)
);

OAI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_998),
.A2(n_1009),
.B1(n_1016),
.B2(n_991),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_932),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_991),
.B(n_990),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_1039),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_932),
.B(n_941),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_941),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_949),
.A2(n_990),
.B(n_988),
.C(n_983),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_949),
.B(n_988),
.Y(n_1199)
);

CKINVDCx14_ASAP7_75t_R g1200 ( 
.A(n_1046),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_906),
.A2(n_908),
.B(n_909),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1021),
.A2(n_1015),
.B(n_900),
.C(n_973),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1023),
.A2(n_1030),
.B1(n_1039),
.B2(n_1037),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_913),
.B(n_1023),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_977),
.A2(n_974),
.B(n_1030),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_SL g1206 ( 
.A(n_1057),
.B(n_1058),
.Y(n_1206)
);

NOR3xp33_ASAP7_75t_L g1207 ( 
.A(n_1057),
.B(n_1058),
.C(n_1037),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1033),
.A2(n_1038),
.B1(n_1042),
.B2(n_1043),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_961),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_905),
.B(n_553),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_905),
.A2(n_875),
.B(n_714),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_SL g1212 ( 
.A1(n_905),
.A2(n_807),
.B(n_775),
.C(n_681),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_915),
.Y(n_1213)
);

INVx3_ASAP7_75t_L g1214 ( 
.A(n_1061),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1143),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1210),
.B(n_1126),
.Y(n_1216)
);

BUFx4f_ASAP7_75t_SL g1217 ( 
.A(n_1137),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1091),
.A2(n_1134),
.B1(n_1148),
.B2(n_1067),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1191),
.A2(n_1194),
.A3(n_1169),
.B(n_1095),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1211),
.A2(n_1095),
.B(n_1169),
.Y(n_1220)
);

OAI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1102),
.A2(n_1062),
.B1(n_1093),
.B2(n_1063),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1171),
.A2(n_1205),
.B(n_1201),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1189),
.B(n_1061),
.Y(n_1223)
);

BUFx10_ASAP7_75t_L g1224 ( 
.A(n_1128),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1171),
.A2(n_1205),
.B(n_1201),
.Y(n_1225)
);

INVxp67_ASAP7_75t_SL g1226 ( 
.A(n_1070),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_SL g1227 ( 
.A1(n_1199),
.A2(n_1151),
.B(n_1112),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1108),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1105),
.B(n_1117),
.Y(n_1229)
);

INVx4_ASAP7_75t_L g1230 ( 
.A(n_1114),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1077),
.B(n_1076),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1158),
.A2(n_1153),
.B1(n_1157),
.B2(n_1064),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1211),
.A2(n_1147),
.B(n_1170),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1130),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1082),
.B(n_1146),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1089),
.A2(n_1098),
.B(n_1174),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1209),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1074),
.B(n_1110),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1152),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1083),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1170),
.A2(n_1066),
.B(n_1174),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1089),
.A2(n_1098),
.B(n_1078),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1212),
.B(n_1172),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1066),
.A2(n_1204),
.B(n_1196),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1155),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1213),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1178),
.A2(n_1075),
.A3(n_1122),
.B(n_1156),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1075),
.A2(n_1122),
.A3(n_1184),
.B(n_1193),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_SL g1249 ( 
.A1(n_1166),
.A2(n_1183),
.B(n_1185),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1167),
.A2(n_1202),
.B(n_1187),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1101),
.A2(n_1175),
.B(n_1068),
.Y(n_1251)
);

AND2x6_ASAP7_75t_SL g1252 ( 
.A(n_1100),
.B(n_1119),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1101),
.A2(n_1078),
.B(n_1080),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1123),
.A2(n_1092),
.B(n_1121),
.C(n_1181),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_SL g1255 ( 
.A1(n_1079),
.A2(n_1084),
.B(n_1115),
.C(n_1163),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_SL g1256 ( 
.A1(n_1115),
.A2(n_1111),
.B(n_1113),
.C(n_1164),
.Y(n_1256)
);

INVx4_ASAP7_75t_L g1257 ( 
.A(n_1114),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1192),
.A2(n_1198),
.B(n_1189),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_SL g1259 ( 
.A(n_1186),
.B(n_1069),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1162),
.A2(n_1200),
.B1(n_1118),
.B2(n_1132),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1197),
.A2(n_1195),
.B(n_1206),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1116),
.A2(n_1096),
.B(n_1131),
.C(n_1149),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1080),
.A2(n_1125),
.B(n_1139),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_1073),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1120),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1145),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1141),
.A2(n_1203),
.B(n_1208),
.Y(n_1267)
);

AOI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1107),
.A2(n_1144),
.B(n_1138),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1209),
.A2(n_1173),
.B(n_1190),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1159),
.A2(n_1180),
.A3(n_1168),
.B(n_1104),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1135),
.A2(n_1188),
.B(n_1090),
.C(n_1142),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1207),
.A2(n_1106),
.B(n_1097),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1190),
.A2(n_1160),
.B(n_1109),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1129),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1190),
.A2(n_1168),
.B(n_1088),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1133),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1165),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1103),
.A2(n_1124),
.B1(n_1099),
.B2(n_1086),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1179),
.A2(n_1161),
.B(n_1168),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1177),
.A2(n_1135),
.B1(n_1085),
.B2(n_1114),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1094),
.A2(n_1150),
.B(n_1176),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1071),
.B(n_1081),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1140),
.A2(n_1127),
.B(n_1154),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1140),
.A2(n_1136),
.B(n_1154),
.C(n_1127),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1071),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1071),
.A2(n_1081),
.B1(n_1087),
.B2(n_1182),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_SL g1287 ( 
.A1(n_1140),
.A2(n_1127),
.B(n_1081),
.C(n_1087),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1087),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1065),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1140),
.A2(n_1191),
.A3(n_1194),
.B(n_1169),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1140),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1140),
.A2(n_1171),
.B(n_1205),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1210),
.A2(n_905),
.B(n_899),
.C(n_775),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1210),
.A2(n_905),
.B(n_899),
.C(n_775),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1210),
.A2(n_905),
.B(n_899),
.C(n_775),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_SL g1296 ( 
.A(n_1067),
.B(n_1210),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1171),
.A2(n_1205),
.B(n_1201),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1210),
.B(n_945),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1191),
.A2(n_1194),
.A3(n_1169),
.B(n_1095),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1072),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1067),
.B(n_1210),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1082),
.B(n_710),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1171),
.A2(n_1205),
.B(n_1201),
.Y(n_1303)
);

INVxp67_ASAP7_75t_L g1304 ( 
.A(n_1070),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1095),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1061),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_1067),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1146),
.B(n_963),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1067),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1210),
.A2(n_553),
.B1(n_780),
.B2(n_905),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1077),
.A2(n_951),
.B(n_877),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_SL g1312 ( 
.A1(n_1212),
.A2(n_905),
.B(n_1054),
.C(n_1062),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1210),
.A2(n_553),
.B1(n_780),
.B2(n_905),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1095),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1066),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1210),
.A2(n_780),
.B1(n_905),
.B2(n_569),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1066),
.Y(n_1317)
);

INVx4_ASAP7_75t_L g1318 ( 
.A(n_1143),
.Y(n_1318)
);

AOI221xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1115),
.A2(n_1062),
.B1(n_1123),
.B2(n_1148),
.C(n_905),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1072),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1171),
.A2(n_1205),
.B(n_1201),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1210),
.B(n_905),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1072),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1095),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1070),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1210),
.A2(n_905),
.B(n_553),
.C(n_775),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1095),
.Y(n_1327)
);

AOI31xp67_ASAP7_75t_L g1328 ( 
.A1(n_1184),
.A2(n_1197),
.A3(n_1204),
.B(n_1188),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1070),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1066),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1210),
.B(n_905),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1171),
.A2(n_1205),
.B(n_1201),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1191),
.A2(n_1194),
.A3(n_1169),
.B(n_1095),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1191),
.A2(n_1194),
.A3(n_1169),
.B(n_1095),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1061),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1095),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1071),
.Y(n_1337)
);

INVxp67_ASAP7_75t_SL g1338 ( 
.A(n_1070),
.Y(n_1338)
);

OAI22x1_ASAP7_75t_L g1339 ( 
.A1(n_1210),
.A2(n_1148),
.B1(n_1134),
.B2(n_1049),
.Y(n_1339)
);

NAND3xp33_ASAP7_75t_SL g1340 ( 
.A(n_1210),
.B(n_553),
.C(n_780),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1210),
.A2(n_553),
.B1(n_780),
.B2(n_905),
.Y(n_1341)
);

NOR2xp67_ASAP7_75t_L g1342 ( 
.A(n_1158),
.B(n_708),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1171),
.A2(n_1205),
.B(n_1201),
.Y(n_1343)
);

AND2x2_ASAP7_75t_SL g1344 ( 
.A(n_1210),
.B(n_905),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1066),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1072),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1210),
.B(n_553),
.Y(n_1347)
);

AO32x2_ASAP7_75t_L g1348 ( 
.A1(n_1077),
.A2(n_1068),
.A3(n_1049),
.B1(n_772),
.B2(n_782),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1072),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_SL g1350 ( 
.A1(n_1212),
.A2(n_905),
.B(n_1054),
.C(n_1062),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1210),
.B(n_945),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1077),
.A2(n_951),
.B(n_877),
.Y(n_1352)
);

NAND3xp33_ASAP7_75t_SL g1353 ( 
.A(n_1210),
.B(n_553),
.C(n_780),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_1070),
.Y(n_1354)
);

AO21x1_ASAP7_75t_L g1355 ( 
.A1(n_1077),
.A2(n_905),
.B(n_807),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1210),
.A2(n_905),
.B(n_899),
.C(n_775),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_SL g1357 ( 
.A1(n_1138),
.A2(n_1144),
.B(n_1131),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1210),
.A2(n_905),
.B(n_899),
.C(n_775),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1210),
.A2(n_905),
.B(n_553),
.C(n_775),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1091),
.B(n_582),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1082),
.B(n_710),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1211),
.A2(n_905),
.B(n_1095),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1171),
.A2(n_1205),
.B(n_1201),
.Y(n_1363)
);

AO31x2_ASAP7_75t_L g1364 ( 
.A1(n_1191),
.A2(n_1194),
.A3(n_1169),
.B(n_1095),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1072),
.Y(n_1365)
);

OAI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1347),
.A2(n_1341),
.B1(n_1313),
.B2(n_1310),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1298),
.A2(n_1351),
.B1(n_1331),
.B2(n_1322),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1322),
.B(n_1331),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1340),
.A2(n_1353),
.B1(n_1231),
.B2(n_1344),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1215),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1339),
.A2(n_1309),
.B1(n_1307),
.B2(n_1216),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1231),
.A2(n_1316),
.B1(n_1355),
.B2(n_1238),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1260),
.A2(n_1224),
.B1(n_1259),
.B2(n_1216),
.Y(n_1373)
);

AOI22xp5_ASAP7_75t_SL g1374 ( 
.A1(n_1260),
.A2(n_1229),
.B1(n_1289),
.B2(n_1338),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1221),
.A2(n_1232),
.B1(n_1251),
.B2(n_1296),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1264),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1251),
.A2(n_1301),
.B1(n_1218),
.B2(n_1361),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1266),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1349),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1302),
.A2(n_1330),
.B1(n_1317),
.B2(n_1345),
.Y(n_1380)
);

OAI21xp33_ASAP7_75t_L g1381 ( 
.A1(n_1326),
.A2(n_1359),
.B(n_1294),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1318),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1318),
.A2(n_1278),
.B1(n_1217),
.B2(n_1329),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_1325),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1360),
.B(n_1235),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1240),
.Y(n_1386)
);

INVx3_ASAP7_75t_L g1387 ( 
.A(n_1223),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1329),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1315),
.A2(n_1317),
.B1(n_1345),
.B2(n_1330),
.Y(n_1389)
);

BUFx10_ASAP7_75t_L g1390 ( 
.A(n_1228),
.Y(n_1390)
);

OAI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1259),
.A2(n_1365),
.B1(n_1320),
.B2(n_1323),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1226),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1315),
.A2(n_1357),
.B1(n_1243),
.B2(n_1224),
.Y(n_1393)
);

CKINVDCx11_ASAP7_75t_R g1394 ( 
.A(n_1252),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1293),
.B(n_1295),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1252),
.A2(n_1280),
.B1(n_1258),
.B2(n_1319),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1308),
.Y(n_1397)
);

BUFx8_ASAP7_75t_SL g1398 ( 
.A(n_1337),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1243),
.A2(n_1319),
.B1(n_1246),
.B2(n_1234),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1277),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1230),
.Y(n_1401)
);

INVx6_ASAP7_75t_L g1402 ( 
.A(n_1257),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1356),
.B(n_1358),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1239),
.A2(n_1245),
.B1(n_1276),
.B2(n_1265),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1337),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1271),
.A2(n_1342),
.B1(n_1304),
.B2(n_1354),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1257),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1346),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1282),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1274),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1311),
.A2(n_1352),
.B1(n_1291),
.B2(n_1249),
.Y(n_1411)
);

OAI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1223),
.A2(n_1261),
.B1(n_1233),
.B2(n_1273),
.Y(n_1412)
);

CKINVDCx11_ASAP7_75t_R g1413 ( 
.A(n_1285),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1286),
.A2(n_1281),
.B1(n_1255),
.B2(n_1237),
.Y(n_1414)
);

NAND2x1p5_ASAP7_75t_L g1415 ( 
.A(n_1283),
.B(n_1214),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1286),
.A2(n_1214),
.B1(n_1306),
.B2(n_1335),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1282),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1250),
.A2(n_1362),
.B1(n_1327),
.B2(n_1324),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1288),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1287),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1305),
.A2(n_1314),
.B1(n_1336),
.B2(n_1272),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1306),
.Y(n_1422)
);

CKINVDCx11_ASAP7_75t_R g1423 ( 
.A(n_1284),
.Y(n_1423)
);

OAI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1269),
.A2(n_1335),
.B1(n_1272),
.B2(n_1275),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1244),
.A2(n_1220),
.B1(n_1241),
.B2(n_1256),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1262),
.A2(n_1348),
.B1(n_1267),
.B2(n_1292),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1348),
.A2(n_1363),
.B1(n_1222),
.B2(n_1225),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1328),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1279),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_1312),
.Y(n_1430)
);

OAI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1268),
.A2(n_1348),
.B1(n_1350),
.B2(n_1253),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1248),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1279),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1227),
.Y(n_1434)
);

CKINVDCx6p67_ASAP7_75t_R g1435 ( 
.A(n_1254),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1247),
.A2(n_1219),
.B1(n_1364),
.B2(n_1334),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1219),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1290),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1299),
.Y(n_1439)
);

INVx6_ASAP7_75t_L g1440 ( 
.A(n_1290),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1297),
.A2(n_1303),
.B1(n_1343),
.B2(n_1332),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1321),
.A2(n_1236),
.B1(n_1242),
.B2(n_1247),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1263),
.A2(n_1299),
.B1(n_1333),
.B2(n_1334),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1299),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1333),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1334),
.B(n_1364),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1270),
.A2(n_1347),
.B1(n_1210),
.B2(n_1313),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1270),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1307),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1329),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1217),
.Y(n_1451)
);

CKINVDCx20_ASAP7_75t_R g1452 ( 
.A(n_1217),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1353),
.B2(n_1340),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1310),
.A2(n_1313),
.B1(n_1341),
.B2(n_780),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1347),
.B(n_1210),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1215),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1353),
.B2(n_1340),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1353),
.B2(n_1340),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1347),
.B(n_1210),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1300),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1347),
.B(n_1210),
.Y(n_1461)
);

AOI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_553),
.B2(n_780),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1300),
.Y(n_1463)
);

INVx6_ASAP7_75t_L g1464 ( 
.A(n_1230),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1337),
.Y(n_1465)
);

BUFx4f_ASAP7_75t_SL g1466 ( 
.A(n_1307),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1347),
.A2(n_780),
.B1(n_1210),
.B2(n_1056),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1310),
.A2(n_1313),
.B1(n_1341),
.B2(n_780),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1347),
.B(n_1210),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1329),
.Y(n_1470)
);

INVx6_ASAP7_75t_L g1471 ( 
.A(n_1230),
.Y(n_1471)
);

INVx4_ASAP7_75t_L g1472 ( 
.A(n_1217),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1310),
.A2(n_1313),
.B1(n_1341),
.B2(n_780),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1264),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1353),
.B2(n_1340),
.Y(n_1475)
);

NAND2x1p5_ASAP7_75t_L g1476 ( 
.A(n_1283),
.B(n_1189),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1313),
.B2(n_1310),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1353),
.B2(n_1340),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1353),
.B2(n_1340),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1347),
.A2(n_780),
.B1(n_1210),
.B2(n_1056),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1217),
.Y(n_1481)
);

BUFx2_ASAP7_75t_SL g1482 ( 
.A(n_1215),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1353),
.B2(n_1340),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1353),
.B2(n_1340),
.Y(n_1484)
);

BUFx8_ASAP7_75t_L g1485 ( 
.A(n_1264),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1300),
.Y(n_1486)
);

CKINVDCx11_ASAP7_75t_R g1487 ( 
.A(n_1307),
.Y(n_1487)
);

BUFx2_ASAP7_75t_SL g1488 ( 
.A(n_1215),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_1217),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1300),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1215),
.Y(n_1491)
);

CKINVDCx11_ASAP7_75t_R g1492 ( 
.A(n_1307),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1215),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1347),
.A2(n_1210),
.B1(n_1353),
.B2(n_1340),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1310),
.A2(n_1313),
.B1(n_1341),
.B2(n_780),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1329),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1432),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1462),
.A2(n_1455),
.B1(n_1461),
.B2(n_1459),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1438),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1439),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1445),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1438),
.Y(n_1502)
);

INVxp67_ASAP7_75t_R g1503 ( 
.A(n_1383),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1437),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_L g1505 ( 
.A(n_1477),
.B(n_1469),
.Y(n_1505)
);

AND2x4_ASAP7_75t_L g1506 ( 
.A(n_1444),
.B(n_1387),
.Y(n_1506)
);

OR2x6_ASAP7_75t_L g1507 ( 
.A(n_1444),
.B(n_1440),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1446),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1380),
.B(n_1389),
.Y(n_1509)
);

CKINVDCx14_ASAP7_75t_R g1510 ( 
.A(n_1449),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1367),
.B(n_1368),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_SL g1512 ( 
.A(n_1485),
.Y(n_1512)
);

AOI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1395),
.A2(n_1403),
.B(n_1411),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_SL g1514 ( 
.A(n_1485),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1380),
.B(n_1389),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1417),
.B(n_1393),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1453),
.B(n_1457),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1393),
.B(n_1372),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1433),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1392),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1454),
.A2(n_1495),
.B1(n_1468),
.B2(n_1473),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1381),
.A2(n_1478),
.B(n_1494),
.C(n_1453),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1433),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1454),
.A2(n_1473),
.B1(n_1495),
.B2(n_1468),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1442),
.A2(n_1418),
.B(n_1425),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1398),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1436),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1436),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1420),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1428),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1408),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1418),
.A2(n_1421),
.B(n_1425),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1401),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1442),
.A2(n_1421),
.B(n_1443),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1448),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1429),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1420),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1431),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1431),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1424),
.A2(n_1412),
.B(n_1447),
.Y(n_1540)
);

INVx4_ASAP7_75t_L g1541 ( 
.A(n_1420),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1443),
.A2(n_1476),
.B(n_1415),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1379),
.Y(n_1543)
);

AO31x2_ASAP7_75t_L g1544 ( 
.A1(n_1427),
.A2(n_1426),
.A3(n_1410),
.B(n_1422),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1424),
.A2(n_1412),
.B(n_1391),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1366),
.B(n_1385),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1415),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1486),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1490),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1430),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1460),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1409),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1463),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1476),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1377),
.B(n_1375),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1399),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1399),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1373),
.A2(n_1375),
.B1(n_1396),
.B2(n_1480),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1404),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1369),
.B(n_1377),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1404),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1435),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1474),
.B(n_1466),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1369),
.A2(n_1400),
.B(n_1386),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1374),
.B(n_1371),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1441),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1419),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1401),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1467),
.A2(n_1457),
.B1(n_1458),
.B2(n_1479),
.Y(n_1570)
);

AO21x2_ASAP7_75t_L g1571 ( 
.A1(n_1406),
.A2(n_1414),
.B(n_1434),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1416),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1397),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1397),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1423),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1450),
.Y(n_1576)
);

INVxp67_ASAP7_75t_SL g1577 ( 
.A(n_1378),
.Y(n_1577)
);

AOI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1458),
.A2(n_1494),
.B(n_1475),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1470),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1401),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1496),
.B(n_1483),
.Y(n_1581)
);

AOI21x1_ASAP7_75t_L g1582 ( 
.A1(n_1475),
.A2(n_1479),
.B(n_1478),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1402),
.Y(n_1583)
);

AO21x2_ASAP7_75t_L g1584 ( 
.A1(n_1483),
.A2(n_1484),
.B(n_1465),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1482),
.B(n_1488),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1376),
.Y(n_1586)
);

AO21x2_ASAP7_75t_L g1587 ( 
.A1(n_1484),
.A2(n_1465),
.B(n_1394),
.Y(n_1587)
);

INVx6_ASAP7_75t_L g1588 ( 
.A(n_1390),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1376),
.B(n_1456),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1402),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1464),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1456),
.B(n_1491),
.Y(n_1592)
);

OAI21x1_ASAP7_75t_L g1593 ( 
.A1(n_1471),
.A2(n_1382),
.B(n_1405),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1497),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1522),
.A2(n_1570),
.B(n_1505),
.Y(n_1595)
);

AOI221xp5_ASAP7_75t_L g1596 ( 
.A1(n_1517),
.A2(n_1491),
.B1(n_1493),
.B2(n_1370),
.C(n_1472),
.Y(n_1596)
);

AOI221xp5_ASAP7_75t_L g1597 ( 
.A1(n_1498),
.A2(n_1561),
.B1(n_1559),
.B2(n_1524),
.C(n_1521),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1520),
.B(n_1451),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1588),
.Y(n_1599)
);

AND2x2_ASAP7_75t_SL g1600 ( 
.A(n_1561),
.B(n_1492),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1581),
.B(n_1481),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1556),
.A2(n_1452),
.B(n_1489),
.C(n_1413),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1511),
.B(n_1466),
.Y(n_1603)
);

AO32x2_ASAP7_75t_L g1604 ( 
.A1(n_1541),
.A2(n_1390),
.A3(n_1407),
.B1(n_1487),
.B2(n_1580),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1578),
.A2(n_1582),
.B(n_1556),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_R g1606 ( 
.A(n_1563),
.B(n_1550),
.Y(n_1606)
);

AOI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1546),
.A2(n_1518),
.B1(n_1572),
.B2(n_1558),
.C(n_1557),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1503),
.A2(n_1550),
.B1(n_1566),
.B2(n_1581),
.Y(n_1608)
);

OR2x6_ASAP7_75t_L g1609 ( 
.A(n_1585),
.B(n_1593),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1576),
.B(n_1579),
.Y(n_1610)
);

NAND2xp33_ASAP7_75t_L g1611 ( 
.A(n_1529),
.B(n_1537),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1497),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1551),
.B(n_1564),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1516),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1566),
.A2(n_1571),
.B1(n_1503),
.B2(n_1587),
.Y(n_1615)
);

AO32x2_ASAP7_75t_L g1616 ( 
.A1(n_1541),
.A2(n_1580),
.A3(n_1535),
.B1(n_1528),
.B2(n_1527),
.Y(n_1616)
);

OA21x2_ASAP7_75t_L g1617 ( 
.A1(n_1534),
.A2(n_1525),
.B(n_1539),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_SL g1618 ( 
.A1(n_1510),
.A2(n_1575),
.B1(n_1589),
.B2(n_1592),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1506),
.B(n_1553),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1516),
.B(n_1543),
.Y(n_1620)
);

OAI221xp5_ASAP7_75t_L g1621 ( 
.A1(n_1578),
.A2(n_1582),
.B1(n_1515),
.B2(n_1509),
.C(n_1572),
.Y(n_1621)
);

BUFx12f_ASAP7_75t_L g1622 ( 
.A(n_1526),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1571),
.A2(n_1587),
.B1(n_1584),
.B2(n_1540),
.Y(n_1623)
);

AOI221xp5_ASAP7_75t_L g1624 ( 
.A1(n_1557),
.A2(n_1562),
.B1(n_1560),
.B2(n_1538),
.C(n_1528),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1586),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1509),
.B(n_1515),
.Y(n_1626)
);

BUFx4f_ASAP7_75t_SL g1627 ( 
.A(n_1526),
.Y(n_1627)
);

AO32x2_ASAP7_75t_L g1628 ( 
.A1(n_1541),
.A2(n_1527),
.A3(n_1544),
.B1(n_1536),
.B2(n_1508),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1506),
.B(n_1568),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1587),
.B(n_1592),
.Y(n_1630)
);

INVx4_ASAP7_75t_L g1631 ( 
.A(n_1585),
.Y(n_1631)
);

BUFx3_ASAP7_75t_L g1632 ( 
.A(n_1588),
.Y(n_1632)
);

AO32x2_ASAP7_75t_L g1633 ( 
.A1(n_1544),
.A2(n_1536),
.A3(n_1508),
.B1(n_1499),
.B2(n_1502),
.Y(n_1633)
);

OAI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1513),
.A2(n_1565),
.B(n_1585),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1563),
.A2(n_1575),
.B(n_1560),
.C(n_1562),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1563),
.B(n_1590),
.Y(n_1636)
);

A2O1A1Ixp33_ASAP7_75t_L g1637 ( 
.A1(n_1567),
.A2(n_1529),
.B(n_1537),
.C(n_1573),
.Y(n_1637)
);

O2A1O1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1540),
.A2(n_1545),
.B(n_1584),
.C(n_1567),
.Y(n_1638)
);

AOI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1584),
.A2(n_1540),
.B1(n_1545),
.B2(n_1529),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1500),
.Y(n_1640)
);

A2O1A1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1529),
.A2(n_1537),
.B(n_1573),
.C(n_1542),
.Y(n_1641)
);

AO21x2_ASAP7_75t_L g1642 ( 
.A1(n_1519),
.A2(n_1523),
.B(n_1530),
.Y(n_1642)
);

NAND4xp25_ASAP7_75t_L g1643 ( 
.A(n_1548),
.B(n_1549),
.C(n_1554),
.D(n_1552),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_SL g1644 ( 
.A1(n_1574),
.A2(n_1555),
.B(n_1547),
.C(n_1591),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1617),
.B(n_1544),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1617),
.B(n_1544),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1614),
.B(n_1544),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1633),
.B(n_1532),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1594),
.Y(n_1649)
);

BUFx4f_ASAP7_75t_SL g1650 ( 
.A(n_1622),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1609),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1612),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1620),
.B(n_1519),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_SL g1654 ( 
.A1(n_1595),
.A2(n_1537),
.B(n_1512),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1642),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1633),
.B(n_1532),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1640),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1616),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1628),
.B(n_1532),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1628),
.B(n_1500),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1628),
.B(n_1501),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1626),
.B(n_1501),
.Y(n_1662)
);

NOR2x1_ASAP7_75t_SL g1663 ( 
.A(n_1609),
.B(n_1507),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1616),
.B(n_1542),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1639),
.B(n_1504),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1629),
.B(n_1547),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1630),
.B(n_1623),
.Y(n_1667)
);

INVxp67_ASAP7_75t_SL g1668 ( 
.A(n_1638),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1624),
.B(n_1531),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1634),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1668),
.B(n_1605),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1664),
.B(n_1641),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1663),
.B(n_1631),
.Y(n_1673)
);

AND4x1_ASAP7_75t_L g1674 ( 
.A(n_1650),
.B(n_1615),
.C(n_1597),
.D(n_1635),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1668),
.A2(n_1607),
.B1(n_1621),
.B2(n_1600),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1657),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1660),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1655),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1660),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1658),
.B(n_1610),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1658),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1660),
.B(n_1661),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1662),
.B(n_1653),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1660),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1651),
.Y(n_1685)
);

INVx6_ASAP7_75t_L g1686 ( 
.A(n_1666),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1661),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1647),
.B(n_1645),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1661),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1661),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1667),
.B(n_1629),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1647),
.B(n_1625),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1647),
.B(n_1643),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1649),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1667),
.B(n_1619),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1659),
.A2(n_1611),
.B(n_1644),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1667),
.B(n_1619),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_1667),
.Y(n_1698)
);

AOI32xp33_ASAP7_75t_L g1699 ( 
.A1(n_1669),
.A2(n_1608),
.A3(n_1596),
.B1(n_1613),
.B2(n_1603),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1652),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1681),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1676),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1682),
.B(n_1670),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1674),
.B(n_1670),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1676),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1682),
.B(n_1670),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1682),
.B(n_1648),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1671),
.B(n_1665),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1681),
.B(n_1646),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1671),
.B(n_1665),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1677),
.B(n_1679),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1686),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1677),
.B(n_1648),
.Y(n_1713)
);

OR2x6_ASAP7_75t_L g1714 ( 
.A(n_1673),
.B(n_1696),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1694),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1677),
.B(n_1679),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1685),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1679),
.B(n_1687),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1679),
.B(n_1648),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1694),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1674),
.B(n_1654),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1685),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1687),
.B(n_1656),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1687),
.B(n_1656),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1687),
.B(n_1656),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_1678),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1685),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1690),
.B(n_1645),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1690),
.B(n_1684),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1700),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1690),
.B(n_1656),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1694),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1698),
.B(n_1665),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1708),
.B(n_1693),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1701),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1704),
.A2(n_1674),
.B(n_1675),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1721),
.A2(n_1675),
.B1(n_1654),
.B2(n_1699),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1717),
.Y(n_1738)
);

AOI32xp33_ASAP7_75t_L g1739 ( 
.A1(n_1721),
.A2(n_1672),
.A3(n_1673),
.B1(n_1697),
.B2(n_1695),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1717),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1714),
.B(n_1672),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1708),
.B(n_1693),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1714),
.B(n_1672),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1701),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1714),
.B(n_1684),
.Y(n_1745)
);

NAND4xp25_ASAP7_75t_SL g1746 ( 
.A(n_1704),
.B(n_1699),
.C(n_1696),
.D(n_1602),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1717),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1717),
.B(n_1673),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1714),
.B(n_1689),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1720),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1720),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1710),
.B(n_1693),
.Y(n_1752)
);

OR2x6_ASAP7_75t_L g1753 ( 
.A(n_1717),
.B(n_1654),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1715),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1715),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1717),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1714),
.B(n_1689),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1715),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1710),
.B(n_1698),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1733),
.B(n_1683),
.Y(n_1760)
);

NAND2x1_ASAP7_75t_L g1761 ( 
.A(n_1714),
.B(n_1686),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1730),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1722),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1733),
.B(n_1683),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1722),
.B(n_1680),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1730),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1727),
.B(n_1680),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1730),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1714),
.B(n_1691),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1732),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1714),
.B(n_1691),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1703),
.B(n_1691),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1732),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1727),
.B(n_1680),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1703),
.B(n_1688),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1703),
.B(n_1706),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1732),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1717),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1738),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1738),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1736),
.B(n_1706),
.Y(n_1781)
);

OAI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1746),
.A2(n_1726),
.B(n_1618),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1744),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1740),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1737),
.B(n_1650),
.Y(n_1785)
);

INVxp67_ASAP7_75t_L g1786 ( 
.A(n_1763),
.Y(n_1786)
);

NAND4xp75_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1706),
.C(n_1514),
.D(n_1712),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1740),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1753),
.B(n_1717),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1744),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1747),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1750),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1735),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1772),
.B(n_1734),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1761),
.B(n_1717),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1753),
.B(n_1707),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1742),
.B(n_1688),
.Y(n_1797)
);

NAND2xp33_ASAP7_75t_L g1798 ( 
.A(n_1739),
.B(n_1699),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1772),
.B(n_1695),
.Y(n_1799)
);

OR2x6_ASAP7_75t_L g1800 ( 
.A(n_1753),
.B(n_1712),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1750),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1742),
.B(n_1688),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1751),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1751),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1765),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1753),
.B(n_1707),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1752),
.B(n_1726),
.Y(n_1807)
);

OR2x6_ASAP7_75t_L g1808 ( 
.A(n_1761),
.B(n_1712),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1776),
.B(n_1748),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1741),
.B(n_1707),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1754),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1743),
.B(n_1712),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1754),
.Y(n_1813)
);

NAND2x1_ASAP7_75t_L g1814 ( 
.A(n_1748),
.B(n_1743),
.Y(n_1814)
);

OR2x6_ASAP7_75t_L g1815 ( 
.A(n_1747),
.B(n_1631),
.Y(n_1815)
);

NAND2xp33_ASAP7_75t_SL g1816 ( 
.A(n_1782),
.B(n_1606),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1786),
.B(n_1776),
.Y(n_1817)
);

OAI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1781),
.A2(n_1759),
.B1(n_1775),
.B2(n_1765),
.Y(n_1818)
);

A2O1A1Ixp33_ASAP7_75t_L g1819 ( 
.A1(n_1798),
.A2(n_1749),
.B(n_1757),
.C(n_1745),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1805),
.B(n_1760),
.Y(n_1820)
);

NAND3xp33_ASAP7_75t_L g1821 ( 
.A(n_1798),
.B(n_1756),
.C(n_1767),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1792),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1785),
.Y(n_1823)
);

AND2x2_ASAP7_75t_SL g1824 ( 
.A(n_1789),
.B(n_1601),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1794),
.B(n_1759),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1814),
.A2(n_1774),
.B(n_1778),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1809),
.B(n_1812),
.Y(n_1827)
);

OAI21xp33_ASAP7_75t_L g1828 ( 
.A1(n_1793),
.A2(n_1749),
.B(n_1745),
.Y(n_1828)
);

AOI322xp5_ASAP7_75t_L g1829 ( 
.A1(n_1796),
.A2(n_1731),
.A3(n_1719),
.B1(n_1725),
.B2(n_1713),
.C1(n_1724),
.C2(n_1723),
.Y(n_1829)
);

OAI21xp33_ASAP7_75t_L g1830 ( 
.A1(n_1796),
.A2(n_1757),
.B(n_1769),
.Y(n_1830)
);

OA21x2_ASAP7_75t_L g1831 ( 
.A1(n_1787),
.A2(n_1756),
.B(n_1755),
.Y(n_1831)
);

AO22x1_ASAP7_75t_L g1832 ( 
.A1(n_1789),
.A2(n_1809),
.B1(n_1806),
.B2(n_1790),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1792),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1783),
.B(n_1764),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1806),
.B(n_1769),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1807),
.B(n_1775),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1787),
.A2(n_1748),
.B1(n_1771),
.B2(n_1673),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1801),
.B(n_1771),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1813),
.Y(n_1839)
);

O2A1O1Ixp33_ASAP7_75t_L g1840 ( 
.A1(n_1800),
.A2(n_1678),
.B(n_1637),
.C(n_1709),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1813),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1821),
.A2(n_1814),
.B1(n_1800),
.B2(n_1809),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1821),
.A2(n_1800),
.B1(n_1795),
.B2(n_1799),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1839),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1841),
.Y(n_1845)
);

OAI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1816),
.A2(n_1800),
.B1(n_1807),
.B2(n_1795),
.C(n_1808),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1822),
.Y(n_1847)
);

AOI32xp33_ASAP7_75t_L g1848 ( 
.A1(n_1818),
.A2(n_1827),
.A3(n_1817),
.B1(n_1830),
.B2(n_1828),
.Y(n_1848)
);

OAI222xp33_ASAP7_75t_L g1849 ( 
.A1(n_1840),
.A2(n_1826),
.B1(n_1817),
.B2(n_1820),
.C1(n_1836),
.C2(n_1834),
.Y(n_1849)
);

AOI21xp33_ASAP7_75t_SL g1850 ( 
.A1(n_1831),
.A2(n_1795),
.B(n_1808),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1824),
.B(n_1812),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_R g1852 ( 
.A(n_1823),
.B(n_1627),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1833),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1831),
.B(n_1810),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1832),
.Y(n_1855)
);

AOI32xp33_ASAP7_75t_L g1856 ( 
.A1(n_1835),
.A2(n_1810),
.A3(n_1803),
.B1(n_1804),
.B2(n_1797),
.Y(n_1856)
);

OAI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1837),
.A2(n_1808),
.B1(n_1815),
.B2(n_1797),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1819),
.B(n_1802),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1838),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_SL g1860 ( 
.A1(n_1825),
.A2(n_1673),
.B(n_1802),
.Y(n_1860)
);

NAND2x1_ASAP7_75t_SL g1861 ( 
.A(n_1829),
.B(n_1779),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1858),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1844),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1855),
.B(n_1779),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1848),
.B(n_1780),
.Y(n_1865)
);

XNOR2x1_ASAP7_75t_L g1866 ( 
.A(n_1842),
.B(n_1598),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1858),
.B(n_1780),
.Y(n_1867)
);

OAI21xp33_ASAP7_75t_L g1868 ( 
.A1(n_1861),
.A2(n_1811),
.B(n_1808),
.Y(n_1868)
);

AO22x1_ASAP7_75t_L g1869 ( 
.A1(n_1854),
.A2(n_1791),
.B1(n_1788),
.B2(n_1784),
.Y(n_1869)
);

AOI322xp5_ASAP7_75t_L g1870 ( 
.A1(n_1857),
.A2(n_1719),
.A3(n_1725),
.B1(n_1724),
.B2(n_1723),
.C1(n_1731),
.C2(n_1713),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1845),
.Y(n_1871)
);

AOI32xp33_ASAP7_75t_L g1872 ( 
.A1(n_1843),
.A2(n_1857),
.A3(n_1851),
.B1(n_1846),
.B2(n_1859),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1864),
.Y(n_1873)
);

AOI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1868),
.A2(n_1849),
.B1(n_1850),
.B2(n_1856),
.C(n_1847),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1867),
.Y(n_1875)
);

NAND4xp75_ASAP7_75t_L g1876 ( 
.A(n_1865),
.B(n_1853),
.C(n_1849),
.D(n_1784),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1862),
.B(n_1852),
.Y(n_1877)
);

NOR4xp25_ASAP7_75t_SL g1878 ( 
.A(n_1863),
.B(n_1860),
.C(n_1871),
.D(n_1869),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1872),
.B(n_1788),
.Y(n_1879)
);

NAND5xp2_ASAP7_75t_L g1880 ( 
.A(n_1870),
.B(n_1636),
.C(n_1604),
.D(n_1768),
.E(n_1773),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1866),
.B(n_1815),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1862),
.B(n_1791),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1876),
.A2(n_1815),
.B1(n_1673),
.B2(n_1598),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1879),
.B(n_1815),
.Y(n_1884)
);

AOI21xp33_ASAP7_75t_L g1885 ( 
.A1(n_1877),
.A2(n_1766),
.B(n_1755),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1875),
.Y(n_1886)
);

INVxp67_ASAP7_75t_L g1887 ( 
.A(n_1882),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1886),
.Y(n_1888)
);

NAND5xp2_ASAP7_75t_L g1889 ( 
.A(n_1887),
.B(n_1874),
.C(n_1881),
.D(n_1873),
.E(n_1878),
.Y(n_1889)
);

AOI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1885),
.A2(n_1880),
.B1(n_1766),
.B2(n_1768),
.C(n_1770),
.Y(n_1890)
);

NAND3xp33_ASAP7_75t_L g1891 ( 
.A(n_1884),
.B(n_1773),
.C(n_1770),
.Y(n_1891)
);

OAI22xp5_ASAP7_75t_L g1892 ( 
.A1(n_1883),
.A2(n_1709),
.B1(n_1777),
.B2(n_1758),
.Y(n_1892)
);

OAI211xp5_ASAP7_75t_SL g1893 ( 
.A1(n_1887),
.A2(n_1762),
.B(n_1709),
.C(n_1692),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1888),
.B(n_1729),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1891),
.Y(n_1895)
);

NAND4xp75_ASAP7_75t_L g1896 ( 
.A(n_1890),
.B(n_1889),
.C(n_1892),
.D(n_1893),
.Y(n_1896)
);

XOR2xp5_ASAP7_75t_L g1897 ( 
.A(n_1888),
.B(n_1663),
.Y(n_1897)
);

NOR2x1_ASAP7_75t_L g1898 ( 
.A(n_1889),
.B(n_1711),
.Y(n_1898)
);

AOI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1898),
.A2(n_1588),
.B1(n_1729),
.B2(n_1599),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1894),
.Y(n_1900)
);

NAND3xp33_ASAP7_75t_L g1901 ( 
.A(n_1895),
.B(n_1537),
.C(n_1702),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1900),
.A2(n_1897),
.B1(n_1899),
.B2(n_1901),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1902),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1903),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1903),
.B(n_1896),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1904),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1905),
.A2(n_1588),
.B1(n_1711),
.B2(n_1728),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1906),
.A2(n_1729),
.B1(n_1718),
.B2(n_1716),
.Y(n_1908)
);

AOI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1907),
.B(n_1705),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1909),
.A2(n_1705),
.B(n_1702),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1910),
.Y(n_1911)
);

OAI221xp5_ASAP7_75t_L g1912 ( 
.A1(n_1911),
.A2(n_1632),
.B1(n_1583),
.B2(n_1569),
.C(n_1533),
.Y(n_1912)
);

AOI211xp5_ASAP7_75t_L g1913 ( 
.A1(n_1912),
.A2(n_1583),
.B(n_1569),
.C(n_1533),
.Y(n_1913)
);


endmodule