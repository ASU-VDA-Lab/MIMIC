module fake_netlist_6_313_n_2129 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2129);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2129;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1832;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2017;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_61),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_87),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_152),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_134),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_47),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_127),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_143),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_58),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_118),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_4),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_30),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_98),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_81),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_147),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_158),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_194),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_189),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_23),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_24),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_86),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_110),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_64),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_156),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_49),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_106),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_103),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_29),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_175),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_79),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_56),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_95),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_195),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_58),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_61),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_157),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_17),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_208),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_150),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_65),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_159),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_15),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_174),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_146),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_13),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_115),
.Y(n_268)
);

BUFx8_ASAP7_75t_SL g269 ( 
.A(n_130),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_188),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_140),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_2),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_203),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_37),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_10),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_52),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_26),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_99),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_56),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_101),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_199),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_144),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_64),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_13),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_190),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_114),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_31),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_49),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_40),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_54),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_122),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_100),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_186),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_30),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_162),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_88),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_17),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_39),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_41),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_85),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_173),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_4),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_126),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_183),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_39),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_18),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_6),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_2),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_102),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_44),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_70),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_117),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_10),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_167),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_200),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_155),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_42),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_1),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_182),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_67),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_78),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_196),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_192),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_70),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_170),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_63),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_154),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_46),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_94),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_84),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_133),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_67),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_73),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_38),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_141),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_109),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_191),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_27),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_43),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_40),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_45),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_35),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_57),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_38),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_53),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_128),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_136),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_107),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_169),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_46),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_33),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_149),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_26),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_18),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_210),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_29),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_151),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_112),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_41),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_15),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_137),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_97),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_23),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_33),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_37),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_43),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_50),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_8),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_76),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_179),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_59),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_7),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_5),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_165),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_131),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_16),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_181),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_19),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_21),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_52),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_105),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_65),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_89),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_36),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_5),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_7),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_75),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_123),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_116),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_82),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_34),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_20),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_83),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_36),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_60),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_111),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_68),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_121),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_205),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_92),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_168),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_129),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_163),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_180),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_93),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_96),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_45),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_145),
.Y(n_409)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_80),
.Y(n_410)
);

BUFx5_ASAP7_75t_L g411 ( 
.A(n_197),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_44),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_204),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_63),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_209),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_42),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_90),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_218),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_218),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_220),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_245),
.B(n_0),
.Y(n_421)
);

INVxp33_ASAP7_75t_L g422 ( 
.A(n_298),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_218),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_269),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_261),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_233),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_295),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_216),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_218),
.Y(n_429)
);

INVxp33_ASAP7_75t_SL g430 ( 
.A(n_212),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_266),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_218),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_265),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_275),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_275),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_297),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_275),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_275),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_280),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_281),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_270),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_303),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_282),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_292),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_295),
.B(n_0),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_302),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_356),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_362),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_305),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_219),
.B(n_1),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_275),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_316),
.Y(n_454)
);

BUFx2_ASAP7_75t_SL g455 ( 
.A(n_271),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_350),
.B(n_3),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_371),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_290),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_324),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_328),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_320),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_290),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_290),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_290),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_411),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_290),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_411),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_404),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_410),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_223),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_330),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_340),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_340),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_340),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_340),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_340),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_351),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_295),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_331),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_351),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_351),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_351),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_332),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_351),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_337),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_392),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_347),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_277),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_212),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_L g490 ( 
.A(n_219),
.B(n_3),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_356),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_348),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_349),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_353),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_359),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_417),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_277),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_219),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_262),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_411),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_274),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_276),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_307),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_R g504 ( 
.A(n_217),
.B(n_221),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_279),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_283),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_307),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_411),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_217),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_314),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_398),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_284),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_285),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_314),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_321),
.B(n_6),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_346),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_291),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_293),
.B(n_213),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_293),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_221),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_299),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_312),
.Y(n_522)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_398),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_418),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_420),
.B(n_398),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_418),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_490),
.B(n_293),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_434),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_321),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_498),
.B(n_226),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_419),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_441),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_515),
.B(n_213),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_441),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_465),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_423),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_429),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_490),
.B(n_238),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_465),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_429),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_432),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_515),
.B(n_238),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_432),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_435),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_435),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_427),
.B(n_447),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_519),
.B(n_286),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_491),
.B(n_226),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_427),
.B(n_286),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_467),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_436),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_425),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_421),
.B(n_223),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_467),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_436),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_447),
.B(n_310),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_500),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_438),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_439),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_439),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_453),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_453),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_458),
.B(n_230),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_500),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_458),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_462),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_500),
.Y(n_575)
);

BUFx8_ASAP7_75t_L g576 ( 
.A(n_444),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_462),
.B(n_310),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_508),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_463),
.B(n_464),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_489),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_508),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_463),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_449),
.B(n_336),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_508),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_464),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_466),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_466),
.B(n_336),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_472),
.B(n_338),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_473),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_473),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_474),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_474),
.B(n_230),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_449),
.B(n_338),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_475),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_475),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_422),
.A2(n_308),
.B1(n_300),
.B2(n_240),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_476),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_476),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_477),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_449),
.B(n_477),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_480),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_486),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_480),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_481),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_481),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_482),
.B(n_231),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_484),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_484),
.B(n_214),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_518),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_529),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_L g613 ( 
.A(n_611),
.B(n_452),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_553),
.B(n_426),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_529),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_525),
.A2(n_576),
.B1(n_470),
.B2(n_523),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_579),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_603),
.B(n_420),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_579),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_553),
.B(n_433),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_559),
.B(n_431),
.Y(n_621)
);

AND2x4_ASAP7_75t_L g622 ( 
.A(n_601),
.B(n_488),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_611),
.B(n_440),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_579),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_579),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_601),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_538),
.A2(n_548),
.B1(n_553),
.B2(n_611),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_583),
.B(n_488),
.Y(n_628)
);

AND2x2_ASAP7_75t_SL g629 ( 
.A(n_563),
.B(n_456),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_601),
.Y(n_630)
);

AND2x6_ASAP7_75t_L g631 ( 
.A(n_527),
.B(n_229),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_579),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_559),
.A2(n_525),
.B1(n_306),
.B2(n_334),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_533),
.B(n_442),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_552),
.B(n_497),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_524),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_565),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_580),
.A2(n_343),
.B1(n_255),
.B2(n_222),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_565),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_524),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_524),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_611),
.B(n_445),
.Y(n_642)
);

CKINVDCx14_ASAP7_75t_R g643 ( 
.A(n_558),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_524),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_554),
.B(n_470),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_533),
.B(n_446),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_554),
.B(n_448),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_529),
.Y(n_648)
);

INVx5_ASAP7_75t_L g649 ( 
.A(n_529),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_529),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_600),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_611),
.B(n_538),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_532),
.B(n_455),
.Y(n_653)
);

BUFx4f_ASAP7_75t_L g654 ( 
.A(n_611),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_565),
.Y(n_655)
);

INVxp33_ASAP7_75t_L g656 ( 
.A(n_603),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_573),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_573),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_529),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_573),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_597),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_600),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_600),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_538),
.A2(n_444),
.B1(n_357),
.B2(n_365),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_548),
.A2(n_357),
.B1(n_365),
.B2(n_346),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_600),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_532),
.B(n_451),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_611),
.B(n_548),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_528),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_552),
.B(n_454),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_563),
.A2(n_387),
.B1(n_430),
.B2(n_224),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_571),
.B(n_229),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_528),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_563),
.A2(n_387),
.B1(n_251),
.B2(n_264),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_563),
.A2(n_258),
.B1(n_272),
.B2(n_267),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_576),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_576),
.B(n_437),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_576),
.Y(n_678)
);

OR2x6_ASAP7_75t_L g679 ( 
.A(n_543),
.B(n_455),
.Y(n_679)
);

BUFx10_ASAP7_75t_L g680 ( 
.A(n_563),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_528),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_610),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_552),
.B(n_459),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_583),
.B(n_594),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_528),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_530),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_530),
.Y(n_687)
);

CKINVDCx6p67_ASAP7_75t_R g688 ( 
.A(n_580),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_552),
.B(n_497),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_530),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_526),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_552),
.B(n_460),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_529),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_583),
.B(n_503),
.Y(n_694)
);

AND2x6_ASAP7_75t_L g695 ( 
.A(n_527),
.B(n_229),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_526),
.Y(n_696)
);

INVxp33_ASAP7_75t_L g697 ( 
.A(n_597),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_594),
.B(n_471),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_530),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_610),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_527),
.A2(n_222),
.B1(n_235),
.B2(n_225),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_529),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_531),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_543),
.A2(n_325),
.B1(n_327),
.B2(n_319),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_576),
.B(n_437),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_571),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_539),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_536),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_531),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_539),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_L g711 ( 
.A(n_593),
.B(n_501),
.C(n_499),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_610),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_527),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_608),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_536),
.Y(n_715)
);

BUFx4f_ASAP7_75t_L g716 ( 
.A(n_543),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_555),
.B(n_503),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_534),
.Y(n_718)
);

OR2x6_ASAP7_75t_L g719 ( 
.A(n_543),
.B(n_288),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_608),
.B(n_479),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_534),
.B(n_483),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_539),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_537),
.B(n_492),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_537),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_610),
.B(n_457),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_536),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_541),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_541),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_542),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_543),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_542),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_543),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_536),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_536),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_545),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_539),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_610),
.B(n_457),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_555),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_540),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_555),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_540),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_545),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_546),
.B(n_493),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_540),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_543),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_540),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_536),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_546),
.B(n_494),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_536),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_536),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_544),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_549),
.B(n_495),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_544),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_L g754 ( 
.A(n_564),
.B(n_229),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_549),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_564),
.B(n_229),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_544),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_544),
.Y(n_758)
);

AO22x2_ASAP7_75t_L g759 ( 
.A1(n_555),
.A2(n_309),
.B1(n_311),
.B2(n_289),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_564),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_716),
.B(n_273),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_738),
.Y(n_762)
);

BUFx5_ASAP7_75t_L g763 ( 
.A(n_680),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_628),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_716),
.B(n_680),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_627),
.B(n_502),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_622),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_714),
.B(n_505),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_634),
.B(n_506),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_620),
.B(n_614),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_629),
.A2(n_329),
.B1(n_333),
.B2(n_318),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_646),
.B(n_512),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_691),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_626),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_684),
.B(n_513),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_626),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_630),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_684),
.B(n_507),
.Y(n_778)
);

INVx8_ASAP7_75t_L g779 ( 
.A(n_653),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_652),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_622),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_630),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_620),
.B(n_517),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_647),
.B(n_521),
.Y(n_784)
);

AOI221xp5_ASAP7_75t_L g785 ( 
.A1(n_697),
.A2(n_408),
.B1(n_246),
.B2(n_243),
.C(n_254),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_629),
.A2(n_341),
.B1(n_342),
.B2(n_339),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_716),
.B(n_273),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_L g788 ( 
.A(n_706),
.B(n_411),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_L g789 ( 
.A(n_633),
.B(n_522),
.C(n_511),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_717),
.Y(n_790)
);

BUFx4_ASAP7_75t_L g791 ( 
.A(n_643),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_720),
.B(n_450),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_682),
.Y(n_793)
);

BUFx6f_ASAP7_75t_SL g794 ( 
.A(n_653),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_717),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_668),
.B(n_564),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_682),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_691),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_740),
.B(n_564),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_680),
.B(n_273),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_629),
.B(n_667),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_622),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_621),
.B(n_424),
.C(n_315),
.Y(n_803)
);

AND2x6_ASAP7_75t_SL g804 ( 
.A(n_653),
.B(n_344),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_614),
.B(n_428),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_669),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_654),
.B(n_713),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_635),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_696),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_623),
.B(n_572),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_618),
.B(n_225),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_642),
.B(n_572),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_721),
.B(n_572),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_700),
.Y(n_814)
);

AO22x2_ASAP7_75t_L g815 ( 
.A1(n_661),
.A2(n_705),
.B1(n_677),
.B2(n_732),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_696),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_635),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_656),
.B(n_443),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_654),
.B(n_273),
.Y(n_819)
);

BUFx6f_ASAP7_75t_SL g820 ( 
.A(n_653),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_723),
.B(n_572),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_700),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_712),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_712),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_703),
.Y(n_825)
);

OAI22xp33_ASAP7_75t_L g826 ( 
.A1(n_633),
.A2(n_360),
.B1(n_372),
.B2(n_354),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_671),
.B(n_487),
.C(n_485),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_743),
.B(n_575),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_698),
.B(n_575),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_617),
.B(n_575),
.Y(n_830)
);

NAND3xp33_ASAP7_75t_L g831 ( 
.A(n_664),
.B(n_496),
.C(n_509),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_654),
.B(n_273),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_617),
.B(n_575),
.Y(n_833)
);

INVx8_ASAP7_75t_L g834 ( 
.A(n_679),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_613),
.A2(n_373),
.B(n_379),
.C(n_377),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_L g836 ( 
.A(n_730),
.B(n_411),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_635),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_703),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_628),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_619),
.B(n_575),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_732),
.B(n_296),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_619),
.B(n_575),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_689),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_645),
.B(n_711),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_689),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_624),
.B(n_575),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_730),
.A2(n_520),
.B1(n_468),
.B2(n_461),
.Y(n_847)
);

BUFx6f_ASAP7_75t_SL g848 ( 
.A(n_679),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_689),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_624),
.A2(n_469),
.B1(n_384),
.B2(n_232),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_709),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_694),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_670),
.B(n_231),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_709),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_718),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_688),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_759),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_718),
.Y(n_858)
);

AND2x6_ASAP7_75t_L g859 ( 
.A(n_625),
.B(n_296),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_632),
.B(n_296),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_724),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_632),
.B(n_296),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_636),
.B(n_578),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_636),
.B(n_578),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_676),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_694),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_724),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_701),
.A2(n_388),
.B(n_386),
.C(n_227),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_SL g869 ( 
.A(n_678),
.B(n_676),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_727),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_640),
.B(n_578),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_683),
.B(n_692),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_725),
.B(n_507),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_640),
.B(n_578),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_688),
.B(n_504),
.Y(n_875)
);

BUFx5_ASAP7_75t_L g876 ( 
.A(n_631),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_748),
.B(n_234),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_641),
.B(n_644),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_727),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_759),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_641),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_618),
.B(n_550),
.Y(n_882)
);

INVxp33_ASAP7_75t_L g883 ( 
.A(n_638),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_644),
.B(n_651),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_728),
.Y(n_885)
);

NOR3xp33_ASAP7_75t_L g886 ( 
.A(n_616),
.B(n_345),
.C(n_335),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_728),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_651),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_662),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_752),
.B(n_234),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_679),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_663),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_638),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_663),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_704),
.B(n_244),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_729),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_SL g897 ( 
.A(n_678),
.B(n_223),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_759),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_701),
.B(n_510),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_666),
.B(n_729),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_745),
.B(n_296),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_613),
.A2(n_737),
.B1(n_679),
.B2(n_719),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_731),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_731),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_745),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_735),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_719),
.A2(n_382),
.B1(n_375),
.B2(n_370),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_735),
.B(n_578),
.Y(n_908)
);

NOR3xp33_ASAP7_75t_L g909 ( 
.A(n_742),
.B(n_355),
.C(n_352),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_665),
.B(n_510),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_742),
.B(n_755),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_755),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_637),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_745),
.B(n_304),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_726),
.B(n_577),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_759),
.Y(n_916)
);

INVx5_ASAP7_75t_L g917 ( 
.A(n_631),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_650),
.B(n_304),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_637),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_773),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_801),
.A2(n_771),
.B1(n_786),
.B2(n_902),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_780),
.A2(n_715),
.B(n_693),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_770),
.B(n_650),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_872),
.B(n_760),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_773),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_771),
.A2(n_786),
.B1(n_880),
.B2(n_857),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_796),
.A2(n_715),
.B(n_693),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_793),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_810),
.A2(n_812),
.B(n_799),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_L g930 ( 
.A(n_827),
.B(n_249),
.C(n_244),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_793),
.B(n_650),
.Y(n_931)
);

OAI22xp5_ASAP7_75t_L g932 ( 
.A1(n_766),
.A2(n_719),
.B1(n_674),
.B2(n_675),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_872),
.B(n_615),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_863),
.A2(n_659),
.B(n_615),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_895),
.A2(n_672),
.B(n_228),
.C(n_236),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_915),
.A2(n_747),
.B(n_702),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_779),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_793),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_829),
.A2(n_702),
.B(n_650),
.Y(n_939)
);

OAI21xp5_ASAP7_75t_L g940 ( 
.A1(n_830),
.A2(n_760),
.B(n_659),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_783),
.B(n_719),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_793),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_798),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_798),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_813),
.A2(n_702),
.B(n_650),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_844),
.A2(n_672),
.B1(n_695),
.B2(n_631),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_809),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_821),
.A2(n_750),
.B(n_708),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_809),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_833),
.A2(n_760),
.B(n_659),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_814),
.B(n_708),
.Y(n_951)
);

OAI21xp5_ASAP7_75t_L g952 ( 
.A1(n_840),
.A2(n_733),
.B(n_615),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_828),
.A2(n_750),
.B(n_708),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_842),
.A2(n_734),
.B(n_733),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_895),
.A2(n_239),
.B(n_241),
.C(n_215),
.Y(n_955)
);

OAI21xp33_ASAP7_75t_L g956 ( 
.A1(n_768),
.A2(n_237),
.B(n_235),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_769),
.B(n_772),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_814),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_762),
.B(n_733),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_846),
.A2(n_749),
.B(n_734),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_768),
.B(n_514),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_784),
.B(n_673),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_826),
.A2(n_756),
.B(n_754),
.C(n_655),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_816),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_816),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_826),
.A2(n_756),
.B(n_754),
.C(n_655),
.Y(n_966)
);

BUFx4f_ASAP7_75t_L g967 ( 
.A(n_779),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_807),
.A2(n_648),
.B(n_612),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_825),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_868),
.A2(n_657),
.B(n_658),
.C(n_639),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_883),
.B(n_361),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_805),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_775),
.B(n_364),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_814),
.B(n_681),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_814),
.B(n_681),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_818),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_774),
.B(n_685),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_776),
.B(n_685),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_823),
.Y(n_979)
);

INVxp67_ASAP7_75t_L g980 ( 
.A(n_882),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_822),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_825),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_777),
.B(n_686),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_807),
.A2(n_648),
.B(n_612),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_893),
.B(n_237),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_838),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_856),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_779),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_L g989 ( 
.A(n_831),
.B(n_250),
.C(n_249),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_765),
.A2(n_648),
.B(n_612),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_823),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_822),
.Y(n_992)
);

AOI22x1_ASAP7_75t_L g993 ( 
.A1(n_838),
.A2(n_639),
.B1(n_657),
.B2(n_658),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_857),
.A2(n_631),
.B1(n_695),
.B2(n_400),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_765),
.A2(n_648),
.B(n_612),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_767),
.A2(n_313),
.B1(n_301),
.B2(n_294),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_864),
.A2(n_687),
.B(n_686),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_908),
.A2(n_690),
.B(n_687),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_782),
.B(n_690),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_851),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_824),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_854),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_SL g1003 ( 
.A(n_865),
.B(n_250),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_844),
.A2(n_376),
.B(n_247),
.C(n_248),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_763),
.B(n_905),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_854),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_877),
.B(n_699),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_855),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_871),
.A2(n_758),
.B(n_710),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_877),
.B(n_707),
.Y(n_1010)
);

AO21x1_ASAP7_75t_L g1011 ( 
.A1(n_761),
.A2(n_252),
.B(n_242),
.Y(n_1011)
);

O2A1O1Ixp5_ASAP7_75t_L g1012 ( 
.A1(n_819),
.A2(n_832),
.B(n_761),
.C(n_787),
.Y(n_1012)
);

NAND2x1_ASAP7_75t_L g1013 ( 
.A(n_797),
.B(n_631),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_868),
.A2(n_660),
.B(n_268),
.C(n_278),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_815),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_800),
.A2(n_649),
.B(n_535),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_SL g1017 ( 
.A(n_785),
.B(n_246),
.C(n_243),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_764),
.B(n_514),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_855),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_874),
.A2(n_710),
.B(n_707),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_858),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_858),
.Y(n_1022)
);

NOR2x2_ASAP7_75t_L g1023 ( 
.A(n_897),
.B(n_254),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_890),
.B(n_722),
.Y(n_1024)
);

NOR2xp67_ASAP7_75t_L g1025 ( 
.A(n_847),
.B(n_660),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_890),
.B(n_259),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_797),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_903),
.B(n_736),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_824),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_839),
.B(n_516),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_767),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_861),
.Y(n_1032)
);

O2A1O1Ixp5_ASAP7_75t_L g1033 ( 
.A1(n_819),
.A2(n_263),
.B(n_287),
.C(n_256),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_861),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_852),
.B(n_516),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_904),
.B(n_736),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_788),
.A2(n_378),
.B(n_322),
.C(n_323),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_867),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_867),
.Y(n_1039)
);

OAI21xp33_ASAP7_75t_L g1040 ( 
.A1(n_899),
.A2(n_366),
.B(n_259),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_906),
.B(n_739),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_870),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_787),
.A2(n_741),
.B(n_739),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_835),
.A2(n_317),
.B(n_326),
.C(n_358),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_832),
.A2(n_744),
.B(n_741),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_811),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_878),
.A2(n_649),
.B(n_535),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_880),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_884),
.A2(n_649),
.B(n_556),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_870),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_802),
.B(n_790),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_898),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_853),
.B(n_744),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_853),
.B(n_746),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_900),
.A2(n_556),
.B(n_547),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_879),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_836),
.A2(n_556),
.B(n_547),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_911),
.A2(n_556),
.B(n_547),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_905),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_875),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_866),
.B(n_366),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_804),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_879),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_885),
.B(n_751),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_791),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_885),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_901),
.A2(n_560),
.B(n_547),
.Y(n_1067)
);

CKINVDCx10_ASAP7_75t_R g1068 ( 
.A(n_794),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_887),
.B(n_896),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_887),
.B(n_751),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_912),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_901),
.A2(n_914),
.B(n_841),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_912),
.B(n_753),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_841),
.A2(n_562),
.B(n_560),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_919),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_781),
.B(n_795),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_898),
.B(n_367),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_781),
.B(n_757),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_881),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_917),
.A2(n_562),
.B(n_560),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_778),
.B(n_757),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_916),
.A2(n_363),
.B(n_391),
.C(n_397),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_916),
.B(n_367),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_888),
.A2(n_399),
.B(n_401),
.C(n_409),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_778),
.B(n_758),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_763),
.B(n_304),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_910),
.B(n_631),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_873),
.B(n_631),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_917),
.A2(n_562),
.B(n_581),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_873),
.A2(n_415),
.B(n_369),
.C(n_374),
.Y(n_1090)
);

BUFx8_ASAP7_75t_SL g1091 ( 
.A(n_794),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_808),
.B(n_577),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_905),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_957),
.B(n_792),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1026),
.A2(n_789),
.B(n_803),
.C(n_817),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_1091),
.Y(n_1096)
);

O2A1O1Ixp5_ASAP7_75t_L g1097 ( 
.A1(n_1012),
.A2(n_862),
.B(n_860),
.C(n_918),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_961),
.B(n_869),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_991),
.B(n_1001),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_991),
.B(n_905),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_925),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_976),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_925),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_929),
.A2(n_843),
.B(n_837),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_1059),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_R g1106 ( 
.A(n_1017),
.B(n_820),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1026),
.B(n_815),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_943),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_926),
.A2(n_849),
.B1(n_845),
.B2(n_815),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_937),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_921),
.A2(n_1015),
.B1(n_1051),
.B2(n_926),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_991),
.B(n_763),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_985),
.B(n_891),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_SL g1114 ( 
.A1(n_1062),
.A2(n_383),
.B1(n_368),
.B2(n_369),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_SL g1115 ( 
.A(n_987),
.B(n_820),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_943),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_955),
.A2(n_894),
.B(n_889),
.C(n_892),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_973),
.B(n_850),
.Y(n_1118)
);

AOI221xp5_ASAP7_75t_L g1119 ( 
.A1(n_985),
.A2(n_886),
.B1(n_909),
.B2(n_416),
.C(n_393),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_973),
.B(n_919),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_924),
.A2(n_862),
.B(n_860),
.Y(n_1121)
);

O2A1O1Ixp5_ASAP7_75t_L g1122 ( 
.A1(n_1011),
.A2(n_918),
.B(n_913),
.C(n_806),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1068),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_933),
.A2(n_917),
.B(n_834),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_971),
.A2(n_907),
.B(n_834),
.C(n_577),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1079),
.B(n_859),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_942),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_941),
.A2(n_848),
.B1(n_876),
.B2(n_413),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_944),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_980),
.A2(n_570),
.B(n_550),
.C(n_568),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_972),
.B(n_848),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_937),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_971),
.B(n_368),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_962),
.A2(n_581),
.B(n_584),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1087),
.A2(n_260),
.B1(n_257),
.B2(n_370),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_SL g1136 ( 
.A1(n_930),
.A2(n_551),
.B(n_557),
.C(n_561),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_L g1137 ( 
.A1(n_935),
.A2(n_587),
.B(n_577),
.C(n_589),
.Y(n_1137)
);

NOR3xp33_ASAP7_75t_SL g1138 ( 
.A(n_1040),
.B(n_408),
.C(n_374),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_991),
.B(n_876),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_989),
.A2(n_876),
.B1(n_253),
.B2(n_257),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_939),
.A2(n_581),
.B(n_584),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1048),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1025),
.A2(n_589),
.B(n_587),
.C(n_577),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_988),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1046),
.B(n_380),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_949),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1018),
.B(n_859),
.Y(n_1147)
);

BUFx2_ASAP7_75t_SL g1148 ( 
.A(n_988),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_936),
.A2(n_876),
.B(n_589),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1072),
.A2(n_589),
.B(n_587),
.C(n_253),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_955),
.A2(n_551),
.B(n_557),
.C(n_561),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_992),
.A2(n_260),
.B1(n_402),
.B2(n_375),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1030),
.B(n_859),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_1065),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1051),
.B(n_859),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_956),
.B(n_380),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1001),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1048),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_SL g1159 ( 
.A1(n_1004),
.A2(n_566),
.B(n_567),
.C(n_568),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1052),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_982),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1076),
.A2(n_589),
.B(n_587),
.C(n_382),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_932),
.A2(n_587),
.B(n_413),
.C(n_407),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1035),
.Y(n_1164)
);

BUFx10_ASAP7_75t_L g1165 ( 
.A(n_1077),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_SL g1166 ( 
.A1(n_1004),
.A2(n_591),
.B(n_567),
.C(n_569),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1060),
.A2(n_876),
.B1(n_394),
.B2(n_402),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1082),
.A2(n_389),
.B(n_407),
.C(n_406),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_1052),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_986),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_986),
.B(n_859),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1000),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1037),
.A2(n_389),
.B(n_406),
.C(n_405),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_945),
.A2(n_590),
.B(n_588),
.Y(n_1174)
);

OR2x6_ASAP7_75t_SL g1175 ( 
.A(n_996),
.B(n_381),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1090),
.A2(n_405),
.B(n_403),
.C(n_390),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1002),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_1077),
.Y(n_1178)
);

AO21x1_ASAP7_75t_L g1179 ( 
.A1(n_1086),
.A2(n_591),
.B(n_607),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1092),
.A2(n_390),
.B1(n_394),
.B2(n_403),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_997),
.A2(n_934),
.B(n_948),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_1083),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1003),
.B(n_381),
.Y(n_1183)
);

INVx3_ASAP7_75t_SL g1184 ( 
.A(n_1023),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1008),
.B(n_695),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_953),
.A2(n_590),
.B(n_588),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1059),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_981),
.A2(n_1010),
.B1(n_1024),
.B2(n_1007),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_979),
.B(n_77),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1083),
.B(n_383),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1019),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_922),
.A2(n_590),
.B(n_588),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1001),
.B(n_385),
.Y(n_1193)
);

AOI21xp33_ASAP7_75t_L g1194 ( 
.A1(n_1088),
.A2(n_396),
.B(n_385),
.Y(n_1194)
);

NOR3xp33_ASAP7_75t_SL g1195 ( 
.A(n_1090),
.B(n_395),
.C(n_393),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1061),
.B(n_395),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_927),
.A2(n_590),
.B(n_586),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1001),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1092),
.A2(n_695),
.B1(n_566),
.B2(n_607),
.Y(n_1199)
);

INVx5_ASAP7_75t_L g1200 ( 
.A(n_1059),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1019),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1032),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_959),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1032),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_959),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_981),
.A2(n_304),
.B1(n_400),
.B2(n_396),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_923),
.A2(n_695),
.B1(n_400),
.B2(n_596),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_979),
.B(n_412),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1029),
.Y(n_1209)
);

INVx4_ASAP7_75t_L g1210 ( 
.A(n_1059),
.Y(n_1210)
);

AO21x1_ASAP7_75t_L g1211 ( 
.A1(n_1053),
.A2(n_574),
.B(n_582),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1031),
.A2(n_400),
.B1(n_412),
.B2(n_414),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1093),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1054),
.A2(n_1044),
.B(n_1014),
.C(n_1084),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1029),
.B(n_414),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_SL g1216 ( 
.A(n_967),
.B(n_416),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1034),
.B(n_695),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1034),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1031),
.A2(n_695),
.B1(n_400),
.B2(n_596),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_1081),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1069),
.A2(n_569),
.B(n_582),
.C(n_585),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1093),
.Y(n_1222)
);

AO22x1_ASAP7_75t_L g1223 ( 
.A1(n_1027),
.A2(n_585),
.B1(n_602),
.B2(n_11),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1093),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1039),
.B(n_602),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1027),
.A2(n_586),
.B1(n_588),
.B2(n_605),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_920),
.A2(n_599),
.B(n_592),
.C(n_605),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1039),
.Y(n_1228)
);

AOI22x1_ASAP7_75t_L g1229 ( 
.A1(n_1021),
.A2(n_599),
.B1(n_592),
.B2(n_605),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_940),
.A2(n_599),
.B(n_592),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_942),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_950),
.A2(n_599),
.B(n_592),
.Y(n_1232)
);

AO21x2_ASAP7_75t_L g1233 ( 
.A1(n_952),
.A2(n_586),
.B(n_595),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_947),
.A2(n_595),
.B(n_606),
.C(n_604),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_964),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_954),
.A2(n_595),
.B(n_606),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_938),
.B(n_148),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_965),
.B(n_8),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1056),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_969),
.B(n_609),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1093),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_960),
.A2(n_606),
.B(n_604),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_967),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_942),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_942),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1006),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1235),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1094),
.B(n_1022),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1101),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1125),
.A2(n_1005),
.B(n_963),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1118),
.A2(n_946),
.B(n_966),
.C(n_1038),
.Y(n_1251)
);

NAND2x2_ASAP7_75t_L g1252 ( 
.A(n_1243),
.B(n_1013),
.Y(n_1252)
);

INVx3_ASAP7_75t_SL g1253 ( 
.A(n_1123),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1211),
.A2(n_1071),
.A3(n_1063),
.B(n_1042),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1102),
.Y(n_1255)
);

AOI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1133),
.A2(n_1050),
.B1(n_1066),
.B2(n_1085),
.Y(n_1256)
);

OAI22x1_ASAP7_75t_L g1257 ( 
.A1(n_1178),
.A2(n_931),
.B1(n_951),
.B2(n_958),
.Y(n_1257)
);

AND2x6_ASAP7_75t_SL g1258 ( 
.A(n_1183),
.B(n_977),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1190),
.A2(n_970),
.B(n_1033),
.C(n_994),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1111),
.A2(n_994),
.B1(n_928),
.B2(n_958),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1178),
.A2(n_928),
.B1(n_951),
.B2(n_931),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1182),
.B(n_1075),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1182),
.B(n_978),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1246),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1095),
.A2(n_1119),
.B(n_1156),
.C(n_1107),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1163),
.A2(n_1078),
.B(n_1058),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1103),
.Y(n_1267)
);

BUFx2_ASAP7_75t_R g1268 ( 
.A(n_1096),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1188),
.A2(n_1064),
.B(n_1070),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1203),
.B(n_974),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1146),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1197),
.A2(n_993),
.B(n_1009),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1161),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1220),
.B(n_983),
.Y(n_1274)
);

O2A1O1Ixp5_ASAP7_75t_L g1275 ( 
.A1(n_1098),
.A2(n_974),
.B(n_975),
.C(n_1043),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1119),
.A2(n_999),
.B(n_1028),
.C(n_1036),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1197),
.A2(n_1020),
.B(n_998),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1108),
.Y(n_1278)
);

AND2x4_ASAP7_75t_SL g1279 ( 
.A(n_1210),
.B(n_598),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1110),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1113),
.B(n_1041),
.Y(n_1281)
);

AOI221x1_ASAP7_75t_L g1282 ( 
.A1(n_1109),
.A2(n_1047),
.B1(n_1049),
.B2(n_1045),
.C(n_1057),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_SL g1283 ( 
.A(n_1106),
.B(n_1073),
.C(n_1055),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1121),
.A2(n_975),
.B(n_995),
.Y(n_1284)
);

AOI21xp33_ASAP7_75t_L g1285 ( 
.A1(n_1164),
.A2(n_1215),
.B(n_1208),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1157),
.B(n_990),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1170),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1160),
.Y(n_1288)
);

CKINVDCx16_ASAP7_75t_R g1289 ( 
.A(n_1115),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1121),
.A2(n_968),
.B(n_984),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1165),
.B(n_1067),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1172),
.Y(n_1292)
);

NOR2x1_ASAP7_75t_SL g1293 ( 
.A(n_1200),
.B(n_598),
.Y(n_1293)
);

AOI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1124),
.A2(n_1242),
.B(n_1236),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1149),
.A2(n_1016),
.B(n_1074),
.Y(n_1295)
);

AO31x2_ASAP7_75t_L g1296 ( 
.A1(n_1179),
.A2(n_1089),
.A3(n_1080),
.B(n_12),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1097),
.A2(n_609),
.B(n_606),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1196),
.B(n_9),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1142),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1214),
.A2(n_142),
.B(n_104),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1149),
.A2(n_609),
.B(n_606),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1116),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1200),
.Y(n_1303)
);

AO32x2_ASAP7_75t_L g1304 ( 
.A1(n_1206),
.A2(n_1135),
.A3(n_1212),
.B1(n_1226),
.B2(n_1152),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1158),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1191),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1129),
.Y(n_1307)
);

OA22x2_ASAP7_75t_L g1308 ( 
.A1(n_1114),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1220),
.B(n_14),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1205),
.B(n_14),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1201),
.Y(n_1311)
);

AO21x1_ASAP7_75t_L g1312 ( 
.A1(n_1117),
.A2(n_16),
.B(n_20),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1169),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1228),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1132),
.Y(n_1315)
);

AO31x2_ASAP7_75t_L g1316 ( 
.A1(n_1150),
.A2(n_21),
.A3(n_22),
.B(n_24),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1154),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1194),
.B(n_22),
.Y(n_1318)
);

CKINVDCx8_ASAP7_75t_R g1319 ( 
.A(n_1148),
.Y(n_1319)
);

NAND2x1p5_ASAP7_75t_L g1320 ( 
.A(n_1200),
.B(n_609),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1198),
.Y(n_1321)
);

INVx4_ASAP7_75t_L g1322 ( 
.A(n_1200),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1144),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1145),
.B(n_25),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1184),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1097),
.A2(n_139),
.B(n_108),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1231),
.Y(n_1327)
);

NOR2xp67_ASAP7_75t_L g1328 ( 
.A(n_1140),
.B(n_207),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1176),
.A2(n_604),
.B1(n_598),
.B2(n_31),
.C(n_32),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1112),
.A2(n_604),
.B(n_598),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1131),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1242),
.A2(n_160),
.B(n_113),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1233),
.A2(n_604),
.B(n_598),
.Y(n_1333)
);

AOI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1236),
.A2(n_604),
.B(n_598),
.Y(n_1334)
);

AOI221xp5_ASAP7_75t_L g1335 ( 
.A1(n_1138),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.C(n_35),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_R g1336 ( 
.A(n_1216),
.B(n_206),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1165),
.B(n_28),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1192),
.A2(n_198),
.B(n_187),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1117),
.A2(n_47),
.B(n_48),
.C(n_50),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1239),
.B(n_48),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1233),
.A2(n_184),
.B(n_178),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1195),
.B(n_51),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1234),
.A2(n_51),
.A3(n_53),
.B(n_54),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1177),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1105),
.Y(n_1345)
);

AOI221xp5_ASAP7_75t_L g1346 ( 
.A1(n_1238),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.C(n_60),
.Y(n_1346)
);

NOR2xp67_ASAP7_75t_L g1347 ( 
.A(n_1210),
.B(n_91),
.Y(n_1347)
);

INVx5_ASAP7_75t_L g1348 ( 
.A(n_1105),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1128),
.A2(n_1193),
.B1(n_1189),
.B2(n_1180),
.Y(n_1349)
);

AO31x2_ASAP7_75t_L g1350 ( 
.A1(n_1162),
.A2(n_55),
.A3(n_62),
.B(n_66),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1189),
.A2(n_62),
.B1(n_66),
.B2(n_68),
.Y(n_1351)
);

AOI221x1_ASAP7_75t_L g1352 ( 
.A1(n_1168),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.C(n_73),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1202),
.B(n_69),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1147),
.A2(n_124),
.B(n_172),
.Y(n_1354)
);

O2A1O1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1136),
.A2(n_71),
.B(n_72),
.C(n_74),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1209),
.Y(n_1356)
);

INVx6_ASAP7_75t_SL g1357 ( 
.A(n_1237),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1105),
.Y(n_1358)
);

NOR2x1_ASAP7_75t_L g1359 ( 
.A(n_1245),
.B(n_125),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1204),
.B(n_74),
.Y(n_1360)
);

BUFx3_ASAP7_75t_L g1361 ( 
.A(n_1187),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1192),
.A2(n_119),
.B(n_120),
.Y(n_1362)
);

INVx6_ASAP7_75t_L g1363 ( 
.A(n_1187),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1187),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1218),
.B(n_75),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1237),
.B(n_132),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1225),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1151),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1213),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1167),
.B(n_1153),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1230),
.A2(n_135),
.B(n_138),
.Y(n_1371)
);

INVx5_ASAP7_75t_L g1372 ( 
.A(n_1213),
.Y(n_1372)
);

AND2x2_ASAP7_75t_SL g1373 ( 
.A(n_1213),
.B(n_176),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1173),
.A2(n_1137),
.B(n_1122),
.C(n_1143),
.Y(n_1374)
);

AO21x1_ASAP7_75t_L g1375 ( 
.A1(n_1221),
.A2(n_1126),
.B(n_1151),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1137),
.A2(n_1122),
.B(n_1221),
.C(n_1199),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1229),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1223),
.A2(n_1155),
.B1(n_1099),
.B2(n_1100),
.Y(n_1378)
);

AO31x2_ASAP7_75t_L g1379 ( 
.A1(n_1230),
.A2(n_1232),
.A3(n_1227),
.B(n_1186),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1232),
.A2(n_1186),
.A3(n_1174),
.B(n_1141),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1155),
.A2(n_1139),
.B1(n_1244),
.B2(n_1127),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1171),
.A2(n_1217),
.B1(n_1185),
.B2(n_1207),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1175),
.B(n_1127),
.Y(n_1383)
);

OAI21xp33_ASAP7_75t_L g1384 ( 
.A1(n_1219),
.A2(n_1240),
.B(n_1134),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1244),
.B(n_1245),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1159),
.A2(n_1166),
.B(n_1130),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1222),
.A2(n_1224),
.B(n_1241),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1222),
.A2(n_1224),
.B(n_1241),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1222),
.A2(n_1224),
.B(n_1241),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1181),
.A2(n_997),
.B(n_934),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1118),
.A2(n_1121),
.B(n_1104),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1120),
.A2(n_654),
.B(n_957),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1113),
.B(n_805),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1118),
.A2(n_801),
.B1(n_1094),
.B2(n_957),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1181),
.A2(n_997),
.B(n_934),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1133),
.A2(n_1026),
.B1(n_1118),
.B2(n_1190),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1211),
.A2(n_1179),
.A3(n_1188),
.B(n_1150),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1101),
.Y(n_1398)
);

NOR2xp67_ASAP7_75t_L g1399 ( 
.A(n_1200),
.B(n_980),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1118),
.A2(n_1094),
.B(n_801),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1102),
.B(n_768),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1308),
.A2(n_1373),
.B1(n_1336),
.B2(n_1300),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1396),
.A2(n_1393),
.B1(n_1318),
.B2(n_1394),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1253),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1400),
.B(n_1396),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1248),
.B(n_1265),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1348),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1348),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1346),
.A2(n_1328),
.B1(n_1401),
.B2(n_1335),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1280),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1328),
.A2(n_1324),
.B1(n_1285),
.B2(n_1349),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1289),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1249),
.Y(n_1413)
);

CKINVDCx11_ASAP7_75t_R g1414 ( 
.A(n_1319),
.Y(n_1414)
);

INVx6_ASAP7_75t_L g1415 ( 
.A(n_1348),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1298),
.A2(n_1342),
.B1(n_1326),
.B2(n_1366),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_SL g1417 ( 
.A1(n_1366),
.A2(n_1354),
.B1(n_1281),
.B2(n_1260),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1367),
.B(n_1274),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1251),
.B(n_1263),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1349),
.A2(n_1351),
.B1(n_1312),
.B2(n_1337),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1255),
.B(n_1270),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1247),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1351),
.A2(n_1352),
.B1(n_1366),
.B2(n_1309),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1325),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1383),
.A2(n_1331),
.B1(n_1317),
.B2(n_1255),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1270),
.A2(n_1370),
.B1(n_1368),
.B2(n_1317),
.Y(n_1426)
);

BUFx2_ASAP7_75t_SL g1427 ( 
.A(n_1315),
.Y(n_1427)
);

BUFx8_ASAP7_75t_L g1428 ( 
.A(n_1313),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1391),
.A2(n_1299),
.B1(n_1332),
.B2(n_1305),
.Y(n_1429)
);

CKINVDCx11_ASAP7_75t_R g1430 ( 
.A(n_1258),
.Y(n_1430)
);

INVx6_ASAP7_75t_L g1431 ( 
.A(n_1372),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1291),
.A2(n_1283),
.B1(n_1357),
.B2(n_1310),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1357),
.A2(n_1391),
.B1(n_1288),
.B2(n_1340),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1252),
.A2(n_1375),
.B1(n_1360),
.B2(n_1365),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1278),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1264),
.Y(n_1436)
);

INVx6_ASAP7_75t_L g1437 ( 
.A(n_1372),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1302),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1303),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1305),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1307),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1268),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1344),
.Y(n_1443)
);

INVx6_ASAP7_75t_L g1444 ( 
.A(n_1372),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1353),
.A2(n_1256),
.B1(n_1257),
.B2(n_1327),
.Y(n_1445)
);

BUFx2_ASAP7_75t_SL g1446 ( 
.A(n_1323),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1378),
.A2(n_1356),
.B1(n_1256),
.B2(n_1262),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1267),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1321),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1339),
.A2(n_1259),
.B1(n_1378),
.B2(n_1376),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1271),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1356),
.B(n_1398),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1258),
.Y(n_1453)
);

BUFx2_ASAP7_75t_SL g1454 ( 
.A(n_1361),
.Y(n_1454)
);

INVx6_ASAP7_75t_L g1455 ( 
.A(n_1345),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1392),
.A2(n_1286),
.B1(n_1292),
.B2(n_1306),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1273),
.B(n_1287),
.Y(n_1457)
);

OAI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1311),
.A2(n_1314),
.B1(n_1382),
.B2(n_1261),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1332),
.A2(n_1329),
.B1(n_1250),
.B2(n_1355),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1374),
.A2(n_1381),
.B1(n_1276),
.B2(n_1399),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1388),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1254),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1350),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1363),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1286),
.A2(n_1266),
.B1(n_1384),
.B2(n_1359),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1350),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1386),
.A2(n_1347),
.B1(n_1341),
.B2(n_1385),
.Y(n_1467)
);

OAI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1382),
.A2(n_1347),
.B1(n_1329),
.B2(n_1269),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1364),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1363),
.Y(n_1470)
);

CKINVDCx11_ASAP7_75t_R g1471 ( 
.A(n_1369),
.Y(n_1471)
);

INVx5_ASAP7_75t_L g1472 ( 
.A(n_1358),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1369),
.A2(n_1389),
.B1(n_1320),
.B2(n_1387),
.Y(n_1473)
);

OAI21xp33_ASAP7_75t_L g1474 ( 
.A1(n_1371),
.A2(n_1294),
.B(n_1297),
.Y(n_1474)
);

INVx6_ASAP7_75t_L g1475 ( 
.A(n_1279),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1350),
.Y(n_1476)
);

BUFx2_ASAP7_75t_SL g1477 ( 
.A(n_1377),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1293),
.A2(n_1362),
.B1(n_1338),
.B2(n_1277),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1316),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1316),
.Y(n_1480)
);

INVx6_ASAP7_75t_L g1481 ( 
.A(n_1275),
.Y(n_1481)
);

OAI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1282),
.A2(n_1284),
.B1(n_1297),
.B2(n_1304),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1334),
.A2(n_1290),
.B1(n_1304),
.B2(n_1295),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1316),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1343),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1343),
.Y(n_1486)
);

OAI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1304),
.A2(n_1301),
.B1(n_1333),
.B2(n_1330),
.Y(n_1487)
);

CKINVDCx11_ASAP7_75t_R g1488 ( 
.A(n_1343),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1296),
.Y(n_1489)
);

INVx3_ASAP7_75t_L g1490 ( 
.A(n_1296),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1397),
.B(n_1380),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1397),
.A2(n_1379),
.B1(n_1380),
.B2(n_1390),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1395),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1380),
.Y(n_1494)
);

BUFx8_ASAP7_75t_L g1495 ( 
.A(n_1397),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1272),
.A2(n_525),
.B1(n_921),
.B2(n_1133),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1379),
.A2(n_525),
.B1(n_921),
.B2(n_1133),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1379),
.A2(n_1396),
.B1(n_1026),
.B2(n_1133),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1247),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1348),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1396),
.A2(n_1026),
.B1(n_1133),
.B2(n_1118),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1396),
.A2(n_1351),
.B1(n_1118),
.B2(n_633),
.Y(n_1502)
);

CKINVDCx6p67_ASAP7_75t_R g1503 ( 
.A(n_1253),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1396),
.A2(n_771),
.B1(n_786),
.B2(n_926),
.Y(n_1504)
);

INVx4_ASAP7_75t_L g1505 ( 
.A(n_1348),
.Y(n_1505)
);

INVx6_ASAP7_75t_L g1506 ( 
.A(n_1348),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1247),
.Y(n_1507)
);

BUFx10_ASAP7_75t_L g1508 ( 
.A(n_1325),
.Y(n_1508)
);

INVx8_ASAP7_75t_L g1509 ( 
.A(n_1348),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1280),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1249),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1249),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1288),
.Y(n_1513)
);

CKINVDCx12_ASAP7_75t_R g1514 ( 
.A(n_1366),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1396),
.A2(n_1026),
.B1(n_1133),
.B2(n_1118),
.Y(n_1515)
);

CKINVDCx6p67_ASAP7_75t_R g1516 ( 
.A(n_1253),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1396),
.A2(n_616),
.B(n_633),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1396),
.A2(n_1026),
.B1(n_1133),
.B2(n_1118),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1348),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1280),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1250),
.A2(n_1391),
.B(n_1392),
.Y(n_1521)
);

CKINVDCx6p67_ASAP7_75t_R g1522 ( 
.A(n_1253),
.Y(n_1522)
);

NAND2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1322),
.B(n_1200),
.Y(n_1523)
);

OAI22x1_ASAP7_75t_L g1524 ( 
.A1(n_1396),
.A2(n_1351),
.B1(n_633),
.B2(n_1349),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1322),
.Y(n_1525)
);

BUFx2_ASAP7_75t_SL g1526 ( 
.A(n_1319),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_1253),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1247),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1396),
.A2(n_771),
.B1(n_786),
.B2(n_926),
.Y(n_1529)
);

OAI22x1_ASAP7_75t_L g1530 ( 
.A1(n_1396),
.A2(n_1351),
.B1(n_633),
.B2(n_1349),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1247),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1249),
.Y(n_1532)
);

BUFx8_ASAP7_75t_L g1533 ( 
.A(n_1313),
.Y(n_1533)
);

INVx6_ASAP7_75t_L g1534 ( 
.A(n_1348),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1253),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1396),
.A2(n_1026),
.B1(n_1133),
.B2(n_1118),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1308),
.A2(n_525),
.B1(n_921),
.B2(n_1133),
.Y(n_1537)
);

BUFx8_ASAP7_75t_L g1538 ( 
.A(n_1313),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1249),
.Y(n_1539)
);

INVx5_ASAP7_75t_L g1540 ( 
.A(n_1322),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1280),
.Y(n_1541)
);

BUFx8_ASAP7_75t_SL g1542 ( 
.A(n_1325),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1348),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1396),
.A2(n_771),
.B1(n_786),
.B2(n_926),
.Y(n_1544)
);

AO22x1_ASAP7_75t_L g1545 ( 
.A1(n_1281),
.A2(n_676),
.B1(n_1026),
.B2(n_1133),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1396),
.A2(n_1026),
.B1(n_1133),
.B2(n_1118),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1255),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1348),
.Y(n_1548)
);

INVx6_ASAP7_75t_L g1549 ( 
.A(n_1348),
.Y(n_1549)
);

INVx6_ASAP7_75t_L g1550 ( 
.A(n_1348),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1393),
.B(n_805),
.Y(n_1551)
);

BUFx12f_ASAP7_75t_L g1552 ( 
.A(n_1325),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1393),
.B(n_805),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_SL g1554 ( 
.A1(n_1308),
.A2(n_525),
.B1(n_921),
.B2(n_1133),
.Y(n_1554)
);

INVx4_ASAP7_75t_L g1555 ( 
.A(n_1348),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1396),
.A2(n_1118),
.B1(n_1026),
.B2(n_1190),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1396),
.A2(n_1026),
.B1(n_1133),
.B2(n_1118),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1249),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1280),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1253),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1495),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1462),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1495),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1463),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1418),
.B(n_1556),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1422),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1448),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1451),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1491),
.B(n_1479),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1491),
.B(n_1480),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1497),
.B(n_1466),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1440),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1513),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1494),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1436),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1501),
.A2(n_1518),
.B(n_1515),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1499),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1497),
.B(n_1476),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1485),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_R g1580 ( 
.A(n_1442),
.B(n_1414),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1484),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1486),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1489),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1490),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1507),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1461),
.Y(n_1586)
);

OR2x6_ASAP7_75t_L g1587 ( 
.A(n_1521),
.B(n_1450),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1528),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1481),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1481),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1405),
.B(n_1421),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1493),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1492),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1405),
.B(n_1406),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1418),
.B(n_1536),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1531),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1457),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1457),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1481),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1496),
.B(n_1498),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1452),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1493),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1546),
.B(n_1557),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1509),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1403),
.B(n_1502),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1547),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1443),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1551),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1493),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1458),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1406),
.B(n_1419),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1413),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1435),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1449),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1438),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1514),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1441),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1511),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1512),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_SL g1620 ( 
.A(n_1428),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1532),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1502),
.B(n_1419),
.Y(n_1622)
);

A2O1A1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1517),
.A2(n_1529),
.B(n_1504),
.C(n_1544),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1539),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1558),
.Y(n_1625)
);

AO21x2_ASAP7_75t_L g1626 ( 
.A1(n_1468),
.A2(n_1474),
.B(n_1482),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1411),
.B(n_1402),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1412),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1483),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1458),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1496),
.B(n_1524),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1530),
.B(n_1488),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1477),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1447),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1509),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1450),
.B(n_1460),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1439),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1428),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1439),
.Y(n_1639)
);

AO21x2_ASAP7_75t_L g1640 ( 
.A1(n_1468),
.A2(n_1482),
.B(n_1487),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1467),
.A2(n_1456),
.B(n_1465),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1426),
.B(n_1429),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1429),
.B(n_1416),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1460),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1509),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1473),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1473),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1537),
.B(n_1554),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1540),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1459),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1537),
.B(n_1554),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1434),
.A2(n_1445),
.B(n_1432),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1420),
.A2(n_1433),
.B(n_1409),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1540),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1459),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1478),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1540),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1533),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1525),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1523),
.A2(n_1478),
.B(n_1529),
.Y(n_1660)
);

O2A1O1Ixp5_ASAP7_75t_L g1661 ( 
.A1(n_1545),
.A2(n_1544),
.B(n_1504),
.C(n_1423),
.Y(n_1661)
);

AO32x1_ASAP7_75t_L g1662 ( 
.A1(n_1423),
.A2(n_1416),
.A3(n_1555),
.B1(n_1519),
.B2(n_1408),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1472),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1417),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1417),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1540),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1533),
.Y(n_1667)
);

INVx2_ASAP7_75t_SL g1668 ( 
.A(n_1407),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1472),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1523),
.Y(n_1670)
);

OR2x6_ASAP7_75t_L g1671 ( 
.A(n_1526),
.B(n_1427),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1407),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1542),
.Y(n_1673)
);

AOI222xp33_ASAP7_75t_L g1674 ( 
.A1(n_1553),
.A2(n_1453),
.B1(n_1430),
.B2(n_1425),
.C1(n_1402),
.C2(n_1538),
.Y(n_1674)
);

AO31x2_ASAP7_75t_L g1675 ( 
.A1(n_1408),
.A2(n_1505),
.A3(n_1548),
.B(n_1519),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1538),
.A2(n_1446),
.B1(n_1407),
.B2(n_1534),
.Y(n_1676)
);

BUFx2_ASAP7_75t_SL g1677 ( 
.A(n_1505),
.Y(n_1677)
);

AOI222xp33_ASAP7_75t_L g1678 ( 
.A1(n_1424),
.A2(n_1552),
.B1(n_1471),
.B2(n_1559),
.C1(n_1410),
.C2(n_1541),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1415),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1475),
.A2(n_1510),
.B1(n_1520),
.B2(n_1431),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1415),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1415),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1431),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1469),
.B(n_1455),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1454),
.B(n_1469),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1437),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1548),
.B(n_1555),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1470),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1469),
.B(n_1464),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1437),
.Y(n_1690)
);

AO21x1_ASAP7_75t_L g1691 ( 
.A1(n_1437),
.A2(n_1549),
.B(n_1444),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1503),
.B(n_1522),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1444),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1444),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1500),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1475),
.A2(n_1543),
.B1(n_1534),
.B2(n_1500),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1609),
.B(n_1592),
.Y(n_1697)
);

OR2x6_ASAP7_75t_L g1698 ( 
.A(n_1587),
.B(n_1475),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1609),
.B(n_1527),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1627),
.B(n_1534),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1578),
.B(n_1455),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1578),
.B(n_1516),
.Y(n_1702)
);

OAI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1636),
.A2(n_1543),
.B1(n_1506),
.B2(n_1550),
.Y(n_1703)
);

INVx4_ASAP7_75t_L g1704 ( 
.A(n_1649),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1571),
.B(n_1543),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1601),
.B(n_1404),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1634),
.B(n_1506),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1573),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1581),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1661),
.A2(n_1560),
.B1(n_1535),
.B2(n_1508),
.C(n_1550),
.Y(n_1710)
);

AO21x2_ASAP7_75t_L g1711 ( 
.A1(n_1623),
.A2(n_1549),
.B(n_1550),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1591),
.B(n_1508),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1591),
.B(n_1632),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1576),
.A2(n_1648),
.B(n_1651),
.C(n_1652),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1632),
.B(n_1631),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1594),
.B(n_1611),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1592),
.B(n_1602),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1674),
.A2(n_1631),
.B(n_1603),
.C(n_1665),
.Y(n_1718)
);

INVx5_ASAP7_75t_SL g1719 ( 
.A(n_1671),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1628),
.Y(n_1720)
);

NOR2x1_ASAP7_75t_SL g1721 ( 
.A(n_1587),
.B(n_1636),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1643),
.B(n_1600),
.Y(n_1722)
);

NAND2xp33_ASAP7_75t_L g1723 ( 
.A(n_1605),
.B(n_1622),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1587),
.B(n_1636),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1600),
.B(n_1608),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1664),
.B(n_1665),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1571),
.B(n_1656),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1636),
.A2(n_1595),
.B1(n_1587),
.B2(n_1664),
.Y(n_1728)
);

NOR2x1_ASAP7_75t_SL g1729 ( 
.A(n_1599),
.B(n_1671),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1565),
.A2(n_1676),
.B1(n_1653),
.B2(n_1671),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1597),
.B(n_1598),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1599),
.B(n_1644),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_1604),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_SL g1734 ( 
.A(n_1673),
.B(n_1628),
.Y(n_1734)
);

O2A1O1Ixp33_ASAP7_75t_SL g1735 ( 
.A1(n_1633),
.A2(n_1655),
.B(n_1650),
.C(n_1696),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1602),
.B(n_1567),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1652),
.A2(n_1641),
.B(n_1653),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1568),
.B(n_1575),
.Y(n_1738)
);

INVxp67_ASAP7_75t_L g1739 ( 
.A(n_1606),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1589),
.B(n_1590),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1671),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1590),
.B(n_1691),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1607),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1616),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1581),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1630),
.B(n_1647),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1653),
.A2(n_1610),
.B1(n_1642),
.B2(n_1655),
.Y(n_1747)
);

AOI21x1_ASAP7_75t_L g1748 ( 
.A1(n_1691),
.A2(n_1680),
.B(n_1650),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1577),
.B(n_1585),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1662),
.A2(n_1640),
.B(n_1626),
.Y(n_1750)
);

OA21x2_ASAP7_75t_L g1751 ( 
.A1(n_1660),
.A2(n_1641),
.B(n_1593),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1673),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1662),
.A2(n_1640),
.B(n_1626),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1596),
.B(n_1607),
.Y(n_1754)
);

OA21x2_ASAP7_75t_L g1755 ( 
.A1(n_1660),
.A2(n_1593),
.B(n_1629),
.Y(n_1755)
);

OR2x6_ASAP7_75t_L g1756 ( 
.A(n_1646),
.B(n_1610),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1566),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1637),
.Y(n_1758)
);

INVx4_ASAP7_75t_L g1759 ( 
.A(n_1649),
.Y(n_1759)
);

OAI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1653),
.A2(n_1688),
.B(n_1670),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_SL g1761 ( 
.A1(n_1668),
.A2(n_1685),
.B(n_1663),
.C(n_1670),
.Y(n_1761)
);

OAI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1614),
.A2(n_1572),
.B(n_1687),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1612),
.B(n_1613),
.Y(n_1763)
);

OA21x2_ASAP7_75t_L g1764 ( 
.A1(n_1629),
.A2(n_1582),
.B(n_1579),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1588),
.B(n_1561),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1687),
.A2(n_1672),
.B(n_1693),
.Y(n_1766)
);

O2A1O1Ixp33_ASAP7_75t_L g1767 ( 
.A1(n_1626),
.A2(n_1640),
.B(n_1672),
.C(n_1693),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1586),
.B(n_1564),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1564),
.Y(n_1769)
);

OA21x2_ASAP7_75t_L g1770 ( 
.A1(n_1579),
.A2(n_1582),
.B(n_1583),
.Y(n_1770)
);

NOR4xp25_ASAP7_75t_SL g1771 ( 
.A(n_1561),
.B(n_1563),
.C(n_1662),
.D(n_1586),
.Y(n_1771)
);

OAI211xp5_ASAP7_75t_L g1772 ( 
.A1(n_1678),
.A2(n_1563),
.B(n_1615),
.C(n_1619),
.Y(n_1772)
);

A2O1A1Ixp33_ASAP7_75t_L g1773 ( 
.A1(n_1662),
.A2(n_1668),
.B(n_1657),
.C(n_1666),
.Y(n_1773)
);

CKINVDCx20_ASAP7_75t_R g1774 ( 
.A(n_1580),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1679),
.B(n_1690),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1569),
.B(n_1570),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1770),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1715),
.B(n_1727),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1776),
.B(n_1570),
.Y(n_1779)
);

INVxp67_ASAP7_75t_SL g1780 ( 
.A(n_1764),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1738),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1770),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1776),
.B(n_1584),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1718),
.A2(n_1658),
.B1(n_1667),
.B2(n_1638),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1713),
.B(n_1562),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1714),
.A2(n_1620),
.B1(n_1662),
.B2(n_1638),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1738),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1770),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1716),
.B(n_1574),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1764),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1714),
.A2(n_1773),
.B1(n_1747),
.B2(n_1753),
.Y(n_1791)
);

INVx4_ASAP7_75t_L g1792 ( 
.A(n_1711),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1756),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1723),
.A2(n_1658),
.B1(n_1667),
.B2(n_1617),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1769),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1722),
.B(n_1639),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1706),
.B(n_1692),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1769),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_SL g1799 ( 
.A1(n_1710),
.A2(n_1772),
.B(n_1728),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1709),
.B(n_1618),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1736),
.B(n_1697),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_SL g1802 ( 
.A(n_1703),
.B(n_1604),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1723),
.A2(n_1621),
.B1(n_1624),
.B2(n_1625),
.Y(n_1803)
);

AND2x4_ASAP7_75t_SL g1804 ( 
.A(n_1698),
.B(n_1657),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1700),
.A2(n_1695),
.B1(n_1694),
.B2(n_1683),
.Y(n_1805)
);

CKINVDCx14_ASAP7_75t_R g1806 ( 
.A(n_1720),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1725),
.B(n_1669),
.Y(n_1807)
);

BUFx2_ASAP7_75t_SL g1808 ( 
.A(n_1741),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1756),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1745),
.Y(n_1810)
);

BUFx2_ASAP7_75t_L g1811 ( 
.A(n_1741),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1731),
.B(n_1749),
.Y(n_1812)
);

INVx3_ASAP7_75t_L g1813 ( 
.A(n_1738),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1717),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1701),
.B(n_1659),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1700),
.A2(n_1695),
.B1(n_1694),
.B2(n_1683),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1724),
.A2(n_1692),
.B1(n_1689),
.B2(n_1686),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1801),
.B(n_1751),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1795),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1793),
.B(n_1729),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1801),
.B(n_1751),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1790),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1779),
.B(n_1755),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1793),
.B(n_1721),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1790),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1810),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1791),
.A2(n_1750),
.B1(n_1767),
.B2(n_1737),
.C(n_1760),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1801),
.B(n_1751),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1812),
.B(n_1768),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1812),
.B(n_1754),
.Y(n_1830)
);

OAI321xp33_ASAP7_75t_L g1831 ( 
.A1(n_1786),
.A2(n_1730),
.A3(n_1748),
.B1(n_1773),
.B2(n_1742),
.C(n_1707),
.Y(n_1831)
);

BUFx3_ASAP7_75t_L g1832 ( 
.A(n_1811),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1801),
.B(n_1724),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1778),
.B(n_1724),
.Y(n_1834)
);

INVxp67_ASAP7_75t_L g1835 ( 
.A(n_1807),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_R g1836 ( 
.A(n_1806),
.B(n_1720),
.Y(n_1836)
);

OAI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1799),
.A2(n_1744),
.B1(n_1762),
.B2(n_1707),
.C(n_1735),
.Y(n_1837)
);

OR2x6_ASAP7_75t_L g1838 ( 
.A(n_1808),
.B(n_1724),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1798),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1783),
.B(n_1754),
.Y(n_1840)
);

CKINVDCx20_ASAP7_75t_R g1841 ( 
.A(n_1784),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1798),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1786),
.A2(n_1771),
.B1(n_1746),
.B2(n_1732),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1783),
.B(n_1754),
.Y(n_1844)
);

INVxp67_ASAP7_75t_SL g1845 ( 
.A(n_1810),
.Y(n_1845)
);

XNOR2xp5_ASAP7_75t_L g1846 ( 
.A(n_1784),
.B(n_1774),
.Y(n_1846)
);

OA21x2_ASAP7_75t_L g1847 ( 
.A1(n_1777),
.A2(n_1742),
.B(n_1766),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1799),
.A2(n_1746),
.B1(n_1732),
.B2(n_1739),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1777),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1778),
.B(n_1755),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1782),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1782),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1781),
.B(n_1702),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1809),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1791),
.A2(n_1702),
.B1(n_1698),
.B2(n_1711),
.Y(n_1855)
);

INVx4_ASAP7_75t_L g1856 ( 
.A(n_1804),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1781),
.B(n_1708),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1779),
.B(n_1758),
.Y(n_1858)
);

AO21x2_ASAP7_75t_L g1859 ( 
.A1(n_1780),
.A2(n_1761),
.B(n_1743),
.Y(n_1859)
);

INVx5_ASAP7_75t_L g1860 ( 
.A(n_1792),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1781),
.B(n_1705),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_SL g1862 ( 
.A1(n_1802),
.A2(n_1719),
.B1(n_1712),
.B2(n_1705),
.Y(n_1862)
);

INVx4_ASAP7_75t_L g1863 ( 
.A(n_1804),
.Y(n_1863)
);

AO21x2_ASAP7_75t_L g1864 ( 
.A1(n_1780),
.A2(n_1761),
.B(n_1757),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1817),
.A2(n_1698),
.B1(n_1726),
.B2(n_1699),
.Y(n_1865)
);

OAI211xp5_ASAP7_75t_SL g1866 ( 
.A1(n_1805),
.A2(n_1735),
.B(n_1775),
.C(n_1763),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1817),
.A2(n_1698),
.B1(n_1699),
.B2(n_1740),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1814),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1781),
.B(n_1765),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1788),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1859),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1850),
.B(n_1814),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1839),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1849),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1850),
.B(n_1814),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1826),
.B(n_1785),
.Y(n_1876)
);

NOR2x1_ASAP7_75t_SL g1877 ( 
.A(n_1838),
.B(n_1808),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1839),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1818),
.B(n_1787),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1842),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1845),
.B(n_1785),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1842),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1849),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1818),
.B(n_1787),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1848),
.A2(n_1802),
.B1(n_1797),
.B2(n_1809),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1846),
.B(n_1734),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1830),
.B(n_1796),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1849),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1830),
.B(n_1796),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1851),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1851),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1851),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1852),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1824),
.B(n_1792),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1852),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1852),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1858),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1824),
.B(n_1792),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1836),
.B(n_1805),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1832),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1821),
.B(n_1787),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1870),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1870),
.Y(n_1903)
);

INVx3_ASAP7_75t_SL g1904 ( 
.A(n_1838),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1823),
.B(n_1800),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1858),
.B(n_1807),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1821),
.B(n_1787),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1829),
.B(n_1815),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1823),
.B(n_1800),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1870),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1847),
.B(n_1789),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1822),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1829),
.B(n_1848),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1864),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1819),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1828),
.B(n_1813),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1819),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1847),
.B(n_1789),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1857),
.B(n_1815),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1904),
.B(n_1872),
.Y(n_1920)
);

INVxp67_ASAP7_75t_L g1921 ( 
.A(n_1899),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1873),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1904),
.B(n_1828),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1871),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1900),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1905),
.B(n_1847),
.Y(n_1926)
);

NAND2x2_ASAP7_75t_L g1927 ( 
.A(n_1913),
.B(n_1832),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1905),
.B(n_1847),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1904),
.B(n_1820),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1873),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1885),
.A2(n_1827),
.B1(n_1837),
.B2(n_1841),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1900),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1878),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1878),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1871),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1897),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1871),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1886),
.B(n_1752),
.Y(n_1938)
);

OAI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1881),
.A2(n_1837),
.B1(n_1831),
.B2(n_1843),
.Y(n_1939)
);

NOR4xp75_ASAP7_75t_L g1940 ( 
.A(n_1876),
.B(n_1843),
.C(n_1868),
.D(n_1831),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1880),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1880),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1872),
.B(n_1820),
.Y(n_1943)
);

AOI21xp33_ASAP7_75t_L g1944 ( 
.A1(n_1911),
.A2(n_1855),
.B(n_1866),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1882),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1875),
.B(n_1877),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1906),
.B(n_1857),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1882),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1909),
.B(n_1840),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1915),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1887),
.B(n_1834),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1915),
.Y(n_1952)
);

HB1xp67_ASAP7_75t_L g1953 ( 
.A(n_1914),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1909),
.B(n_1840),
.Y(n_1954)
);

INVxp67_ASAP7_75t_L g1955 ( 
.A(n_1911),
.Y(n_1955)
);

BUFx2_ASAP7_75t_L g1956 ( 
.A(n_1894),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1874),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1917),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1917),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1883),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1889),
.B(n_1834),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1875),
.B(n_1820),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1908),
.B(n_1752),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1883),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1877),
.B(n_1824),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1919),
.B(n_1835),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1932),
.B(n_1894),
.Y(n_1967)
);

NOR2x1_ASAP7_75t_L g1968 ( 
.A(n_1932),
.B(n_1774),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1921),
.B(n_1846),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1936),
.B(n_1918),
.Y(n_1970)
);

BUFx2_ASAP7_75t_L g1971 ( 
.A(n_1965),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1936),
.B(n_1918),
.Y(n_1972)
);

NAND4xp25_ASAP7_75t_L g1973 ( 
.A(n_1931),
.B(n_1794),
.C(n_1867),
.D(n_1862),
.Y(n_1973)
);

INVxp67_ASAP7_75t_L g1974 ( 
.A(n_1963),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1946),
.B(n_1894),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1949),
.B(n_1888),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1939),
.B(n_1854),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1933),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1965),
.B(n_1824),
.Y(n_1979)
);

INVxp67_ASAP7_75t_SL g1980 ( 
.A(n_1925),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1933),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1949),
.B(n_1888),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1924),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1934),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1924),
.Y(n_1985)
);

OAI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1927),
.A2(n_1865),
.B1(n_1794),
.B2(n_1854),
.C(n_1816),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1944),
.B(n_1951),
.Y(n_1987)
);

NOR2x1_ASAP7_75t_L g1988 ( 
.A(n_1965),
.B(n_1832),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1927),
.A2(n_1920),
.B1(n_1946),
.B2(n_1929),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1935),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1954),
.B(n_1947),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1934),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1920),
.B(n_1943),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1956),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1961),
.B(n_1861),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1943),
.B(n_1894),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1966),
.B(n_1861),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1935),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1922),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1962),
.B(n_1898),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1962),
.B(n_1898),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1938),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1923),
.B(n_1853),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1954),
.B(n_1890),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1930),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1994),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1968),
.A2(n_1929),
.B1(n_1923),
.B2(n_1956),
.Y(n_2007)
);

AOI222xp33_ASAP7_75t_L g2008 ( 
.A1(n_1977),
.A2(n_1940),
.B1(n_1955),
.B2(n_1898),
.C1(n_1953),
.C2(n_1792),
.Y(n_2008)
);

AOI32xp33_ASAP7_75t_L g2009 ( 
.A1(n_1987),
.A2(n_1898),
.A3(n_1820),
.B1(n_1928),
.B2(n_1926),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_SL g2010 ( 
.A1(n_1969),
.A2(n_1860),
.B1(n_1864),
.B2(n_1926),
.Y(n_2010)
);

OAI211xp5_ASAP7_75t_L g2011 ( 
.A1(n_1980),
.A2(n_1928),
.B(n_1860),
.C(n_1803),
.Y(n_2011)
);

OAI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1973),
.A2(n_1838),
.B1(n_1860),
.B2(n_1856),
.Y(n_2012)
);

AOI221xp5_ASAP7_75t_L g2013 ( 
.A1(n_1986),
.A2(n_1942),
.B1(n_1941),
.B2(n_1945),
.C(n_1948),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1971),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1971),
.Y(n_2015)
);

NAND2xp33_ASAP7_75t_SL g2016 ( 
.A(n_2002),
.B(n_1856),
.Y(n_2016)
);

O2A1O1Ixp33_ASAP7_75t_L g2017 ( 
.A1(n_1974),
.A2(n_1959),
.B(n_1950),
.C(n_1958),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1989),
.A2(n_1993),
.B1(n_2002),
.B2(n_1979),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1991),
.B(n_1699),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1993),
.A2(n_1988),
.B1(n_1975),
.B2(n_2001),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1994),
.A2(n_1991),
.B1(n_1972),
.B2(n_1970),
.Y(n_2021)
);

NOR3xp33_ASAP7_75t_L g2022 ( 
.A(n_1999),
.B(n_1964),
.C(n_1960),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_2005),
.B(n_1952),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1981),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_1970),
.Y(n_2025)
);

AOI21xp33_ASAP7_75t_L g2026 ( 
.A1(n_1972),
.A2(n_1967),
.B(n_1978),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1981),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1984),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1992),
.A2(n_1860),
.B(n_1937),
.Y(n_2029)
);

INVx3_ASAP7_75t_L g2030 ( 
.A(n_1967),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1983),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1983),
.Y(n_2032)
);

AOI22x1_ASAP7_75t_L g2033 ( 
.A1(n_1967),
.A2(n_1957),
.B1(n_1856),
.B2(n_1863),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1975),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_2019),
.B(n_1997),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2025),
.Y(n_2036)
);

NAND4xp25_ASAP7_75t_SL g2037 ( 
.A(n_2008),
.B(n_2001),
.C(n_2000),
.D(n_1996),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2006),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_2021),
.B(n_1995),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_2034),
.B(n_1996),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2024),
.Y(n_2041)
);

INVx1_ASAP7_75t_SL g2042 ( 
.A(n_2030),
.Y(n_2042)
);

OAI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_2007),
.A2(n_2003),
.B1(n_1860),
.B2(n_1838),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_SL g2044 ( 
.A1(n_2030),
.A2(n_2000),
.B1(n_1985),
.B2(n_1998),
.Y(n_2044)
);

NAND2x1p5_ASAP7_75t_L g2045 ( 
.A(n_2014),
.B(n_1604),
.Y(n_2045)
);

AOI32xp33_ASAP7_75t_L g2046 ( 
.A1(n_2012),
.A2(n_2004),
.A3(n_1982),
.B1(n_1976),
.B2(n_1985),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2015),
.B(n_1990),
.Y(n_2047)
);

OAI21xp33_ASAP7_75t_L g2048 ( 
.A1(n_2018),
.A2(n_1982),
.B(n_1976),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_2020),
.B(n_1879),
.Y(n_2049)
);

NAND2x1_ASAP7_75t_SL g2050 ( 
.A(n_2031),
.B(n_1990),
.Y(n_2050)
);

OAI222xp33_ASAP7_75t_L g2051 ( 
.A1(n_2009),
.A2(n_2004),
.B1(n_1838),
.B2(n_1860),
.C1(n_1863),
.C2(n_1856),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2026),
.B(n_1998),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_2027),
.Y(n_2053)
);

AOI221xp5_ASAP7_75t_L g2054 ( 
.A1(n_2013),
.A2(n_1964),
.B1(n_1960),
.B2(n_1957),
.C(n_1937),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_2023),
.B(n_1844),
.Y(n_2055)
);

OAI21xp5_ASAP7_75t_SL g2056 ( 
.A1(n_2011),
.A2(n_1816),
.B(n_1803),
.Y(n_2056)
);

NOR4xp25_ASAP7_75t_SL g2057 ( 
.A(n_2016),
.B(n_1902),
.C(n_1910),
.D(n_1895),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_2017),
.B(n_1853),
.Y(n_2058)
);

NAND3xp33_ASAP7_75t_L g2059 ( 
.A(n_2046),
.B(n_2036),
.C(n_2052),
.Y(n_2059)
);

OAI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_2056),
.A2(n_2011),
.B(n_2010),
.Y(n_2060)
);

O2A1O1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_2038),
.A2(n_2017),
.B(n_2028),
.C(n_2022),
.Y(n_2061)
);

INVx2_ASAP7_75t_SL g2062 ( 
.A(n_2050),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_2040),
.B(n_2032),
.Y(n_2063)
);

OAI21xp33_ASAP7_75t_SL g2064 ( 
.A1(n_2037),
.A2(n_2029),
.B(n_2010),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2042),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2042),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2047),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2048),
.B(n_2029),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2047),
.B(n_1874),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2041),
.Y(n_2070)
);

NAND3xp33_ASAP7_75t_L g2071 ( 
.A(n_2044),
.B(n_2033),
.C(n_1775),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2053),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_2043),
.B(n_1863),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2055),
.Y(n_2074)
);

NOR3xp33_ASAP7_75t_L g2075 ( 
.A(n_2059),
.B(n_2039),
.C(n_2035),
.Y(n_2075)
);

OAI221xp5_ASAP7_75t_L g2076 ( 
.A1(n_2060),
.A2(n_2058),
.B1(n_2054),
.B2(n_2045),
.C(n_2049),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2065),
.Y(n_2077)
);

OAI211xp5_ASAP7_75t_L g2078 ( 
.A1(n_2064),
.A2(n_2057),
.B(n_2051),
.C(n_2045),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2066),
.B(n_1879),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_2063),
.B(n_1884),
.Y(n_2080)
);

A2O1A1Ixp33_ASAP7_75t_L g2081 ( 
.A1(n_2061),
.A2(n_1868),
.B(n_1740),
.C(n_1907),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2067),
.Y(n_2082)
);

NOR2x1p5_ASAP7_75t_SL g2083 ( 
.A(n_2070),
.B(n_1892),
.Y(n_2083)
);

NAND4xp25_ASAP7_75t_L g2084 ( 
.A(n_2068),
.B(n_1863),
.C(n_1833),
.D(n_1689),
.Y(n_2084)
);

NAND3xp33_ASAP7_75t_SL g2085 ( 
.A(n_2068),
.B(n_1811),
.C(n_1833),
.Y(n_2085)
);

NAND3xp33_ASAP7_75t_L g2086 ( 
.A(n_2062),
.B(n_1689),
.C(n_1686),
.Y(n_2086)
);

NOR2x1_ASAP7_75t_L g2087 ( 
.A(n_2072),
.B(n_1890),
.Y(n_2087)
);

NAND4xp25_ASAP7_75t_L g2088 ( 
.A(n_2074),
.B(n_1684),
.C(n_1884),
.D(n_1916),
.Y(n_2088)
);

OAI211xp5_ASAP7_75t_SL g2089 ( 
.A1(n_2073),
.A2(n_1895),
.B(n_1902),
.C(n_1891),
.Y(n_2089)
);

AOI21xp5_ASAP7_75t_L g2090 ( 
.A1(n_2071),
.A2(n_1892),
.B(n_1893),
.Y(n_2090)
);

AOI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_2075),
.A2(n_2078),
.B(n_2076),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_R g2092 ( 
.A(n_2077),
.B(n_2069),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2079),
.Y(n_2093)
);

NOR3xp33_ASAP7_75t_SL g2094 ( 
.A(n_2085),
.B(n_2069),
.C(n_1910),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2083),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_R g2096 ( 
.A(n_2082),
.B(n_1604),
.Y(n_2096)
);

NAND3xp33_ASAP7_75t_L g2097 ( 
.A(n_2081),
.B(n_2086),
.C(n_2089),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2080),
.B(n_1901),
.Y(n_2098)
);

AND4x1_ASAP7_75t_L g2099 ( 
.A(n_2091),
.B(n_2087),
.C(n_2090),
.D(n_2084),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2093),
.A2(n_2088),
.B1(n_1719),
.B2(n_1916),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2095),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2092),
.Y(n_2102)
);

AOI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_2097),
.A2(n_1912),
.B(n_1893),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2098),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_2096),
.A2(n_1719),
.B1(n_2094),
.B2(n_1733),
.Y(n_2105)
);

AOI222xp33_ASAP7_75t_L g2106 ( 
.A1(n_2097),
.A2(n_1903),
.B1(n_1896),
.B2(n_1891),
.C1(n_1901),
.C2(n_1907),
.Y(n_2106)
);

AND2x4_ASAP7_75t_L g2107 ( 
.A(n_2102),
.B(n_1869),
.Y(n_2107)
);

NOR2x1_ASAP7_75t_L g2108 ( 
.A(n_2101),
.B(n_1896),
.Y(n_2108)
);

NOR3xp33_ASAP7_75t_L g2109 ( 
.A(n_2104),
.B(n_1704),
.C(n_1759),
.Y(n_2109)
);

OAI221xp5_ASAP7_75t_SL g2110 ( 
.A1(n_2105),
.A2(n_2099),
.B1(n_2100),
.B2(n_2103),
.C(n_2106),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2102),
.B(n_1869),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2102),
.B(n_1912),
.Y(n_2112)
);

XNOR2xp5_ASAP7_75t_L g2113 ( 
.A(n_2099),
.B(n_1682),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_2110),
.B(n_1903),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2107),
.B(n_1822),
.Y(n_2115)
);

OAI321xp33_ASAP7_75t_L g2116 ( 
.A1(n_2112),
.A2(n_1604),
.A3(n_1635),
.B1(n_1645),
.B2(n_1733),
.C(n_1681),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2114),
.B(n_2111),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2117),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2118),
.Y(n_2119)
);

INVx2_ASAP7_75t_SL g2120 ( 
.A(n_2118),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_SL g2121 ( 
.A1(n_2119),
.A2(n_2113),
.B1(n_2108),
.B2(n_2115),
.Y(n_2121)
);

OAI22xp5_ASAP7_75t_SL g2122 ( 
.A1(n_2120),
.A2(n_2109),
.B1(n_2116),
.B2(n_1635),
.Y(n_2122)
);

INVxp67_ASAP7_75t_L g2123 ( 
.A(n_2121),
.Y(n_2123)
);

AOI21x1_ASAP7_75t_L g2124 ( 
.A1(n_2122),
.A2(n_1825),
.B(n_1822),
.Y(n_2124)
);

XNOR2xp5_ASAP7_75t_L g2125 ( 
.A(n_2123),
.B(n_2124),
.Y(n_2125)
);

OAI22xp5_ASAP7_75t_SL g2126 ( 
.A1(n_2125),
.A2(n_1635),
.B1(n_1645),
.B2(n_1677),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_2126),
.A2(n_1635),
.B(n_1645),
.Y(n_2127)
);

OAI221xp5_ASAP7_75t_R g2128 ( 
.A1(n_2127),
.A2(n_1677),
.B1(n_1864),
.B2(n_1859),
.C(n_1675),
.Y(n_2128)
);

AOI211xp5_ASAP7_75t_L g2129 ( 
.A1(n_2128),
.A2(n_1635),
.B(n_1645),
.C(n_1654),
.Y(n_2129)
);


endmodule