module real_jpeg_9131_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_295, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_295;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_243;
wire n_105;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_216;
wire n_167;
wire n_179;
wire n_133;
wire n_202;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_1),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_2),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_2),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_2),
.A2(n_12),
.B(n_34),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_7),
.A2(n_33),
.B(n_44),
.C(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_33),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_9),
.A2(n_28),
.B1(n_36),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_9),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_111),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_111),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_111),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_10),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_128),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_128),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_10),
.A2(n_28),
.B1(n_36),
.B2(n_128),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_12),
.A2(n_46),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_12),
.B(n_46),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_12),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_12),
.A2(n_83),
.B1(n_86),
.B2(n_146),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_12),
.A2(n_33),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_12),
.B(n_33),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_12),
.B(n_193),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_12),
.A2(n_28),
.B1(n_36),
.B2(n_148),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_13),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_137),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_137),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_13),
.A2(n_28),
.B1(n_36),
.B2(n_137),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_14),
.A2(n_28),
.B1(n_36),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_14),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_93),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_93),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_93),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_15),
.A2(n_28),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_15),
.A2(n_39),
.B1(n_46),
.B2(n_47),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_15),
.A2(n_39),
.B1(n_60),
.B2(n_61),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_16),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_17),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_17),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_17),
.A2(n_37),
.B1(n_60),
.B2(n_61),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_17),
.A2(n_37),
.B1(n_46),
.B2(n_47),
.Y(n_225)
);

HAxp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_117),
.CON(n_18),
.SN(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_115),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_94),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_21),
.B(n_94),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_79),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_66),
.B2(n_67),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_40),
.B2(n_41),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_27),
.A2(n_32),
.B1(n_35),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_27),
.A2(n_32),
.B1(n_92),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_27),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_27),
.A2(n_32),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_27),
.A2(n_32),
.B1(n_110),
.B2(n_244),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_30),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_28),
.A2(n_30),
.B(n_148),
.C(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_32),
.Y(n_193)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_54),
.B1(n_55),
.B2(n_65),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_49),
.B2(n_52),
.Y(n_42)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_43),
.A2(n_45),
.B1(n_71),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_43),
.A2(n_45),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_43),
.A2(n_45),
.B1(n_173),
.B2(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_43),
.A2(n_45),
.B1(n_189),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_43),
.A2(n_45),
.B1(n_228),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_43),
.A2(n_45),
.B1(n_114),
.B2(n_240),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_44),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_45),
.B(n_148),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_46),
.B(n_48),
.Y(n_177)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_47),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_59),
.B(n_63),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_59),
.B1(n_75),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_56),
.A2(n_59),
.B1(n_89),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_56),
.A2(n_59),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_56),
.A2(n_59),
.B1(n_136),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_56),
.A2(n_59),
.B1(n_161),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_56),
.A2(n_59),
.B1(n_169),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_56),
.A2(n_59),
.B1(n_107),
.B2(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_59),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_60),
.B(n_62),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_60),
.B(n_152),
.Y(n_151)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_61),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_68),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_76),
.A2(n_78),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_90),
.B(n_91),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_81),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_90),
.B1(n_91),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_82),
.A2(n_88),
.B1(n_90),
.B2(n_275),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B(n_87),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_86),
.B1(n_87),
.B2(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_83),
.A2(n_86),
.B1(n_127),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_83),
.A2(n_86),
.B1(n_130),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_83),
.A2(n_86),
.B1(n_163),
.B2(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_83),
.A2(n_86),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_83),
.A2(n_86),
.B1(n_105),
.B2(n_216),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_85),
.B1(n_126),
.B2(n_129),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_84),
.A2(n_85),
.B1(n_181),
.B2(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_148),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_88),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_101),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_95),
.Y(n_280)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_101),
.A2(n_102),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.C(n_112),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_103),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_104),
.B(n_106),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI321xp33_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_269),
.A3(n_281),
.B1(n_287),
.B2(n_292),
.C(n_295),
.Y(n_117)
);

NOR3xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_234),
.C(n_265),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_205),
.B(n_233),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_183),
.B(n_204),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_165),
.B(n_182),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_155),
.B(n_164),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_143),
.B(n_154),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_131),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_138),
.B2(n_142),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_132),
.B(n_142),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_135),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_138),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_149),
.B(n_153),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_157),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_160),
.C(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_167),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.CI(n_174),
.CON(n_167),
.SN(n_167)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_172),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_179),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_185),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_197),
.B2(n_198),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_200),
.C(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_190),
.B1(n_191),
.B2(n_196),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_188),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_194),
.C(n_196),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_199),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_200),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_206),
.B(n_207),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_220),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_209),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_209),
.B(n_219),
.C(n_220),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_214),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_217),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_226),
.C(n_229),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_232),
.Y(n_243)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_235),
.A2(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_252),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_236),
.B(n_252),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_247),
.C(n_251),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_246),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_241),
.B1(n_242),
.B2(n_245),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_SL g263 ( 
.A(n_241),
.B(n_245),
.C(n_246),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_251),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_249),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_263),
.B2(n_264),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_256),
.C(n_264),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_260),
.C(n_262),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_259),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_267),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_277),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_274),
.C(n_276),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_274),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_288),
.B(n_291),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_284),
.Y(n_291)
);


endmodule