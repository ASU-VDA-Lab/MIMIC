module real_jpeg_6570_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_1),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_2),
.Y(n_111)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_2),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_3),
.A2(n_45),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_45),
.B1(n_115),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_3),
.A2(n_45),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_3),
.B(n_148),
.C(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_3),
.B(n_247),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_3),
.A2(n_254),
.B(n_256),
.C(n_257),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_3),
.B(n_267),
.C(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_3),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_3),
.B(n_213),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_3),
.B(n_24),
.Y(n_293)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_4),
.Y(n_63)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_5),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_5),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_5),
.Y(n_280)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_6),
.Y(n_236)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_9),
.Y(n_128)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_9),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_10),
.A2(n_49),
.B1(n_53),
.B2(n_56),
.Y(n_48)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_10),
.A2(n_41),
.B1(n_56),
.B2(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_10),
.A2(n_56),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_10),
.A2(n_56),
.B1(n_74),
.B2(n_186),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_83),
.B1(n_87),
.B2(n_90),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_90),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_11),
.A2(n_90),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_90),
.B1(n_161),
.B2(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_12),
.Y(n_97)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_364),
.B(n_366),
.Y(n_17)
);

AO21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_136),
.B(n_363),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_131),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_20),
.B(n_131),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_119),
.C(n_130),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_21),
.A2(n_22),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_47),
.C(n_91),
.Y(n_22)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_23),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_23),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_23),
.B(n_201),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_23),
.A2(n_178),
.B1(n_179),
.B2(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_23),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_23),
.A2(n_220),
.B1(n_250),
.B2(n_260),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_23),
.B(n_170),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_23),
.A2(n_220),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_23),
.A2(n_178),
.B(n_216),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_23),
.A2(n_220),
.B1(n_348),
.B2(n_349),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_23),
.A2(n_220),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

OA21x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_34),
.B(n_43),
.Y(n_23)
);

NOR2x1_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_24),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_30),
.Y(n_147)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_35)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_36),
.Y(n_133)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_45),
.A2(n_71),
.B(n_74),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_47),
.A2(n_91),
.B1(n_92),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_47),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_57),
.B1(n_70),
.B2(n_82),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_48),
.A2(n_57),
.B1(n_70),
.B2(n_145),
.Y(n_341)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AO21x1_ASAP7_75t_L g130 ( 
.A1(n_57),
.A2(n_70),
.B(n_82),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AO21x2_ASAP7_75t_SL g144 ( 
.A1(n_58),
.A2(n_70),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_70),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_59)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_60),
.Y(n_255)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_70),
.Y(n_247)
);

OA22x2_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_79),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_89),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_91),
.A2(n_92),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_92),
.B(n_220),
.C(n_341),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_102),
.B(n_113),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_93),
.B(n_102),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_93),
.A2(n_102),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_93),
.Y(n_211)
);

NAND2x1_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_102),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_101),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_97),
.Y(n_268)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B1(n_108),
.B2(n_112),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_103),
.B(n_277),
.Y(n_276)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_105),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_113),
.Y(n_212)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g269 ( 
.A(n_116),
.Y(n_269)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_119),
.B(n_130),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_129),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_122),
.B1(n_129),
.B2(n_132),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g365 ( 
.A1(n_121),
.A2(n_129),
.B(n_132),
.Y(n_365)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_131),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_131),
.B(n_365),
.Y(n_367)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_357),
.B(n_362),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_335),
.B(n_354),
.Y(n_137)
);

OAI211xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_240),
.B(n_329),
.C(n_334),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_222),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g329 ( 
.A1(n_140),
.A2(n_222),
.B(n_330),
.C(n_333),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_204),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_141),
.B(n_204),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_177),
.C(n_189),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_142),
.B(n_177),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_149),
.B1(n_175),
.B2(n_176),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_143),
.B(n_190),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_143),
.A2(n_175),
.B1(n_229),
.B2(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_144),
.B(n_210),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_144),
.A2(n_203),
.B(n_220),
.C(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_144),
.A2(n_170),
.B1(n_201),
.B2(n_226),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_144),
.A2(n_201),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_149),
.A2(n_200),
.B(n_202),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_170),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_150),
.A2(n_170),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_150),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_157),
.B1(n_163),
.B2(n_167),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_155),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_157),
.B1(n_192),
.B2(n_198),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_153),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_167),
.B(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_170),
.B(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_170),
.A2(n_226),
.B1(n_246),
.B2(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_170),
.A2(n_226),
.B1(n_264),
.B2(n_265),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_170),
.A2(n_226),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_L g297 ( 
.A1(n_170),
.A2(n_201),
.B(n_252),
.C(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_170),
.B(n_201),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_170),
.A2(n_191),
.B1(n_226),
.B2(n_320),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_188),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_182),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_193),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_210)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_189),
.B(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_200),
.B(n_202),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_191),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_209),
.B(n_214),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_201),
.B(n_237),
.C(n_292),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AND3x1_ASAP7_75t_L g322 ( 
.A(n_203),
.B(n_299),
.C(n_323),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_221),
.Y(n_204)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_208),
.B(n_215),
.C(n_221),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

FAx1_ASAP7_75t_L g337 ( 
.A(n_214),
.B(n_338),
.CI(n_343),
.CON(n_337),
.SN(n_337)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_220),
.B(n_349),
.C(n_353),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_238),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_223),
.B(n_238),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.C(n_228),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_224),
.B(n_225),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_246),
.C(n_248),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_226),
.B(n_289),
.C(n_296),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_228),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_237),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_230),
.A2(n_231),
.B1(n_237),
.B2(n_248),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_237),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_248),
.B1(n_253),
.B2(n_259),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_237),
.B(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_237),
.A2(n_248),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_237),
.B(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_311),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_301),
.B(n_310),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_287),
.B(n_300),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_261),
.B(n_286),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_245),
.B(n_249),
.Y(n_286)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_246),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_248),
.B(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_260),
.Y(n_249)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_253),
.Y(n_259)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_273),
.B(n_285),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_270),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_283),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_281),
.Y(n_274)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_297),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_297),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_307),
.C(n_308),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_324),
.Y(n_311)
);

NOR2x1_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_314),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_317),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_321),
.B2(n_322),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_321),
.C(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_324),
.A2(n_331),
.B(n_332),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_327),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_345),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_344),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_337),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_344),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_337),
.B(n_346),
.Y(n_356)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_345),
.A2(n_355),
.B(n_356),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_353),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_361),
.Y(n_362)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_367),
.Y(n_366)
);


endmodule