module real_jpeg_33016_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g12 ( 
.A(n_0),
.B(n_1),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_4),
.B(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx2_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

AOI322xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_10),
.A3(n_11),
.B1(n_15),
.B2(n_17),
.C1(n_22),
.C2(n_29),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NAND2xp33_ASAP7_75t_SL g27 ( 
.A(n_10),
.B(n_20),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_10),
.B(n_21),
.Y(n_28)
);

AND2x4_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

NAND3xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_27),
.C(n_28),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);


endmodule