module real_jpeg_7497_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_61),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_1),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_1),
.B(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_1),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_1),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_1),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_2),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_2),
.B(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_2),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_2),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_2),
.B(n_183),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_2),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_2),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_3),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_3),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_3),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_3),
.B(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_4),
.Y(n_193)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_4),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_5),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_5),
.B(n_202),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_5),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g301 ( 
.A(n_5),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_5),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_5),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_5),
.B(n_401),
.Y(n_400)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_7),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_7),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_7),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_7),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_7),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_7),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_7),
.B(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_8),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_8),
.Y(n_158)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_9),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_9),
.B(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_9),
.B(n_121),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_9),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_9),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_9),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_9),
.B(n_89),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_12),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_12),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_12),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_12),
.B(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_12),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_12),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_12),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_12),
.B(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_13),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_13),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_13),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_13),
.Y(n_332)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_14),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_15),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_16),
.Y(n_165)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_16),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_16),
.Y(n_433)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_17),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_17),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_17),
.B(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_504),
.B(n_507),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_72),
.B(n_105),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_21),
.B(n_72),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.C(n_35),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_24),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_24),
.A2(n_35),
.B1(n_49),
.B2(n_58),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_24),
.B(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_28),
.Y(n_118)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_29),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_29),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_30),
.A2(n_31),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_30),
.A2(n_31),
.B1(n_337),
.B2(n_343),
.Y(n_336)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_31),
.B(n_338),
.C(n_342),
.Y(n_485)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_35),
.A2(n_58),
.B1(n_63),
.B2(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_35),
.A2(n_58),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_35),
.B(n_146),
.C(n_150),
.Y(n_254)
);

OR2x2_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_36),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_38),
.Y(n_277)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_39),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_39),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_64),
.Y(n_63)
);

OR2x2_ASAP7_75t_SL g77 ( 
.A(n_40),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_40),
.B(n_331),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_44),
.A2(n_45),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_44),
.A2(n_45),
.B1(n_355),
.B2(n_356),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_44),
.B(n_351),
.C(n_356),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_45),
.B(n_313),
.C(n_318),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_46),
.Y(n_168)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_47),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_49),
.B(n_229),
.C(n_232),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_50),
.A2(n_51),
.B1(n_76),
.B2(n_77),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_63),
.C(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.C(n_62),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_55),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_63),
.C(n_69),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_62),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_99),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_63),
.B(n_117),
.C(n_120),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_63),
.A2(n_99),
.B1(n_480),
.B2(n_481),
.Y(n_479)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_67),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_67),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_67),
.Y(n_378)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_68),
.Y(n_253)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_68),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_70),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_69),
.A2(n_70),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_69),
.B(n_191),
.C(n_296),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_100),
.C(n_101),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_73),
.B(n_501),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_87),
.C(n_96),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_74),
.B(n_492),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_83),
.C(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_76),
.A2(n_77),
.B1(n_130),
.B2(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_76),
.A2(n_77),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_77),
.B(n_127),
.C(n_130),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_77),
.B(n_191),
.C(n_330),
.Y(n_484)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_79),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_83),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_87),
.B(n_96),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.C(n_95),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_88),
.A2(n_91),
.B1(n_92),
.B2(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_88),
.Y(n_475)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_91),
.A2(n_92),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_92),
.B(n_135),
.C(n_238),
.Y(n_318)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_94),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_95),
.B(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_100),
.B(n_101),
.Y(n_501)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_499),
.B(n_503),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_467),
.B(n_496),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_357),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_285),
.B(n_320),
.C(n_321),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_255),
.B(n_284),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_111),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_221),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_112),
.B(n_221),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_169),
.C(n_205),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_113),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_142),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_114),
.B(n_143),
.C(n_151),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_126),
.C(n_133),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_115),
.B(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_124),
.B(n_172),
.Y(n_425)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_126),
.A2(n_133),
.B1(n_134),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_126),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_127),
.B(n_263),
.Y(n_262)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_130),
.Y(n_264)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_135),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_135),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_240),
.Y(n_278)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_151),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_147),
.B(n_191),
.Y(n_373)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_148),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_153),
.B(n_155),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_152),
.B(n_160),
.C(n_166),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_167),
.B(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_169),
.B(n_205),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_186),
.C(n_188),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_170),
.A2(n_186),
.B1(n_187),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_175),
.C(n_180),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_172),
.B(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_179),
.B1(n_180),
.B2(n_185),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_179),
.A2(n_180),
.B1(n_300),
.B2(n_304),
.Y(n_299)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_180),
.B(n_238),
.C(n_301),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_188),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_194),
.C(n_200),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_189),
.A2(n_190),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_191),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_191),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_191),
.A2(n_293),
.B1(n_330),
.B2(n_333),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g368 ( 
.A(n_193),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_194),
.A2(n_195),
.B1(n_200),
.B2(n_201),
.Y(n_455)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_199),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_199),
.Y(n_429)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_220),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_208),
.C(n_220),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_216),
.C(n_219),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_214),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_214),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_216),
.A2(n_338),
.B1(n_341),
.B2(n_342),
.Y(n_337)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_216),
.Y(n_342)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_222),
.B(n_224),
.C(n_241),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_241),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_234),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_226),
.B(n_227),
.C(n_234),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_237),
.A2(n_238),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_237),
.A2(n_238),
.B1(n_365),
.B2(n_366),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_238),
.B(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_247),
.B(n_249),
.C(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_254),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_282),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_256),
.B(n_282),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.C(n_279),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_257),
.A2(n_258),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_261),
.B(n_279),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_278),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_262),
.B(n_449),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_265),
.B(n_278),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_271),
.C(n_274),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_266),
.A2(n_267),
.B1(n_274),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_271),
.B(n_385),
.Y(n_384)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_273),
.Y(n_410)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_274),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_275),
.B(n_377),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_275),
.B(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_286),
.B(n_322),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_288),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_323),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_288),
.B(n_323),
.Y(n_466)
);

FAx1_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_305),
.CI(n_319),
.CON(n_288),
.SN(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_299),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_292),
.C(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_300),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_301),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_308),
.C(n_310),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_318),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_324),
.B(n_326),
.C(n_344),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_344),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_334),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_327),
.B(n_335),
.C(n_336),
.Y(n_476)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_330),
.Y(n_333)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_337),
.Y(n_343)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_338),
.Y(n_341)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_345),
.B(n_349),
.C(n_350),
.Y(n_486)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

AO22x1_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_355),
.Y(n_356)
);

OAI31xp33_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_463),
.A3(n_464),
.B(n_466),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_457),
.B(n_462),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_444),
.B(n_456),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_404),
.B(n_443),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_387),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_362),
.B(n_387),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_374),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_363),
.B(n_375),
.C(n_384),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_369),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_364),
.B(n_370),
.C(n_373),
.Y(n_452)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_373),
.Y(n_369)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_384),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.C(n_382),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_376),
.B(n_389),
.Y(n_388)
);

INVx11_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_379),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.Y(n_389)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.C(n_403),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_388),
.B(n_440),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_390),
.A2(n_391),
.B1(n_403),
.B2(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_399),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_392),
.A2(n_393),
.B1(n_399),
.B2(n_400),
.Y(n_413)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_405),
.A2(n_437),
.B(n_442),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_423),
.B(n_436),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_414),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_414),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_413),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_409),
.B(n_411),
.C(n_413),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_420),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_415),
.A2(n_416),
.B1(n_420),
.B2(n_421),
.Y(n_434)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_421),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_430),
.B(n_435),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx8_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_434),
.Y(n_435)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_439),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_445),
.B(n_446),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_452),
.C(n_453),
.Y(n_461)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_458),
.B(n_461),
.Y(n_462)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_459),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_493),
.Y(n_467)
);

OAI21xp33_ASAP7_75t_L g496 ( 
.A1(n_468),
.A2(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_487),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_487),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_477),
.C(n_486),
.Y(n_469)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_470),
.B(n_477),
.CI(n_486),
.CON(n_495),
.SN(n_495)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_476),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_473),
.C(n_476),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_482),
.B2(n_483),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_484),
.C(n_485),
.Y(n_490)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_490),
.C(n_491),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_495),
.Y(n_497)
);

BUFx24_ASAP7_75t_SL g510 ( 
.A(n_495),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_502),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_500),
.B(n_502),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx13_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx8_ASAP7_75t_L g508 ( 
.A(n_506),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_509),
.Y(n_507)
);


endmodule