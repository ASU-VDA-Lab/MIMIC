module fake_netlist_1_1878_n_17 (n_1, n_2, n_0, n_17);
input n_1;
input n_2;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
AOI21x1_ASAP7_75t_L g3 ( .A1(n_0), .A2(n_2), .B(n_1), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
NAND2xp5_ASAP7_75t_SL g5 ( .A(n_1), .B(n_2), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
AOI21xp5_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_5), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_0), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
INVx1_ASAP7_75t_SL g11 ( .A(n_8), .Y(n_11) );
NOR2x1_ASAP7_75t_SL g12 ( .A(n_10), .B(n_3), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_10), .B(n_2), .Y(n_13) );
OAI211xp5_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_11), .B(n_1), .C(n_2), .Y(n_14) );
OR2x2_ASAP7_75t_L g15 ( .A(n_12), .B(n_11), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
AOI222xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_12), .C1(n_14), .C2(n_10), .Y(n_17) );
endmodule