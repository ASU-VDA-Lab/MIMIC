module fake_jpeg_276_n_161 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_55),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_62),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_1),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_48),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_42),
.B1(n_49),
.B2(n_50),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_73),
.B1(n_50),
.B2(n_49),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_51),
.B1(n_52),
.B2(n_42),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_49),
.B1(n_51),
.B2(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_47),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_76),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_44),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_46),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_83),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_65),
.B(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_39),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_1),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_45),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_91),
.Y(n_98)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_54),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_65),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_65),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_102),
.C(n_84),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_11),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_68),
.B1(n_5),
.B2(n_7),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_18),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_10),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_118),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_107),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_122),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_88),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_108),
.C(n_99),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_12),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_126),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_14),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_88),
.B(n_16),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_93),
.B(n_19),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_136),
.C(n_137),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g147 ( 
.A(n_134),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_15),
.B1(n_20),
.B2(n_21),
.Y(n_135)
);

NAND2x1p5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_110),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_143),
.B(n_145),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_113),
.C(n_112),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_129),
.CI(n_135),
.CON(n_150),
.SN(n_150)
);

AOI322xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_111),
.A3(n_114),
.B1(n_31),
.B2(n_32),
.C1(n_33),
.C2(n_35),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_138),
.B(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_151),
.B1(n_138),
.B2(n_152),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_132),
.C(n_137),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_154),
.B1(n_130),
.B2(n_150),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_153),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_139),
.B1(n_131),
.B2(n_147),
.Y(n_158)
);

AOI21x1_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_142),
.B(n_127),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_24),
.B(n_25),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_37),
.Y(n_161)
);


endmodule