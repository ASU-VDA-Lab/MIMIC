module fake_jpeg_28976_n_169 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_31),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_34),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_1),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_94),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_70),
.B1(n_60),
.B2(n_64),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_95),
.B(n_29),
.C(n_48),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_89),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_73),
.B(n_62),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_86),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_62),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_59),
.B1(n_67),
.B2(n_65),
.Y(n_90)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_71),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_59),
.B1(n_58),
.B2(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_114),
.B1(n_3),
.B2(n_5),
.Y(n_120)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_106),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_107),
.Y(n_127)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_68),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_66),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_3),
.B(n_4),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_61),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_83),
.A2(n_63),
.B1(n_57),
.B2(n_52),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_83),
.B(n_51),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_124),
.B(n_11),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_83),
.B1(n_4),
.B2(n_5),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_126),
.B1(n_135),
.B2(n_13),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_6),
.B(n_7),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_14),
.C(n_42),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_87),
.B(n_7),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_98),
.B(n_100),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_130),
.C(n_132),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_27),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_9),
.B(n_10),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_47),
.B1(n_28),
.B2(n_30),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_11),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_140),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_141),
.C(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_12),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_33),
.C(n_40),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_143),
.C(n_147),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_25),
.C(n_39),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_23),
.B(n_38),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_13),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_149),
.C(n_144),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_22),
.C(n_35),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_150),
.C(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_37),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_135),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_125),
.A3(n_129),
.B1(n_131),
.B2(n_134),
.C1(n_137),
.C2(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_155),
.B(n_157),
.Y(n_161)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_162),
.Y(n_163)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_164),
.C(n_156),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_160),
.B(n_161),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_153),
.C(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_150),
.Y(n_169)
);


endmodule