module fake_netlist_1_3633_n_34 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_34);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_34;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_30;
wire n_26;
wire n_13;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_6), .B(n_4), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
NAND2xp5_ASAP7_75t_SL g17 ( .A(n_12), .B(n_0), .Y(n_17) );
AND2x6_ASAP7_75t_L g18 ( .A(n_12), .B(n_7), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_18), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_12), .B(n_13), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
AND2x2_ASAP7_75t_SL g24 ( .A(n_22), .B(n_11), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
NAND2xp5_ASAP7_75t_SL g26 ( .A(n_24), .B(n_19), .Y(n_26) );
OAI211xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_15), .B(n_14), .C(n_11), .Y(n_27) );
AO22x2_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_23), .B1(n_24), .B2(n_3), .Y(n_28) );
OAI21xp33_ASAP7_75t_SL g29 ( .A1(n_28), .A2(n_19), .B(n_18), .Y(n_29) );
NOR2x1_ASAP7_75t_L g30 ( .A(n_27), .B(n_11), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
OAI22xp5_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_16), .B1(n_18), .B2(n_3), .Y(n_32) );
OAI22xp5_ASAP7_75t_SL g33 ( .A1(n_31), .A2(n_0), .B1(n_2), .B2(n_8), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_32), .B1(n_2), .B2(n_10), .Y(n_34) );
endmodule