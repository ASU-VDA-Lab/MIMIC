module fake_jpeg_20292_n_154 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_20),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_6),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_78),
.Y(n_90)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_59),
.B1(n_50),
.B2(n_57),
.Y(n_84)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_2),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_69),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_80),
.A2(n_57),
.B1(n_71),
.B2(n_73),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_89),
.B1(n_94),
.B2(n_64),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_60),
.C(n_66),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_87),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_66),
.C(n_61),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_78),
.A2(n_48),
.B1(n_56),
.B2(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_49),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_52),
.B1(n_55),
.B2(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_67),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_58),
.B1(n_61),
.B2(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_86),
.B1(n_92),
.B2(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_104),
.Y(n_113)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_75),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_74),
.C(n_72),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_5),
.Y(n_130)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_120),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_115),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_2),
.Y(n_117)
);

OR2x2_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_119),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_58),
.B(n_4),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_107),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_122),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_133),
.B1(n_9),
.B2(n_121),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_118),
.B1(n_109),
.B2(n_122),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_126),
.A2(n_109),
.B1(n_23),
.B2(n_24),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_131),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_28),
.A3(n_44),
.B1(n_10),
.B2(n_17),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_29),
.B1(n_42),
.B2(n_18),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_132),
.A2(n_129),
.B1(n_134),
.B2(n_108),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_7),
.B1(n_9),
.B2(n_21),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_22),
.B(n_26),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_27),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_140),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_141),
.B1(n_142),
.B2(n_126),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_132),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_125),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_136),
.B1(n_33),
.B2(n_35),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_154)
);


endmodule