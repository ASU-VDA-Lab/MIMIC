module fake_jpeg_11699_n_140 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_8),
.B(n_24),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_60),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_72),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_71),
.B1(n_54),
.B2(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_73),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_55),
.B1(n_61),
.B2(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_23),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_72),
.B(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_56),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_50),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_76),
.A2(n_64),
.B1(n_54),
.B2(n_48),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_0),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_100),
.Y(n_117)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_63),
.B(n_60),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_31),
.B(n_44),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_1),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_63),
.C(n_30),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_12),
.C(n_16),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_2),
.C(n_4),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_113),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_115),
.B(n_34),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_92),
.C(n_88),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_107),
.C(n_35),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_28),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_86),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_5),
.B1(n_9),
.B2(n_11),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_101),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_116),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_46),
.B(n_21),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_20),
.Y(n_116)
);

NOR4xp25_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_22),
.C(n_32),
.D(n_33),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_119),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_123),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_95),
.B1(n_36),
.B2(n_37),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_126),
.B1(n_114),
.B2(n_111),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_43),
.C(n_40),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_127),
.C(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_132),
.C(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

OAI21x1_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_117),
.B(n_121),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_134),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_135),
.B(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_125),
.Y(n_140)
);


endmodule