module real_aes_8339_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_516;
wire n_177;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
INVx1_ASAP7_75t_L g529 ( .A(n_1), .Y(n_529) );
INVx1_ASAP7_75t_L g147 ( .A(n_2), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_3), .A2(n_38), .B1(n_172), .B2(n_475), .Y(n_498) );
AOI21xp33_ASAP7_75t_L g179 ( .A1(n_4), .A2(n_163), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_5), .B(n_161), .Y(n_541) );
AND2x6_ASAP7_75t_L g140 ( .A(n_6), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_7), .A2(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_8), .B(n_39), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_8), .B(n_39), .Y(n_437) );
INVx1_ASAP7_75t_L g185 ( .A(n_9), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_10), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g132 ( .A(n_11), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_12), .B(n_153), .Y(n_484) );
INVx1_ASAP7_75t_L g256 ( .A(n_13), .Y(n_256) );
INVx1_ASAP7_75t_L g523 ( .A(n_14), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_15), .B(n_128), .Y(n_512) );
AO32x2_ASAP7_75t_L g496 ( .A1(n_16), .A2(n_127), .A3(n_161), .B1(n_477), .B2(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_17), .B(n_172), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_18), .B(n_168), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_19), .B(n_128), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_20), .A2(n_50), .B1(n_172), .B2(n_475), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_21), .B(n_163), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_22), .A2(n_97), .B1(n_729), .B2(n_730), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_22), .Y(n_730) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_23), .A2(n_75), .B1(n_153), .B2(n_172), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_24), .B(n_172), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_25), .B(n_175), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_26), .A2(n_254), .B(n_255), .C(n_257), .Y(n_253) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_28), .B(n_158), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_29), .B(n_151), .Y(n_150) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_30), .A2(n_87), .B1(n_118), .B2(n_119), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_30), .Y(n_118) );
INVx1_ASAP7_75t_L g200 ( .A(n_31), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_32), .B(n_158), .Y(n_468) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_33), .A2(n_442), .B1(n_727), .B2(n_728), .C1(n_731), .C2(n_733), .Y(n_441) );
INVx2_ASAP7_75t_L g138 ( .A(n_34), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_35), .B(n_172), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_36), .B(n_158), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_37), .A2(n_140), .B(n_143), .C(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g198 ( .A(n_40), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_41), .B(n_151), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_42), .A2(n_102), .B1(n_103), .B2(n_110), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_43), .B(n_172), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_44), .A2(n_85), .B1(n_220), .B2(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_45), .B(n_172), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_46), .B(n_172), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_47), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_48), .B(n_528), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_49), .B(n_163), .Y(n_244) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_51), .A2(n_60), .B1(n_153), .B2(n_172), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_52), .A2(n_143), .B1(n_153), .B2(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_53), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_54), .B(n_172), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_55), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_56), .B(n_172), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_57), .A2(n_171), .B(n_183), .C(n_184), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_58), .Y(n_233) );
INVx1_ASAP7_75t_L g181 ( .A(n_59), .Y(n_181) );
INVx1_ASAP7_75t_L g141 ( .A(n_61), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_62), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_63), .B(n_172), .Y(n_530) );
INVx1_ASAP7_75t_L g131 ( .A(n_64), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_65), .Y(n_114) );
AO32x2_ASAP7_75t_L g472 ( .A1(n_66), .A2(n_161), .A3(n_236), .B1(n_473), .B2(n_477), .Y(n_472) );
INVx1_ASAP7_75t_L g548 ( .A(n_67), .Y(n_548) );
INVx1_ASAP7_75t_L g463 ( .A(n_68), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_SL g167 ( .A1(n_69), .A2(n_168), .B(n_169), .C(n_171), .Y(n_167) );
INVxp67_ASAP7_75t_L g170 ( .A(n_70), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_71), .B(n_153), .Y(n_464) );
INVx1_ASAP7_75t_L g109 ( .A(n_72), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_73), .Y(n_203) );
INVx1_ASAP7_75t_L g226 ( .A(n_74), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_76), .A2(n_140), .B(n_143), .C(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_77), .B(n_475), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_78), .B(n_153), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_79), .B(n_148), .Y(n_216) );
INVx2_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_81), .B(n_168), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_82), .B(n_153), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_83), .A2(n_140), .B(n_143), .C(n_146), .Y(n_142) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_84), .B(n_106), .C(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g434 ( .A(n_84), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g445 ( .A(n_84), .B(n_436), .Y(n_445) );
INVx2_ASAP7_75t_L g450 ( .A(n_84), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_86), .A2(n_100), .B1(n_153), .B2(n_154), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_87), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_88), .B(n_158), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_89), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_90), .A2(n_140), .B(n_143), .C(n_239), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_91), .Y(n_246) );
INVx1_ASAP7_75t_L g166 ( .A(n_92), .Y(n_166) );
CKINVDCx16_ASAP7_75t_R g252 ( .A(n_93), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_94), .B(n_148), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_95), .B(n_153), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_96), .B(n_161), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_97), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_98), .B(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_99), .A2(n_163), .B(n_164), .Y(n_162) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x2_ASAP7_75t_L g436 ( .A(n_106), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AO21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_115), .B(n_440), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx3_ASAP7_75t_L g736 ( .A(n_112), .Y(n_736) );
INVx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI21xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_432), .B(n_438), .Y(n_115) );
XNOR2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g446 ( .A(n_120), .Y(n_446) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_120), .A2(n_447), .B1(n_452), .B2(n_732), .Y(n_731) );
NAND2x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_348), .Y(n_120) );
NOR5xp2_ASAP7_75t_L g121 ( .A(n_122), .B(n_271), .C(n_303), .D(n_318), .E(n_335), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_187), .B(n_208), .C(n_259), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_159), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_124), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_124), .B(n_323), .Y(n_386) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_125), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_125), .B(n_205), .Y(n_272) );
AND2x2_ASAP7_75t_L g313 ( .A(n_125), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_125), .B(n_282), .Y(n_317) );
OR2x2_ASAP7_75t_L g354 ( .A(n_125), .B(n_193), .Y(n_354) );
INVx3_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g192 ( .A(n_126), .B(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g262 ( .A(n_126), .Y(n_262) );
OR2x2_ASAP7_75t_L g425 ( .A(n_126), .B(n_265), .Y(n_425) );
AO21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_133), .B(n_155), .Y(n_126) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_127), .A2(n_194), .B(n_202), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_127), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g221 ( .A(n_127), .Y(n_221) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_128), .Y(n_161) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_129), .B(n_130), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_135), .B(n_142), .Y(n_133) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_135), .A2(n_173), .B1(n_195), .B2(n_201), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_135), .A2(n_226), .B(n_227), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
AND2x4_ASAP7_75t_L g163 ( .A(n_136), .B(n_140), .Y(n_163) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g528 ( .A(n_137), .Y(n_528) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g144 ( .A(n_138), .Y(n_144) );
INVx1_ASAP7_75t_L g154 ( .A(n_138), .Y(n_154) );
INVx1_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx3_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_139), .Y(n_151) );
INVx1_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_139), .Y(n_197) );
INVx4_ASAP7_75t_SL g173 ( .A(n_140), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_140), .A2(n_462), .B(n_465), .Y(n_461) );
BUFx3_ASAP7_75t_L g477 ( .A(n_140), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_140), .A2(n_482), .B(n_486), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_140), .A2(n_522), .B(n_526), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_140), .A2(n_535), .B(n_538), .Y(n_534) );
INVx5_ASAP7_75t_L g165 ( .A(n_143), .Y(n_165) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
BUFx3_ASAP7_75t_L g220 ( .A(n_144), .Y(n_220) );
INVx1_ASAP7_75t_L g475 ( .A(n_144), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_150), .C(n_152), .Y(n_146) );
O2A1O1Ixp5_ASAP7_75t_SL g462 ( .A1(n_148), .A2(n_171), .B(n_463), .C(n_464), .Y(n_462) );
INVx2_ASAP7_75t_L g499 ( .A(n_148), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_148), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_148), .A2(n_545), .B(n_546), .Y(n_544) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_149), .B(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_149), .B(n_185), .Y(n_184) );
OAI22xp5_ASAP7_75t_SL g473 ( .A1(n_149), .A2(n_151), .B1(n_474), .B2(n_476), .Y(n_473) );
INVx2_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
INVx4_ASAP7_75t_L g242 ( .A(n_151), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_151), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_151), .A2(n_499), .B1(n_515), .B2(n_516), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_152), .A2(n_523), .B(n_524), .C(n_525), .Y(n_522) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_157), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_157), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g236 ( .A(n_158), .Y(n_236) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_158), .A2(n_249), .B(n_258), .Y(n_248) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_158), .A2(n_461), .B(n_468), .Y(n_460) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_158), .A2(n_481), .B(n_489), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g327 ( .A1(n_159), .A2(n_328), .B1(n_329), .B2(n_332), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_159), .B(n_262), .Y(n_411) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_177), .Y(n_159) );
AND2x2_ASAP7_75t_L g207 ( .A(n_160), .B(n_193), .Y(n_207) );
AND2x2_ASAP7_75t_L g264 ( .A(n_160), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g269 ( .A(n_160), .Y(n_269) );
INVx3_ASAP7_75t_L g282 ( .A(n_160), .Y(n_282) );
OR2x2_ASAP7_75t_L g302 ( .A(n_160), .B(n_265), .Y(n_302) );
AND2x2_ASAP7_75t_L g321 ( .A(n_160), .B(n_178), .Y(n_321) );
BUFx2_ASAP7_75t_L g353 ( .A(n_160), .Y(n_353) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_174), .Y(n_160) );
INVx4_ASAP7_75t_L g176 ( .A(n_161), .Y(n_176) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_161), .A2(n_534), .B(n_541), .Y(n_533) );
BUFx2_ASAP7_75t_L g250 ( .A(n_163), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_167), .C(n_173), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_165), .A2(n_173), .B(n_181), .C(n_182), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g251 ( .A1(n_165), .A2(n_173), .B(n_252), .C(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g485 ( .A(n_168), .Y(n_485) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_172), .Y(n_243) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_175), .A2(n_179), .B(n_186), .Y(n_178) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_176), .B(n_223), .Y(n_222) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_176), .B(n_477), .C(n_514), .Y(n_513) );
AO21x1_ASAP7_75t_L g603 ( .A1(n_176), .A2(n_514), .B(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_L g268 ( .A(n_177), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
BUFx2_ASAP7_75t_L g191 ( .A(n_178), .Y(n_191) );
INVx2_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
OR2x2_ASAP7_75t_L g284 ( .A(n_178), .B(n_265), .Y(n_284) );
AND2x2_ASAP7_75t_L g314 ( .A(n_178), .B(n_193), .Y(n_314) );
AND2x2_ASAP7_75t_L g331 ( .A(n_178), .B(n_262), .Y(n_331) );
AND2x2_ASAP7_75t_L g371 ( .A(n_178), .B(n_282), .Y(n_371) );
AND2x2_ASAP7_75t_SL g407 ( .A(n_178), .B(n_207), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_183), .A2(n_487), .B(n_488), .Y(n_486) );
O2A1O1Ixp5_ASAP7_75t_L g547 ( .A1(n_183), .A2(n_527), .B(n_548), .C(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp33_ASAP7_75t_SL g188 ( .A(n_189), .B(n_204), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_192), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_190), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
OAI21xp33_ASAP7_75t_L g345 ( .A1(n_191), .A2(n_207), .B(n_346), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_191), .B(n_193), .Y(n_401) );
AND2x2_ASAP7_75t_L g337 ( .A(n_192), .B(n_338), .Y(n_337) );
INVx3_ASAP7_75t_L g265 ( .A(n_193), .Y(n_265) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_193), .Y(n_363) );
OAI22xp5_ASAP7_75t_SL g196 ( .A1(n_197), .A2(n_198), .B1(n_199), .B2(n_200), .Y(n_196) );
INVx2_ASAP7_75t_L g199 ( .A(n_197), .Y(n_199) );
INVx4_ASAP7_75t_L g254 ( .A(n_197), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_204), .B(n_262), .Y(n_430) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_205), .A2(n_373), .B1(n_374), .B2(n_379), .Y(n_372) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
AND2x2_ASAP7_75t_L g263 ( .A(n_206), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g301 ( .A(n_206), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g338 ( .A(n_206), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_207), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g392 ( .A(n_207), .Y(n_392) );
CKINVDCx16_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_234), .Y(n_209) );
INVx4_ASAP7_75t_L g278 ( .A(n_210), .Y(n_278) );
AND2x2_ASAP7_75t_L g356 ( .A(n_210), .B(n_323), .Y(n_356) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_224), .Y(n_210) );
INVx3_ASAP7_75t_L g275 ( .A(n_211), .Y(n_275) );
AND2x2_ASAP7_75t_L g289 ( .A(n_211), .B(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g293 ( .A(n_211), .Y(n_293) );
INVx2_ASAP7_75t_L g307 ( .A(n_211), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_211), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g364 ( .A(n_211), .B(n_359), .Y(n_364) );
AND2x2_ASAP7_75t_L g429 ( .A(n_211), .B(n_399), .Y(n_429) );
OR2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
AOI21xp5_ASAP7_75t_SL g212 ( .A1(n_213), .A2(n_214), .B(n_221), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_218), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_218), .A2(n_229), .B(n_230), .Y(n_228) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g257 ( .A(n_220), .Y(n_257) );
INVx1_ASAP7_75t_L g231 ( .A(n_221), .Y(n_231) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_221), .A2(n_521), .B(n_531), .Y(n_520) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_221), .A2(n_543), .B(n_550), .Y(n_542) );
AND2x2_ASAP7_75t_L g270 ( .A(n_224), .B(n_248), .Y(n_270) );
INVx2_ASAP7_75t_L g290 ( .A(n_224), .Y(n_290) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_231), .B(n_232), .Y(n_224) );
INVx1_ASAP7_75t_L g295 ( .A(n_234), .Y(n_295) );
AND2x2_ASAP7_75t_L g341 ( .A(n_234), .B(n_289), .Y(n_341) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_247), .Y(n_234) );
INVx2_ASAP7_75t_L g280 ( .A(n_235), .Y(n_280) );
INVx1_ASAP7_75t_L g288 ( .A(n_235), .Y(n_288) );
AND2x2_ASAP7_75t_L g306 ( .A(n_235), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_235), .B(n_290), .Y(n_344) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_245), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_243), .Y(n_239) );
AND2x2_ASAP7_75t_L g323 ( .A(n_247), .B(n_280), .Y(n_323) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g276 ( .A(n_248), .Y(n_276) );
AND2x2_ASAP7_75t_L g359 ( .A(n_248), .B(n_290), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_254), .B(n_256), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_254), .A2(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g525 ( .A(n_254), .Y(n_525) );
OAI21xp5_ASAP7_75t_SL g259 ( .A1(n_260), .A2(n_266), .B(n_270), .Y(n_259) );
INVx1_ASAP7_75t_SL g304 ( .A(n_260), .Y(n_304) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_261), .B(n_268), .Y(n_361) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g310 ( .A(n_262), .B(n_265), .Y(n_310) );
AND2x2_ASAP7_75t_L g339 ( .A(n_262), .B(n_283), .Y(n_339) );
OR2x2_ASAP7_75t_L g342 ( .A(n_262), .B(n_302), .Y(n_342) );
AOI222xp33_ASAP7_75t_L g406 ( .A1(n_263), .A2(n_355), .B1(n_407), .B2(n_408), .C1(n_410), .C2(n_412), .Y(n_406) );
BUFx2_ASAP7_75t_L g320 ( .A(n_265), .Y(n_320) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g309 ( .A(n_268), .B(n_310), .Y(n_309) );
INVx3_ASAP7_75t_SL g326 ( .A(n_268), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_268), .B(n_320), .Y(n_380) );
AND2x2_ASAP7_75t_L g315 ( .A(n_270), .B(n_275), .Y(n_315) );
INVx1_ASAP7_75t_L g334 ( .A(n_270), .Y(n_334) );
OAI221xp5_ASAP7_75t_SL g271 ( .A1(n_272), .A2(n_273), .B1(n_277), .B2(n_281), .C(n_285), .Y(n_271) );
OR2x2_ASAP7_75t_L g343 ( .A(n_273), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x2_ASAP7_75t_L g328 ( .A(n_275), .B(n_298), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_275), .B(n_288), .Y(n_368) );
AND2x2_ASAP7_75t_L g373 ( .A(n_275), .B(n_323), .Y(n_373) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_275), .Y(n_383) );
NAND2x1_ASAP7_75t_SL g394 ( .A(n_275), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g279 ( .A(n_276), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g299 ( .A(n_276), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_276), .B(n_294), .Y(n_325) );
INVx1_ASAP7_75t_L g391 ( .A(n_276), .Y(n_391) );
INVx1_ASAP7_75t_L g366 ( .A(n_277), .Y(n_366) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g378 ( .A(n_278), .Y(n_378) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_278), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g395 ( .A(n_279), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_279), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g298 ( .A(n_280), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_280), .B(n_290), .Y(n_311) );
INVx1_ASAP7_75t_L g377 ( .A(n_280), .Y(n_377) );
INVx1_ASAP7_75t_L g398 ( .A(n_281), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OAI21xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_291), .B(n_300), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
AND2x2_ASAP7_75t_L g431 ( .A(n_287), .B(n_364), .Y(n_431) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g399 ( .A(n_288), .B(n_359), .Y(n_399) );
AOI32xp33_ASAP7_75t_L g312 ( .A1(n_289), .A2(n_295), .A3(n_313), .B1(n_315), .B2(n_316), .Y(n_312) );
AOI322xp5_ASAP7_75t_L g414 ( .A1(n_289), .A2(n_321), .A3(n_404), .B1(n_415), .B2(n_416), .C1(n_417), .C2(n_419), .Y(n_414) );
INVx2_ASAP7_75t_L g294 ( .A(n_290), .Y(n_294) );
INVx1_ASAP7_75t_L g404 ( .A(n_290), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B1(n_296), .B2(n_297), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_292), .B(n_298), .Y(n_347) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_293), .B(n_359), .Y(n_409) );
INVx1_ASAP7_75t_L g296 ( .A(n_294), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_294), .B(n_323), .Y(n_413) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_302), .B(n_397), .Y(n_396) );
OAI221xp5_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_305), .B1(n_308), .B2(n_311), .C(n_312), .Y(n_303) );
OR2x2_ASAP7_75t_L g324 ( .A(n_305), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g333 ( .A(n_305), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g358 ( .A(n_306), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g362 ( .A(n_316), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI221xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B1(n_324), .B2(n_326), .C(n_327), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_320), .A2(n_351), .B1(n_355), .B2(n_356), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_321), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g426 ( .A(n_321), .Y(n_426) );
INVx1_ASAP7_75t_L g420 ( .A(n_323), .Y(n_420) );
INVx1_ASAP7_75t_SL g355 ( .A(n_324), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_326), .B(n_354), .Y(n_416) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_331), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g397 ( .A(n_331), .Y(n_397) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OAI221xp5_ASAP7_75t_SL g335 ( .A1(n_336), .A2(n_340), .B1(n_342), .B2(n_343), .C(n_345), .Y(n_335) );
NOR2xp33_ASAP7_75t_SL g336 ( .A(n_337), .B(n_339), .Y(n_336) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_337), .A2(n_355), .B1(n_401), .B2(n_402), .Y(n_400) );
CKINVDCx14_ASAP7_75t_R g340 ( .A(n_341), .Y(n_340) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_342), .A2(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR3xp33_ASAP7_75t_SL g348 ( .A(n_349), .B(n_381), .C(n_405), .Y(n_348) );
NAND4xp25_ASAP7_75t_L g349 ( .A(n_350), .B(n_357), .C(n_365), .D(n_372), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g428 ( .A(n_353), .Y(n_428) );
INVx3_ASAP7_75t_SL g422 ( .A(n_354), .Y(n_422) );
OR2x2_ASAP7_75t_L g427 ( .A(n_354), .B(n_428), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_362), .B2(n_364), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_359), .B(n_377), .Y(n_418) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI21xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B(n_369), .Y(n_365) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI211xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_384), .B(n_387), .C(n_400), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
AOI222xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_392), .B1(n_393), .B2(n_396), .C1(n_398), .C2(n_399), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND4xp25_ASAP7_75t_SL g424 ( .A(n_397), .B(n_425), .C(n_426), .D(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND3xp33_ASAP7_75t_SL g405 ( .A(n_406), .B(n_414), .C(n_423), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_423) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g439 ( .A(n_434), .Y(n_439) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_435), .B(n_450), .Y(n_735) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g449 ( .A(n_436), .B(n_450), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g440 ( .A1(n_438), .A2(n_441), .B(n_736), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_446), .B1(n_447), .B2(n_451), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g732 ( .A(n_444), .Y(n_732) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_648), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_597), .C(n_639), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_506), .B(n_551), .C(n_573), .Y(n_454) );
OAI211xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_469), .B(n_490), .C(n_501), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_457), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g660 ( .A(n_457), .B(n_577), .Y(n_660) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g562 ( .A(n_458), .B(n_493), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_458), .B(n_480), .Y(n_679) );
INVx1_ASAP7_75t_L g697 ( .A(n_458), .Y(n_697) );
AND2x2_ASAP7_75t_L g706 ( .A(n_458), .B(n_594), .Y(n_706) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g589 ( .A(n_459), .B(n_480), .Y(n_589) );
AND2x2_ASAP7_75t_L g647 ( .A(n_459), .B(n_594), .Y(n_647) );
INVx1_ASAP7_75t_L g691 ( .A(n_459), .Y(n_691) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g568 ( .A(n_460), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g576 ( .A(n_460), .Y(n_576) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_460), .Y(n_616) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_478), .Y(n_470) );
AND2x2_ASAP7_75t_L g555 ( .A(n_471), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g588 ( .A(n_471), .Y(n_588) );
OR2x2_ASAP7_75t_L g714 ( .A(n_471), .B(n_715), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_471), .B(n_480), .Y(n_718) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g493 ( .A(n_472), .Y(n_493) );
INVx1_ASAP7_75t_L g504 ( .A(n_472), .Y(n_504) );
AND2x2_ASAP7_75t_L g577 ( .A(n_472), .B(n_495), .Y(n_577) );
AND2x2_ASAP7_75t_L g617 ( .A(n_472), .B(n_496), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_477), .A2(n_544), .B(n_547), .Y(n_543) );
INVxp67_ASAP7_75t_L g659 ( .A(n_478), .Y(n_659) );
AND2x4_ASAP7_75t_L g684 ( .A(n_478), .B(n_577), .Y(n_684) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_SL g575 ( .A(n_479), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g494 ( .A(n_480), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g563 ( .A(n_480), .B(n_496), .Y(n_563) );
INVx1_ASAP7_75t_L g569 ( .A(n_480), .Y(n_569) );
INVx2_ASAP7_75t_L g595 ( .A(n_480), .Y(n_595) );
AND2x2_ASAP7_75t_L g611 ( .A(n_480), .B(n_612), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_485), .Y(n_482) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_491), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g566 ( .A(n_493), .Y(n_566) );
AND2x2_ASAP7_75t_L g674 ( .A(n_493), .B(n_495), .Y(n_674) );
AND2x2_ASAP7_75t_L g591 ( .A(n_494), .B(n_576), .Y(n_591) );
AND2x2_ASAP7_75t_L g690 ( .A(n_494), .B(n_691), .Y(n_690) );
NOR2xp67_ASAP7_75t_L g612 ( .A(n_495), .B(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g715 ( .A(n_495), .B(n_576), .Y(n_715) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx2_ASAP7_75t_L g505 ( .A(n_496), .Y(n_505) );
AND2x2_ASAP7_75t_L g594 ( .A(n_496), .B(n_595), .Y(n_594) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_499), .A2(n_527), .B(n_529), .C(n_530), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_499), .A2(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
AND2x2_ASAP7_75t_L g640 ( .A(n_503), .B(n_575), .Y(n_640) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_504), .B(n_576), .Y(n_625) );
INVx2_ASAP7_75t_L g624 ( .A(n_505), .Y(n_624) );
OAI222xp33_ASAP7_75t_L g628 ( .A1(n_505), .A2(n_568), .B1(n_629), .B2(n_631), .C1(n_632), .C2(n_635), .Y(n_628) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_517), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g553 ( .A(n_510), .Y(n_553) );
OR2x2_ASAP7_75t_L g664 ( .A(n_510), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g586 ( .A(n_511), .Y(n_586) );
NOR2x1_ASAP7_75t_L g637 ( .A(n_511), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g643 ( .A(n_511), .B(n_557), .Y(n_643) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g604 ( .A(n_512), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_517), .A2(n_607), .B1(n_646), .B2(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_532), .Y(n_517) );
INVx3_ASAP7_75t_L g579 ( .A(n_518), .Y(n_579) );
OR2x2_ASAP7_75t_L g712 ( .A(n_518), .B(n_588), .Y(n_712) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g585 ( .A(n_519), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g601 ( .A(n_519), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g609 ( .A(n_519), .B(n_557), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_519), .B(n_533), .Y(n_665) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g556 ( .A(n_520), .B(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g560 ( .A(n_520), .B(n_533), .Y(n_560) );
AND2x2_ASAP7_75t_L g636 ( .A(n_520), .B(n_583), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_520), .B(n_542), .Y(n_676) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_532), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g592 ( .A(n_532), .B(n_553), .Y(n_592) );
AND2x2_ASAP7_75t_L g596 ( .A(n_532), .B(n_586), .Y(n_596) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_542), .Y(n_532) );
INVx3_ASAP7_75t_L g557 ( .A(n_533), .Y(n_557) );
AND2x2_ASAP7_75t_L g582 ( .A(n_533), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g717 ( .A(n_533), .B(n_700), .Y(n_717) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_542), .Y(n_571) );
INVx2_ASAP7_75t_L g583 ( .A(n_542), .Y(n_583) );
AND2x2_ASAP7_75t_L g627 ( .A(n_542), .B(n_603), .Y(n_627) );
INVx1_ASAP7_75t_L g670 ( .A(n_542), .Y(n_670) );
OR2x2_ASAP7_75t_L g701 ( .A(n_542), .B(n_603), .Y(n_701) );
AND2x2_ASAP7_75t_L g721 ( .A(n_542), .B(n_557), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_554), .B(n_558), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g559 ( .A(n_553), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_553), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g678 ( .A(n_555), .Y(n_678) );
INVx2_ASAP7_75t_SL g572 ( .A(n_556), .Y(n_572) );
AND2x2_ASAP7_75t_L g692 ( .A(n_556), .B(n_586), .Y(n_692) );
INVx2_ASAP7_75t_L g638 ( .A(n_557), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_557), .B(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_561), .B1(n_564), .B2(n_570), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_560), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g726 ( .A(n_560), .Y(n_726) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g651 ( .A(n_562), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_562), .B(n_594), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_563), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g667 ( .A(n_563), .B(n_616), .Y(n_667) );
INVx2_ASAP7_75t_L g723 ( .A(n_563), .Y(n_723) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AND2x2_ASAP7_75t_L g593 ( .A(n_566), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_566), .B(n_611), .Y(n_644) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_568), .B(n_588), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g705 ( .A(n_571), .Y(n_705) );
O2A1O1Ixp33_ASAP7_75t_SL g655 ( .A1(n_572), .A2(n_656), .B(n_658), .C(n_661), .Y(n_655) );
OR2x2_ASAP7_75t_L g682 ( .A(n_572), .B(n_586), .Y(n_682) );
OAI221xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_578), .B1(n_580), .B2(n_587), .C(n_590), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_575), .B(n_624), .Y(n_631) );
AND2x2_ASAP7_75t_L g673 ( .A(n_575), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g709 ( .A(n_575), .Y(n_709) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_576), .Y(n_600) );
INVx1_ASAP7_75t_L g613 ( .A(n_576), .Y(n_613) );
NOR2xp67_ASAP7_75t_L g633 ( .A(n_579), .B(n_634), .Y(n_633) );
INVxp67_ASAP7_75t_L g687 ( .A(n_579), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_579), .B(n_627), .Y(n_703) );
INVx2_ASAP7_75t_L g689 ( .A(n_580), .Y(n_689) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g630 ( .A(n_582), .B(n_601), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_582), .A2(n_598), .B(n_640), .C(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g608 ( .A(n_583), .B(n_603), .Y(n_608) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_587), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
OR2x2_ASAP7_75t_L g656 ( .A(n_588), .B(n_657), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_592), .B1(n_593), .B2(n_596), .Y(n_590) );
INVx1_ASAP7_75t_L g710 ( .A(n_592), .Y(n_710) );
INVx1_ASAP7_75t_L g657 ( .A(n_594), .Y(n_657) );
INVx1_ASAP7_75t_L g708 ( .A(n_596), .Y(n_708) );
AOI211xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_601), .B(n_605), .C(n_628), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g620 ( .A(n_600), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g671 ( .A(n_601), .Y(n_671) );
AND2x2_ASAP7_75t_L g720 ( .A(n_601), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_610), .B(n_618), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx2_ASAP7_75t_L g634 ( .A(n_608), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_608), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g626 ( .A(n_609), .B(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g702 ( .A(n_609), .Y(n_702) );
OAI32xp33_ASAP7_75t_L g713 ( .A1(n_609), .A2(n_661), .A3(n_668), .B1(n_709), .B2(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_SL g610 ( .A(n_611), .B(n_614), .Y(n_610) );
INVx1_ASAP7_75t_SL g681 ( .A(n_611), .Y(n_681) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g621 ( .A(n_617), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B(n_626), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_620), .A2(n_668), .B1(n_694), .B2(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_624), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g661 ( .A(n_627), .Y(n_661) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2x1p5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g654 ( .A(n_638), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_644), .B(n_645), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_647), .A2(n_689), .B1(n_690), .B2(n_692), .C(n_693), .Y(n_688) );
NAND5xp2_ASAP7_75t_L g648 ( .A(n_649), .B(n_672), .C(n_688), .D(n_698), .E(n_716), .Y(n_648) );
AOI211xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_652), .B(n_655), .C(n_662), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g719 ( .A(n_656), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_666), .B2(n_668), .Y(n_662) );
INVx1_ASAP7_75t_SL g695 ( .A(n_665), .Y(n_695) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
OAI322xp33_ASAP7_75t_L g677 ( .A1(n_668), .A2(n_678), .A3(n_679), .B1(n_680), .B2(n_681), .C1(n_682), .C2(n_683), .Y(n_677) );
OR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g680 ( .A(n_670), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_670), .B(n_695), .Y(n_694) );
AOI211xp5_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_675), .B(n_677), .C(n_685), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g707 ( .A1(n_681), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_707) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g724 ( .A(n_691), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_706), .B1(n_707), .B2(n_711), .C(n_713), .Y(n_698) );
OAI211xp5_ASAP7_75t_SL g699 ( .A1(n_700), .A2(n_702), .B(n_703), .C(n_704), .Y(n_699) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g725 ( .A(n_701), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_719), .B2(n_720), .C(n_722), .Y(n_716) );
AOI21xp33_ASAP7_75t_SL g722 ( .A1(n_723), .A2(n_724), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx3_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
endmodule