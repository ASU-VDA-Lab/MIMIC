module fake_jpeg_15870_n_43 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_43);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_43;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_24),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.C(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_34),
.B1(n_5),
.B2(n_6),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_8),
.B(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_12),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_37),
.B1(n_33),
.B2(n_17),
.Y(n_42)
);

AOI321xp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_38),
.A3(n_35),
.B1(n_16),
.B2(n_14),
.C(n_36),
.Y(n_43)
);


endmodule