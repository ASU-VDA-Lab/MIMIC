module fake_jpeg_14155_n_461 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_461);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_461;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_7),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_76),
.Y(n_101)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_63),
.B(n_68),
.Y(n_112)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_48),
.Y(n_98)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_16),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_19),
.B(n_13),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_20),
.A2(n_10),
.B1(n_12),
.B2(n_2),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_18),
.B1(n_38),
.B2(n_41),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_23),
.B(n_24),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_78),
.B(n_81),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_33),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_23),
.B(n_24),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_34),
.B(n_12),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_82),
.B(n_88),
.Y(n_148)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_91),
.Y(n_111)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_34),
.B(n_10),
.Y(n_88)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_37),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_39),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_38),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_45),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_42),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_48),
.B1(n_55),
.B2(n_36),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_96),
.A2(n_83),
.B1(n_69),
.B2(n_59),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_104),
.B(n_116),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_20),
.B1(n_42),
.B2(n_44),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_113),
.A2(n_123),
.B1(n_139),
.B2(n_97),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_41),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_54),
.B(n_32),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_74),
.A2(n_42),
.B1(n_44),
.B2(n_32),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_53),
.B1(n_72),
.B2(n_50),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_56),
.B(n_30),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_143),
.C(n_87),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_49),
.A2(n_20),
.B1(n_36),
.B2(n_18),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_30),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_29),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_147),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_64),
.A2(n_36),
.B1(n_29),
.B2(n_28),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_51),
.A2(n_0),
.B(n_1),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_79),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_58),
.B(n_1),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_164),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_150),
.A2(n_198),
.B1(n_143),
.B2(n_125),
.Y(n_201)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_103),
.Y(n_151)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_151),
.Y(n_235)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_152),
.Y(n_243)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_153),
.Y(n_232)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_156),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_191),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_98),
.A2(n_80),
.B1(n_67),
.B2(n_61),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_168),
.A2(n_175),
.B(n_182),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_104),
.A2(n_84),
.B1(n_75),
.B2(n_57),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_172),
.Y(n_236)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_178),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_124),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_179),
.Y(n_223)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_110),
.B(n_89),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_92),
.Y(n_177)
);

NAND2x1_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_192),
.Y(n_213)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_180),
.B(n_187),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_114),
.A2(n_52),
.B1(n_58),
.B2(n_60),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_184),
.B(n_188),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_110),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_190),
.B(n_199),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_123),
.A2(n_73),
.B1(n_86),
.B2(n_62),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_101),
.B(n_70),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_193),
.Y(n_240)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_148),
.A2(n_85),
.B(n_60),
.C(n_31),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_195),
.A2(n_192),
.B(n_160),
.C(n_164),
.Y(n_231)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_121),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_138),
.B(n_71),
.C(n_93),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_134),
.C(n_117),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_126),
.A2(n_66),
.B1(n_71),
.B2(n_31),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_107),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_167),
.B1(n_177),
.B2(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_200),
.A2(n_228),
.B1(n_234),
.B2(n_182),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_201),
.A2(n_184),
.B1(n_173),
.B2(n_159),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_163),
.B(n_112),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_203),
.B(n_220),
.C(n_226),
.Y(n_263)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_168),
.A2(n_144),
.B1(n_128),
.B2(n_106),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_168),
.B(n_180),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_215),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_118),
.B(n_117),
.Y(n_215)
);

AND2x4_ASAP7_75t_SL g217 ( 
.A(n_163),
.B(n_146),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_231),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_185),
.B(n_140),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_121),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_187),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_160),
.A2(n_114),
.B1(n_99),
.B2(n_108),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_108),
.B1(n_100),
.B2(n_109),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_197),
.A2(n_134),
.B1(n_145),
.B2(n_109),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_25),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_161),
.B(n_1),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_244),
.B(n_2),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_245),
.B(n_277),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_204),
.A2(n_99),
.B1(n_172),
.B2(n_152),
.Y(n_246)
);

AO21x2_ASAP7_75t_L g293 ( 
.A1(n_246),
.A2(n_209),
.B(n_227),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_247),
.B(n_252),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_262),
.Y(n_288)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_251),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_186),
.B1(n_100),
.B2(n_158),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_224),
.A2(n_189),
.B1(n_102),
.B2(n_136),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_253),
.A2(n_258),
.B1(n_276),
.B2(n_221),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_202),
.B(n_188),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_254),
.B(n_255),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_181),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_178),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_256),
.B(n_261),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_224),
.A2(n_136),
.B1(n_193),
.B2(n_154),
.Y(n_258)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

NOR2x1_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_156),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_203),
.Y(n_262)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_209),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_265),
.Y(n_289)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_176),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_242),
.C(n_213),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_221),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_270),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_223),
.B(n_176),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_194),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_271),
.B(n_273),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_220),
.B(n_2),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_274),
.B(n_278),
.C(n_282),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_212),
.A2(n_31),
.B1(n_25),
.B2(n_93),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_242),
.A2(n_31),
.B1(n_25),
.B2(n_4),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_2),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_217),
.B(n_3),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_217),
.B(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_232),
.Y(n_281)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_3),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_243),
.Y(n_283)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_284),
.A2(n_221),
.B(n_230),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_287),
.B(n_301),
.C(n_307),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_293),
.A2(n_305),
.B1(n_252),
.B2(n_269),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_249),
.A2(n_215),
.B(n_216),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_295),
.Y(n_348)
);

AO22x1_ASAP7_75t_SL g296 ( 
.A1(n_250),
.A2(n_216),
.B1(n_213),
.B2(n_207),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_300),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_204),
.B(n_238),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_320),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_222),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_213),
.C(n_219),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_219),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_310),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_211),
.C(n_222),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_251),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_264),
.B(n_211),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_281),
.Y(n_313)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_234),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_268),
.Y(n_325)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_265),
.Y(n_317)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_208),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_268),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_331),
.C(n_336),
.Y(n_356)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_294),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_324),
.B(n_326),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_344),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_311),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_306),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_327),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_248),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_328),
.B(n_342),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_329),
.A2(n_334),
.B1(n_346),
.B2(n_296),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_249),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_309),
.A2(n_253),
.B1(n_272),
.B2(n_258),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_332),
.A2(n_345),
.B1(n_349),
.B2(n_293),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_314),
.A2(n_250),
.B1(n_272),
.B2(n_284),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_280),
.Y(n_336)
);

NAND4xp25_ASAP7_75t_SL g337 ( 
.A(n_285),
.B(n_261),
.C(n_210),
.D(n_209),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_285),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_210),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_340),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_319),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_316),
.B(n_247),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_297),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_279),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_245),
.B1(n_260),
.B2(n_276),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_314),
.A2(n_305),
.B1(n_299),
.B2(n_286),
.Y(n_346)
);

XOR2x2_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_277),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_290),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_293),
.A2(n_259),
.B1(n_240),
.B2(n_275),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_335),
.B(n_313),
.Y(n_352)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_338),
.A2(n_286),
.B1(n_304),
.B2(n_257),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_353),
.A2(n_362),
.B1(n_368),
.B2(n_361),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_357),
.A2(n_365),
.B1(n_334),
.B2(n_347),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_330),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_358),
.B(n_367),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_359),
.B(n_337),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_348),
.A2(n_320),
.B(n_309),
.Y(n_361)
);

OAI31xp33_ASAP7_75t_L g379 ( 
.A1(n_361),
.A2(n_372),
.A3(n_373),
.B(n_333),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_303),
.Y(n_363)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_364),
.B(n_371),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_339),
.A2(n_293),
.B1(n_296),
.B2(n_289),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_333),
.B(n_298),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_369),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_370),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_346),
.B(n_298),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_348),
.A2(n_293),
.B(n_205),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_333),
.A2(n_312),
.B(n_290),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_340),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_370),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g377 ( 
.A(n_354),
.B(n_325),
.CI(n_344),
.CON(n_377),
.SN(n_377)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_364),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_379),
.A2(n_351),
.B(n_257),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_381),
.A2(n_390),
.B1(n_394),
.B2(n_395),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_350),
.C(n_321),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_386),
.C(n_397),
.Y(n_398)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_384),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_363),
.Y(n_385)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_385),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_350),
.C(n_331),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_362),
.A2(n_332),
.B1(n_345),
.B2(n_304),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_387),
.A2(n_376),
.B1(n_351),
.B2(n_374),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_336),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_391),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_371),
.A2(n_291),
.B1(n_240),
.B2(n_218),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_365),
.A2(n_283),
.B1(n_230),
.B2(n_236),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_369),
.A2(n_283),
.B1(n_243),
.B2(n_205),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_396),
.A2(n_376),
.B1(n_372),
.B2(n_355),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_354),
.B(n_214),
.C(n_235),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_369),
.C(n_373),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_404),
.Y(n_426)
);

NOR3xp33_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_388),
.C(n_382),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_375),
.C(n_366),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_385),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_380),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_406),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_370),
.C(n_360),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_407),
.B(n_411),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_370),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_408),
.B(n_414),
.Y(n_417)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_409),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_410),
.A2(n_393),
.B(n_394),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_214),
.C(n_235),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_384),
.A2(n_257),
.B(n_292),
.Y(n_413)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_413),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_232),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_422),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_420),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_381),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_387),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_421),
.B(n_406),
.C(n_403),
.Y(n_436)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_412),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_378),
.C(n_382),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_427),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_425),
.B(n_398),
.C(n_407),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_430),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_426),
.B(n_400),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_431),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_416),
.B(n_411),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_433),
.A2(n_434),
.B(n_438),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_424),
.A2(n_379),
.B(n_408),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_402),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_436),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_421),
.C(n_424),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_417),
.B(n_409),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_439),
.A2(n_395),
.B(n_390),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_417),
.C(n_414),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_441),
.A2(n_444),
.B(n_6),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_442),
.Y(n_452)
);

AOI322xp5_ASAP7_75t_L g443 ( 
.A1(n_429),
.A2(n_292),
.A3(n_377),
.B1(n_210),
.B2(n_232),
.C1(n_4),
.C2(n_8),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_443),
.B(n_446),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_432),
.Y(n_444)
);

AOI322xp5_ASAP7_75t_L g446 ( 
.A1(n_437),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_377),
.C2(n_428),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_448),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_449),
.B(n_451),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_440),
.A2(n_437),
.B(n_6),
.Y(n_450)
);

AOI21x1_ASAP7_75t_L g454 ( 
.A1(n_450),
.A2(n_453),
.B(n_452),
.Y(n_454)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_454),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_449),
.A2(n_444),
.B1(n_445),
.B2(n_447),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_456),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_457),
.B(n_455),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_459),
.B(n_458),
.C(n_441),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_460),
.B(n_8),
.Y(n_461)
);


endmodule