module fake_jpeg_32196_n_306 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_245;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_182;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_300;
wire n_211;
wire n_294;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_48),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_0),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_24),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_50),
.B(n_25),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_26),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_54),
.A2(n_78),
.B(n_95),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_17),
.B1(n_21),
.B2(n_39),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_55),
.A2(n_79),
.B1(n_84),
.B2(n_90),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_32),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_57),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_62),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_75),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_39),
.B1(n_38),
.B2(n_33),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_70),
.B1(n_76),
.B2(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_34),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_67),
.Y(n_123)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_39),
.B1(n_38),
.B2(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_28),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_38),
.B1(n_33),
.B2(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_42),
.B(n_37),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_50),
.A2(n_17),
.B1(n_21),
.B2(n_29),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_51),
.B1(n_43),
.B2(n_27),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_37),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_20),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_20),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_43),
.A2(n_36),
.B1(n_22),
.B2(n_27),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_23),
.B1(n_36),
.B2(n_22),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_94),
.Y(n_106)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_40),
.A2(n_21),
.B1(n_29),
.B2(n_19),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_23),
.B1(n_19),
.B2(n_18),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_103),
.B1(n_25),
.B2(n_5),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_28),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_45),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_100),
.Y(n_127)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_21),
.B1(n_18),
.B2(n_35),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_99),
.B1(n_25),
.B2(n_2),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_50),
.A2(n_35),
.B1(n_11),
.B2(n_3),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_47),
.A2(n_25),
.B1(n_9),
.B2(n_3),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_47),
.B(n_0),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_11),
.B(n_5),
.Y(n_124)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_84),
.B1(n_8),
.B2(n_9),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_124),
.B(n_103),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_56),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_104),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_65),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_58),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_96),
.B(n_71),
.C(n_75),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_118),
.B(n_116),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_141),
.B(n_143),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_106),
.B1(n_110),
.B2(n_131),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_147),
.A2(n_159),
.B1(n_165),
.B2(n_151),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_149),
.B(n_6),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_106),
.B(n_71),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_154),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_94),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_153),
.A2(n_86),
.B1(n_13),
.B2(n_14),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_106),
.B(n_60),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_155),
.B(n_157),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_100),
.A3(n_60),
.B1(n_97),
.B2(n_77),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_156),
.B(n_158),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_95),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_70),
.B1(n_76),
.B2(n_102),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_59),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_161),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_109),
.A2(n_73),
.B1(n_88),
.B2(n_89),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_74),
.B(n_59),
.Y(n_196)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_113),
.B(n_101),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_77),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_112),
.B(n_118),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_72),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_114),
.B1(n_116),
.B2(n_107),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_170),
.A2(n_186),
.B1(n_192),
.B2(n_197),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_178),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_108),
.B(n_135),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_175),
.A2(n_12),
.B(n_14),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_148),
.A2(n_117),
.B1(n_132),
.B2(n_105),
.Y(n_178)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_132),
.B(n_74),
.C(n_69),
.D(n_107),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_194),
.B(n_146),
.Y(n_206)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_189),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_72),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_102),
.B1(n_91),
.B2(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

HAxp5_ASAP7_75t_SL g194 ( 
.A(n_154),
.B(n_105),
.CON(n_194),
.SN(n_194)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_142),
.B(n_61),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_147),
.A2(n_115),
.B1(n_86),
.B2(n_61),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_201),
.Y(n_211)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_149),
.B(n_12),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_160),
.B1(n_138),
.B2(n_145),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_148),
.B1(n_153),
.B2(n_157),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_209),
.B1(n_226),
.B2(n_202),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_151),
.C(n_150),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_171),
.C(n_188),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_178),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_208),
.B(n_213),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_141),
.B1(n_156),
.B2(n_166),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_201),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_210),
.B(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_167),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_197),
.B1(n_192),
.B2(n_176),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_195),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_223),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_218),
.A2(n_196),
.B(n_176),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_74),
.B(n_168),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_183),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_177),
.B(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_222),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_175),
.B(n_190),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_191),
.B(n_160),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_152),
.B1(n_160),
.B2(n_163),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_243),
.B1(n_224),
.B2(n_226),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_241),
.B(n_208),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_213),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_231),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_188),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_235),
.C(n_242),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_187),
.C(n_189),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_215),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_239),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_187),
.C(n_185),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_181),
.Y(n_244)
);

XOR2x2_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_207),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_204),
.A2(n_172),
.B1(n_193),
.B2(n_174),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_246),
.B1(n_203),
.B2(n_214),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_172),
.B1(n_174),
.B2(n_200),
.Y(n_246)
);

OA21x2_ASAP7_75t_SL g247 ( 
.A1(n_227),
.A2(n_216),
.B(n_211),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_248),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g248 ( 
.A(n_240),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_207),
.B(n_223),
.Y(n_249)
);

OAI31xp33_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_254),
.A3(n_221),
.B(n_217),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_234),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_232),
.B(n_203),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_207),
.B(n_218),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_261),
.B(n_229),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_258),
.B1(n_233),
.B2(n_244),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_242),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_236),
.B(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_219),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_257),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_254),
.B1(n_249),
.B2(n_255),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_253),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_270),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_230),
.C(n_235),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_252),
.C(n_259),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_256),
.Y(n_279)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_251),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_231),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_250),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_278),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_282),
.C(n_266),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_280),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_182),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_262),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_283),
.A2(n_268),
.B1(n_272),
.B2(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_289),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_264),
.B1(n_267),
.B2(n_179),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_280),
.A2(n_274),
.B(n_181),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_288),
.B(n_277),
.Y(n_293)
);

AOI221xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_182),
.B1(n_180),
.B2(n_163),
.C(n_16),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_275),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_296),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_282),
.B1(n_275),
.B2(n_152),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_285),
.C(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_292),
.C(n_291),
.Y(n_300)
);

A2O1A1Ixp33_ASAP7_75t_SL g303 ( 
.A1(n_301),
.A2(n_12),
.B(n_14),
.C(n_15),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_303),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_302),
.C(n_298),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_294),
.Y(n_306)
);


endmodule