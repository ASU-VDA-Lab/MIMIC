module fake_netlist_5_206_n_687 (n_137, n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_687);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_687;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_280;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_671;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_668;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_546;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_264;
wire n_669;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_550;
wire n_522;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_638;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_571;
wire n_461;
wire n_333;
wire n_477;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_666;
wire n_538;
wire n_262;
wire n_238;
wire n_639;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

BUFx3_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_52),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_12),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_88),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_48),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_63),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_64),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_28),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_45),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_39),
.Y(n_156)
);

NOR2xp67_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_128),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_21),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_78),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_121),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_54),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_117),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_123),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_83),
.B(n_57),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_1),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_15),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_79),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_42),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_10),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_61),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_40),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_34),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_58),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_33),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_26),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_18),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_112),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_98),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_85),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_7),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_56),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_80),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_15),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_95),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_59),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_192),
.A2(n_0),
.B(n_1),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_141),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_171),
.Y(n_208)
);

AND2x4_ASAP7_75t_L g209 ( 
.A(n_140),
.B(n_19),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_143),
.Y(n_210)
);

OA21x2_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_2),
.B(n_4),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_4),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_5),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_141),
.Y(n_214)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_181),
.A2(n_5),
.B(n_6),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_6),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_218)
);

AOI22x1_ASAP7_75t_SL g219 ( 
.A1(n_176),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_146),
.Y(n_223)
);

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_142),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_149),
.Y(n_225)
);

NOR2x1_ASAP7_75t_L g226 ( 
.A(n_157),
.B(n_20),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_151),
.B(n_11),
.Y(n_227)
);

OAI21x1_ASAP7_75t_L g228 ( 
.A1(n_152),
.A2(n_11),
.B(n_12),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_153),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_156),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_142),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_174),
.B(n_13),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_159),
.B(n_14),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_144),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_174),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_168),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_179),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_179),
.B1(n_182),
.B2(n_164),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_170),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_203),
.Y(n_243)
);

INVxp33_ASAP7_75t_SL g244 ( 
.A(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

NAND2xp33_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_178),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_175),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_220),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_205),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_177),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_196),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_208),
.B(n_145),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_231),
.Y(n_261)
);

OR2x6_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_169),
.Y(n_262)
);

NAND2xp33_ASAP7_75t_SL g263 ( 
.A(n_216),
.B(n_184),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_189),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_208),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_198),
.A2(n_193),
.B1(n_190),
.B2(n_187),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_202),
.B(n_183),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_201),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_234),
.B(n_147),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_202),
.B(n_180),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_148),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_223),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_172),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_150),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_241),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_221),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_198),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_158),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_206),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_206),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_226),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g292 ( 
.A1(n_244),
.A2(n_232),
.B1(n_218),
.B2(n_197),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_206),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

NOR3xp33_ASAP7_75t_L g297 ( 
.A(n_239),
.B(n_207),
.C(n_228),
.Y(n_297)
);

AO221x1_ASAP7_75t_L g298 ( 
.A1(n_263),
.A2(n_228),
.B1(n_230),
.B2(n_229),
.C(n_236),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_L g299 ( 
.A1(n_242),
.A2(n_215),
.B(n_222),
.C(n_207),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_240),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_245),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_257),
.B(n_160),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_240),
.B(n_223),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_SL g304 ( 
.A(n_263),
.B(n_161),
.C(n_162),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_246),
.B(n_223),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_244),
.A2(n_211),
.B1(n_197),
.B2(n_215),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_236),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_237),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_R g311 ( 
.A(n_251),
.B(n_163),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_277),
.B(n_165),
.Y(n_313)
);

A2O1A1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_251),
.A2(n_222),
.B(n_195),
.C(n_229),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_273),
.A2(n_211),
.B(n_197),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_259),
.B(n_195),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_262),
.A2(n_211),
.B1(n_230),
.B2(n_236),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_258),
.B(n_230),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_250),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_266),
.A2(n_236),
.B(n_230),
.C(n_219),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_261),
.B(n_230),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_266),
.B(n_236),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_271),
.B(n_200),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_243),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_258),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_268),
.B(n_22),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_255),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_268),
.B(n_276),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_23),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_270),
.B(n_24),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_252),
.A2(n_224),
.B1(n_219),
.B2(n_16),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_292),
.B(n_262),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_282),
.B(n_270),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_300),
.A2(n_294),
.B(n_315),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_285),
.B(n_255),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_287),
.A2(n_256),
.B(n_262),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_285),
.B(n_256),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_283),
.B(n_17),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_301),
.Y(n_340)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_311),
.B(n_17),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_289),
.A2(n_25),
.B(n_27),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_329),
.A2(n_29),
.B(n_30),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_308),
.A2(n_31),
.B(n_32),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_326),
.Y(n_347)
);

CKINVDCx10_ASAP7_75t_R g348 ( 
.A(n_332),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g349 ( 
.A1(n_297),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_349)
);

AOI21x1_ASAP7_75t_L g350 ( 
.A1(n_303),
.A2(n_38),
.B(n_41),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_311),
.B(n_43),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_308),
.A2(n_44),
.B(n_46),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_310),
.B(n_47),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_309),
.B(n_49),
.Y(n_354)
);

INVxp33_ASAP7_75t_SL g355 ( 
.A(n_281),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_317),
.A2(n_50),
.B(n_51),
.Y(n_356)
);

AO21x1_ASAP7_75t_L g357 ( 
.A1(n_286),
.A2(n_53),
.B(n_55),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_290),
.B(n_293),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_60),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_284),
.B(n_62),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_65),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_327),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_304),
.A2(n_302),
.B1(n_313),
.B2(n_325),
.Y(n_365)
);

O2A1O1Ixp5_ASAP7_75t_L g366 ( 
.A1(n_322),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_366)
);

NOR3xp33_ASAP7_75t_L g367 ( 
.A(n_320),
.B(n_72),
.C(n_73),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_291),
.A2(n_74),
.B(n_75),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_331),
.A2(n_76),
.B(n_77),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_316),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_280),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_314),
.A2(n_323),
.B(n_328),
.C(n_296),
.Y(n_372)
);

AND3x2_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_86),
.C(n_87),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_323),
.B(n_90),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_306),
.B(n_91),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_307),
.B(n_92),
.Y(n_377)
);

AOI21x1_ASAP7_75t_L g378 ( 
.A1(n_318),
.A2(n_96),
.B(n_97),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_306),
.B(n_99),
.Y(n_379)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_312),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_312),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_319),
.B(n_101),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_319),
.B(n_321),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_298),
.B(n_102),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_315),
.A2(n_103),
.B(n_104),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_310),
.A2(n_105),
.B1(n_107),
.B2(n_109),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_335),
.A2(n_110),
.B(n_111),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_346),
.A2(n_113),
.B(n_116),
.Y(n_389)
);

NOR2x1_ASAP7_75t_SL g390 ( 
.A(n_384),
.B(n_118),
.Y(n_390)
);

AO31x2_ASAP7_75t_L g391 ( 
.A1(n_372),
.A2(n_119),
.A3(n_122),
.B(n_126),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_381),
.Y(n_392)
);

AOI21xp33_ASAP7_75t_L g393 ( 
.A1(n_333),
.A2(n_130),
.B(n_132),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_334),
.A2(n_133),
.B(n_134),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_352),
.A2(n_135),
.B1(n_139),
.B2(n_356),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

AO21x2_ASAP7_75t_L g397 ( 
.A1(n_385),
.A2(n_352),
.B(n_354),
.Y(n_397)
);

NOR2x1_ASAP7_75t_SL g398 ( 
.A(n_347),
.B(n_360),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_337),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_340),
.B(n_344),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_375),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_355),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_358),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_342),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_349),
.A2(n_363),
.B1(n_359),
.B2(n_369),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_375),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_380),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_379),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_348),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_341),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_333),
.B(n_365),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_367),
.A2(n_383),
.B(n_353),
.C(n_366),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_341),
.B(n_360),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_350),
.A2(n_378),
.B(n_374),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_347),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_351),
.A2(n_382),
.B(n_376),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_347),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_360),
.A2(n_377),
.B(n_368),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_373),
.B(n_370),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_345),
.A2(n_343),
.B(n_357),
.Y(n_421)
);

AOI221xp5_ASAP7_75t_SL g422 ( 
.A1(n_386),
.A2(n_292),
.B1(n_352),
.B2(n_346),
.C(n_299),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_355),
.B(n_239),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_336),
.B(n_338),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_335),
.A2(n_346),
.B(n_315),
.Y(n_425)
);

NAND2x1p5_ASAP7_75t_L g426 ( 
.A(n_351),
.B(n_375),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_381),
.Y(n_427)
);

O2A1O1Ixp5_ASAP7_75t_L g428 ( 
.A1(n_384),
.A2(n_356),
.B(n_315),
.C(n_346),
.Y(n_428)
);

AO32x2_ASAP7_75t_L g429 ( 
.A1(n_365),
.A2(n_364),
.A3(n_370),
.B1(n_380),
.B2(n_375),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_340),
.B(n_344),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_396),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g432 ( 
.A(n_427),
.Y(n_432)
);

O2A1O1Ixp33_ASAP7_75t_SL g433 ( 
.A1(n_395),
.A2(n_389),
.B(n_411),
.C(n_405),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_402),
.Y(n_434)
);

O2A1O1Ixp33_ASAP7_75t_SL g435 ( 
.A1(n_395),
.A2(n_389),
.B(n_405),
.C(n_425),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_388),
.Y(n_436)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_419),
.A2(n_415),
.B(n_421),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_402),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_403),
.Y(n_440)
);

CKINVDCx6p67_ASAP7_75t_R g441 ( 
.A(n_427),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_420),
.A2(n_397),
.B1(n_393),
.B2(n_387),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_427),
.Y(n_443)
);

AOI21xp33_ASAP7_75t_L g444 ( 
.A1(n_422),
.A2(n_404),
.B(n_397),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_392),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_416),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_408),
.A2(n_425),
.B(n_428),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_410),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_387),
.A2(n_417),
.B1(n_418),
.B2(n_399),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_406),
.A2(n_417),
.B1(n_401),
.B2(n_426),
.Y(n_452)
);

AO31x2_ASAP7_75t_L g453 ( 
.A1(n_413),
.A2(n_390),
.A3(n_398),
.B(n_394),
.Y(n_453)
);

CKINVDCx6p67_ASAP7_75t_R g454 ( 
.A(n_409),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_401),
.A2(n_414),
.B(n_426),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_418),
.B(n_416),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_407),
.A2(n_412),
.B(n_422),
.Y(n_457)
);

AOI21x1_ASAP7_75t_L g458 ( 
.A1(n_429),
.A2(n_391),
.B(n_409),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_429),
.A2(n_428),
.B(n_395),
.Y(n_459)
);

AO21x2_ASAP7_75t_L g460 ( 
.A1(n_429),
.A2(n_425),
.B(n_417),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_391),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_391),
.B(n_430),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_423),
.B(n_355),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_400),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_416),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_416),
.Y(n_466)
);

OA21x2_ASAP7_75t_L g467 ( 
.A1(n_425),
.A2(n_428),
.B(n_422),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_395),
.A2(n_411),
.B1(n_389),
.B2(n_333),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_396),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_438),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_431),
.B(n_469),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_470),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_464),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_463),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_462),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_443),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_462),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_434),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_436),
.Y(n_482)
);

NAND2x1p5_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_467),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_449),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_468),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_439),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_450),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_466),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_443),
.Y(n_490)
);

OAI21xp33_ASAP7_75t_SL g491 ( 
.A1(n_459),
.A2(n_451),
.B(n_442),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_466),
.Y(n_492)
);

AO21x2_ASAP7_75t_L g493 ( 
.A1(n_435),
.A2(n_448),
.B(n_433),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_466),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_439),
.B(n_460),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_469),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_466),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_467),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_431),
.A2(n_466),
.B1(n_442),
.B2(n_447),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_437),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_453),
.Y(n_502)
);

INVxp33_ASAP7_75t_L g503 ( 
.A(n_447),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_465),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_432),
.B(n_446),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_453),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_444),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_496),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_482),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_496),
.B(n_461),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_485),
.B(n_446),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_488),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_488),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_495),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_471),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_479),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_495),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_490),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_499),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_499),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_502),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_473),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_494),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_473),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_478),
.B(n_453),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_476),
.B(n_441),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_472),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_474),
.Y(n_529)
);

OR2x2_ASAP7_75t_SL g530 ( 
.A(n_489),
.B(n_433),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_485),
.B(n_476),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_507),
.B(n_451),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_507),
.B(n_465),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_478),
.B(n_465),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_506),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_480),
.B(n_452),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_474),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_475),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_480),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_475),
.B(n_454),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_491),
.B(n_435),
.C(n_500),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_484),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_505),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_489),
.B(n_498),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_484),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_483),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_526),
.B(n_498),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_516),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_516),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_517),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_513),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_519),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_503),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_513),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_543),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_509),
.B(n_511),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_514),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_509),
.B(n_493),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_518),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_526),
.Y(n_560)
);

INVxp67_ASAP7_75t_SL g561 ( 
.A(n_533),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_526),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_511),
.B(n_491),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_520),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_508),
.B(n_483),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_531),
.B(n_497),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_512),
.B(n_481),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_508),
.B(n_512),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_544),
.B(n_492),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_527),
.B(n_473),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_518),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_521),
.B(n_487),
.Y(n_572)
);

NOR2xp67_ASAP7_75t_L g573 ( 
.A(n_541),
.B(n_501),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_524),
.B(n_505),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_561),
.B(n_532),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_550),
.B(n_552),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_565),
.B(n_521),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_565),
.B(n_536),
.Y(n_578)
);

NAND2x1_ASAP7_75t_L g579 ( 
.A(n_562),
.B(n_535),
.Y(n_579)
);

INVxp33_ASAP7_75t_L g580 ( 
.A(n_570),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_548),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_555),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_548),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_549),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_549),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_568),
.B(n_536),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_568),
.B(n_522),
.Y(n_587)
);

AND2x4_ASAP7_75t_SL g588 ( 
.A(n_569),
.B(n_518),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_556),
.B(n_532),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_558),
.B(n_522),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_551),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_551),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_553),
.B(n_541),
.C(n_540),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_556),
.B(n_543),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_567),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_563),
.A2(n_525),
.B1(n_523),
.B2(n_515),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_554),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_562),
.B(n_546),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_566),
.B(n_528),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_554),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_557),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_557),
.Y(n_602)
);

NAND2x1_ASAP7_75t_SL g603 ( 
.A(n_573),
.B(n_546),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_575),
.B(n_564),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_600),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_578),
.B(n_560),
.Y(n_606)
);

AOI32xp33_ASAP7_75t_L g607 ( 
.A1(n_580),
.A2(n_540),
.A3(n_560),
.B1(n_547),
.B2(n_569),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_583),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_593),
.A2(n_573),
.B1(n_530),
.B2(n_574),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_600),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_577),
.B(n_562),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_582),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_583),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_595),
.A2(n_530),
.B1(n_515),
.B2(n_539),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_577),
.B(n_576),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_584),
.Y(n_616)
);

NAND2x1_ASAP7_75t_L g617 ( 
.A(n_598),
.B(n_564),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_584),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_592),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_592),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_581),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_598),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_613),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_578),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_605),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_604),
.B(n_615),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_604),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_621),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_606),
.B(n_586),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_609),
.A2(n_580),
.B1(n_525),
.B2(n_547),
.Y(n_630)
);

OAI221xp5_ASAP7_75t_L g631 ( 
.A1(n_609),
.A2(n_596),
.B1(n_599),
.B2(n_589),
.C(n_594),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_616),
.B(n_586),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_622),
.B(n_590),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_626),
.B(n_611),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_627),
.B(n_619),
.Y(n_635)
);

AO21x1_ASAP7_75t_L g636 ( 
.A1(n_625),
.A2(n_617),
.B(n_614),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_633),
.B(n_622),
.Y(n_637)
);

AOI31xp33_ASAP7_75t_L g638 ( 
.A1(n_630),
.A2(n_614),
.A3(n_569),
.B(n_559),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_632),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_624),
.B(n_571),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_640),
.B(n_631),
.Y(n_641)
);

OAI221xp5_ASAP7_75t_SL g642 ( 
.A1(n_635),
.A2(n_607),
.B1(n_628),
.B2(n_629),
.C(n_623),
.Y(n_642)
);

AOI221xp5_ASAP7_75t_L g643 ( 
.A1(n_636),
.A2(n_623),
.B1(n_610),
.B2(n_620),
.C(n_608),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_638),
.A2(n_639),
.B(n_634),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_638),
.A2(n_579),
.B(n_585),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_641),
.B(n_639),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_644),
.B(n_637),
.Y(n_647)
);

OAI211xp5_ASAP7_75t_L g648 ( 
.A1(n_643),
.A2(n_603),
.B(n_579),
.C(n_618),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_645),
.B(n_587),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_642),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_646),
.Y(n_651)
);

NOR3x1_ASAP7_75t_L g652 ( 
.A(n_650),
.B(n_559),
.C(n_523),
.Y(n_652)
);

NOR2x1_ASAP7_75t_L g653 ( 
.A(n_648),
.B(n_647),
.Y(n_653)
);

NAND4xp75_ASAP7_75t_L g654 ( 
.A(n_653),
.B(n_649),
.C(n_510),
.D(n_572),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_651),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g656 ( 
.A(n_652),
.B(n_518),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_651),
.B(n_473),
.Y(n_657)
);

AND2x2_ASAP7_75t_SL g658 ( 
.A(n_655),
.B(n_505),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_657),
.Y(n_659)
);

NAND4xp75_ASAP7_75t_L g660 ( 
.A(n_654),
.B(n_510),
.C(n_572),
.D(n_487),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_656),
.B(n_505),
.Y(n_661)
);

NOR2x1_ASAP7_75t_L g662 ( 
.A(n_655),
.B(n_504),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_655),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_663),
.B(n_591),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_662),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_659),
.B(n_597),
.Y(n_666)
);

NAND3xp33_ASAP7_75t_SL g667 ( 
.A(n_660),
.B(n_542),
.C(n_545),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_658),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_661),
.A2(n_569),
.B1(n_547),
.B2(n_571),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_662),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_666),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_664),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_665),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_L g674 ( 
.A(n_670),
.B(n_538),
.Y(n_674)
);

OA22x2_ASAP7_75t_L g675 ( 
.A1(n_668),
.A2(n_588),
.B1(n_602),
.B2(n_601),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_673),
.A2(n_674),
.B1(n_675),
.B2(n_667),
.Y(n_676)
);

AO21x1_ASAP7_75t_L g677 ( 
.A1(n_672),
.A2(n_671),
.B(n_669),
.Y(n_677)
);

AOI31xp33_ASAP7_75t_L g678 ( 
.A1(n_673),
.A2(n_529),
.A3(n_528),
.B(n_537),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_673),
.A2(n_534),
.B(n_544),
.Y(n_679)
);

OAI221xp5_ASAP7_75t_L g680 ( 
.A1(n_673),
.A2(n_603),
.B1(n_525),
.B2(n_537),
.C(n_538),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_677),
.A2(n_571),
.B1(n_518),
.B2(n_547),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_676),
.Y(n_682)
);

AO22x2_ASAP7_75t_L g683 ( 
.A1(n_682),
.A2(n_679),
.B1(n_678),
.B2(n_680),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_681),
.A2(n_544),
.B1(n_598),
.B2(n_515),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_684),
.B(n_477),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_685),
.B(n_683),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_686),
.A2(n_477),
.B1(n_534),
.B2(n_504),
.Y(n_687)
);


endmodule