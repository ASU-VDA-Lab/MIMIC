module fake_netlist_1_6823_n_876 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_876);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_876;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_482;
wire n_394;
wire n_243;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_102), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_69), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_0), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_75), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_29), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_35), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_18), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_64), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_8), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_88), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_78), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_66), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_37), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_24), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_73), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_79), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_39), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_107), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_2), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_87), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_62), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_81), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_30), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_23), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_106), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_77), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_15), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_100), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_46), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_53), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_80), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_76), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_20), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_110), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_1), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_24), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_98), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_7), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_50), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g151 ( .A(n_40), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_92), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_34), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_67), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_136), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_136), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_123), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_154), .B(n_0), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_136), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_154), .B(n_1), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_146), .B(n_2), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_121), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_115), .Y(n_168) );
OR2x2_ASAP7_75t_L g169 ( .A(n_115), .B(n_3), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
AND2x6_ASAP7_75t_L g171 ( .A(n_121), .B(n_135), .Y(n_171) );
BUFx8_ASAP7_75t_SL g172 ( .A(n_116), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_124), .B(n_3), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
BUFx8_ASAP7_75t_L g175 ( .A(n_135), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_165), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_168), .B(n_124), .Y(n_179) );
AOI22xp5_ASAP7_75t_SL g180 ( .A1(n_172), .A2(n_116), .B1(n_151), .B2(n_130), .Y(n_180) );
OAI22xp33_ASAP7_75t_SL g181 ( .A1(n_169), .A2(n_153), .B1(n_113), .B2(n_117), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_168), .B(n_133), .Y(n_182) );
OAI22xp33_ASAP7_75t_SL g183 ( .A1(n_169), .A2(n_129), .B1(n_119), .B2(n_127), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_158), .A2(n_130), .B1(n_138), .B2(n_149), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g185 ( .A1(n_169), .A2(n_151), .B1(n_134), .B2(n_133), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_168), .B(n_144), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_169), .A2(n_134), .B1(n_147), .B2(n_123), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_165), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_158), .B(n_114), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_157), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g191 ( .A1(n_172), .A2(n_152), .B1(n_114), .B2(n_128), .Y(n_191) );
OA22x2_ASAP7_75t_L g192 ( .A1(n_158), .A2(n_152), .B1(n_139), .B2(n_120), .Y(n_192) );
OAI22xp33_ASAP7_75t_L g193 ( .A1(n_161), .A2(n_123), .B1(n_120), .B2(n_122), .Y(n_193) );
INVxp67_ASAP7_75t_SL g194 ( .A(n_161), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_161), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_174), .B(n_122), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_174), .B(n_171), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_158), .A2(n_123), .B1(n_128), .B2(n_137), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g201 ( .A1(n_173), .A2(n_123), .B1(n_137), .B2(n_139), .Y(n_201) );
AO22x2_ASAP7_75t_L g202 ( .A1(n_158), .A2(n_140), .B1(n_142), .B2(n_118), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_158), .A2(n_123), .B1(n_140), .B2(n_142), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_158), .A2(n_118), .B1(n_148), .B2(n_145), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_165), .B(n_111), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_157), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g209 ( .A1(n_173), .A2(n_150), .B1(n_143), .B2(n_141), .Y(n_209) );
OAI22xp5_ASAP7_75t_SL g210 ( .A1(n_173), .A2(n_132), .B1(n_131), .B2(n_126), .Y(n_210) );
AO22x2_ASAP7_75t_L g211 ( .A1(n_165), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_211) );
AO22x2_ASAP7_75t_L g212 ( .A1(n_165), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_165), .A2(n_125), .B1(n_112), .B2(n_9), .Y(n_213) );
AO22x2_ASAP7_75t_L g214 ( .A1(n_170), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_174), .B(n_10), .Y(n_215) );
BUFx10_ASAP7_75t_L g216 ( .A(n_171), .Y(n_216) );
AO22x2_ASAP7_75t_L g217 ( .A1(n_170), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_217) );
OA22x2_ASAP7_75t_L g218 ( .A1(n_170), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_175), .B(n_45), .Y(n_219) );
INVx2_ASAP7_75t_SL g220 ( .A(n_175), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_174), .B(n_13), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_175), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_166), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_178), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_195), .B(n_174), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_180), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_194), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_200), .A2(n_171), .B(n_159), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_184), .Y(n_229) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_220), .B(n_175), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_178), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_202), .B(n_177), .Y(n_232) );
INVxp33_ASAP7_75t_L g233 ( .A(n_186), .Y(n_233) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_189), .B(n_157), .Y(n_234) );
CKINVDCx14_ASAP7_75t_R g235 ( .A(n_184), .Y(n_235) );
XOR2xp5_ASAP7_75t_L g236 ( .A(n_213), .B(n_14), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_178), .Y(n_237) );
BUFx2_ASAP7_75t_R g238 ( .A(n_222), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_188), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_188), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_207), .B(n_175), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_198), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_207), .B(n_175), .Y(n_243) );
NOR2xp33_ASAP7_75t_SL g244 ( .A(n_220), .B(n_175), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_202), .B(n_177), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_189), .B(n_171), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_198), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_189), .Y(n_248) );
NOR2xp33_ASAP7_75t_SL g249 ( .A(n_222), .B(n_171), .Y(n_249) );
INVxp33_ASAP7_75t_SL g250 ( .A(n_210), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_202), .B(n_177), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_202), .B(n_171), .Y(n_252) );
INVxp33_ASAP7_75t_L g253 ( .A(n_179), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
XNOR2x2_ASAP7_75t_L g255 ( .A(n_214), .B(n_159), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_200), .B(n_171), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_192), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_192), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_192), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_179), .B(n_171), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_203), .A2(n_171), .B(n_162), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_190), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_215), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_182), .B(n_171), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_190), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_221), .Y(n_267) );
XOR2xp5_ASAP7_75t_L g268 ( .A(n_213), .B(n_14), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_221), .Y(n_269) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_191), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_209), .B(n_157), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_199), .Y(n_272) );
XOR2xp5_ASAP7_75t_L g273 ( .A(n_185), .B(n_15), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_199), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_182), .B(n_171), .Y(n_275) );
NAND2xp33_ASAP7_75t_R g276 ( .A(n_197), .B(n_16), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_206), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_203), .B(n_171), .Y(n_278) );
INVxp67_ASAP7_75t_SL g279 ( .A(n_223), .Y(n_279) );
NOR2xp67_ASAP7_75t_L g280 ( .A(n_206), .B(n_166), .Y(n_280) );
NOR2xp67_ASAP7_75t_L g281 ( .A(n_196), .B(n_166), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_211), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_216), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_219), .B(n_171), .Y(n_284) );
INVxp33_ASAP7_75t_L g285 ( .A(n_211), .Y(n_285) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_227), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_227), .B(n_187), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_234), .B(n_211), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_234), .B(n_211), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_260), .B(n_166), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_225), .B(n_181), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_224), .Y(n_292) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_239), .A2(n_204), .B(n_205), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_231), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_225), .B(n_183), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_234), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_233), .B(n_193), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_225), .B(n_212), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_231), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_239), .B(n_201), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_240), .B(n_212), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_240), .B(n_212), .Y(n_302) );
BUFx5_ASAP7_75t_L g303 ( .A(n_232), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_237), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_252), .A2(n_218), .B(n_163), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_253), .B(n_204), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_237), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_224), .Y(n_308) );
INVx4_ASAP7_75t_L g309 ( .A(n_252), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_260), .B(n_205), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_242), .B(n_212), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_260), .B(n_214), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_224), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_242), .B(n_214), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_224), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_247), .B(n_214), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_224), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_265), .B(n_217), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_282), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_262), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_262), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_229), .B(n_16), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_282), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_265), .B(n_166), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_265), .B(n_166), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_248), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_248), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_247), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_254), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_262), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_266), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_266), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_275), .B(n_254), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_266), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_272), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_275), .B(n_217), .Y(n_336) );
INVx4_ASAP7_75t_L g337 ( .A(n_323), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_286), .B(n_263), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_321), .Y(n_339) );
AND2x6_ASAP7_75t_L g340 ( .A(n_323), .B(n_252), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_286), .B(n_263), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_323), .B(n_319), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_291), .B(n_277), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_328), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_323), .B(n_279), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_335), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_335), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
OR2x6_ASAP7_75t_L g349 ( .A(n_288), .B(n_264), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_303), .B(n_275), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_303), .B(n_264), .Y(n_351) );
INVx4_ASAP7_75t_L g352 ( .A(n_296), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_322), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_328), .B(n_267), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_328), .B(n_267), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_296), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_329), .B(n_269), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_321), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_303), .B(n_269), .Y(n_360) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_335), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_329), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_319), .Y(n_364) );
NOR2xp33_ASAP7_75t_SL g365 ( .A(n_319), .B(n_230), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_333), .B(n_279), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_303), .B(n_257), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_346), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_337), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_337), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_337), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_289), .B1(n_288), .B2(n_273), .Y(n_373) );
INVx5_ASAP7_75t_SL g374 ( .A(n_345), .Y(n_374) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_346), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_347), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_353), .A2(n_289), .B1(n_288), .B2(n_273), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
NOR2xp67_ASAP7_75t_SL g379 ( .A(n_337), .B(n_288), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_339), .Y(n_380) );
BUFx6f_ASAP7_75t_SL g381 ( .A(n_345), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_361), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_339), .Y(n_383) );
INVx8_ASAP7_75t_L g384 ( .A(n_340), .Y(n_384) );
INVx3_ASAP7_75t_SL g385 ( .A(n_337), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_361), .Y(n_386) );
INVx8_ASAP7_75t_L g387 ( .A(n_340), .Y(n_387) );
OR2x6_ASAP7_75t_L g388 ( .A(n_349), .B(n_289), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_337), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_344), .Y(n_391) );
INVx4_ASAP7_75t_L g392 ( .A(n_345), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_348), .Y(n_393) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_348), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_351), .B(n_289), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_339), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_342), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_385), .Y(n_398) );
CKINVDCx11_ASAP7_75t_R g399 ( .A(n_385), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_385), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_380), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_389), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_381), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_381), .A2(n_235), .B1(n_236), .B2(n_268), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_385), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_373), .A2(n_322), .B1(n_285), .B2(n_364), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_397), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_380), .Y(n_408) );
BUFx10_ASAP7_75t_L g409 ( .A(n_381), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_389), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_373), .A2(n_342), .B1(n_322), .B2(n_345), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_391), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_377), .A2(n_342), .B1(n_322), .B2(n_345), .Y(n_413) );
BUFx10_ASAP7_75t_L g414 ( .A(n_381), .Y(n_414) );
INVx4_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_377), .B(n_343), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_392), .A2(n_235), .B1(n_268), .B2(n_236), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_374), .A2(n_342), .B1(n_345), .B2(n_364), .Y(n_418) );
BUFx4_ASAP7_75t_SL g419 ( .A(n_397), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_391), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_397), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_380), .Y(n_422) );
CKINVDCx11_ASAP7_75t_R g423 ( .A(n_384), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_375), .A2(n_343), .B1(n_367), .B2(n_298), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_383), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_395), .B(n_339), .Y(n_426) );
INVx2_ASAP7_75t_SL g427 ( .A(n_371), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_383), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_375), .A2(n_367), .B1(n_298), .B2(n_349), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_383), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_392), .A2(n_367), .B1(n_298), .B2(n_349), .Y(n_431) );
CKINVDCx11_ASAP7_75t_R g432 ( .A(n_384), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_392), .A2(n_367), .B1(n_298), .B2(n_349), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_392), .A2(n_349), .B1(n_296), .B2(n_226), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_384), .A2(n_364), .B1(n_340), .B2(n_255), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_392), .B(n_352), .Y(n_436) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_384), .A2(n_340), .B1(n_255), .B2(n_342), .Y(n_437) );
OAI22xp33_ASAP7_75t_SL g438 ( .A1(n_370), .A2(n_349), .B1(n_365), .B2(n_352), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_395), .B(n_359), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_384), .A2(n_340), .B1(n_255), .B2(n_365), .Y(n_440) );
INVx6_ASAP7_75t_L g441 ( .A(n_371), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_404), .B(n_250), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_422), .Y(n_443) );
INVx5_ASAP7_75t_SL g444 ( .A(n_419), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_406), .A2(n_388), .B1(n_379), .B2(n_384), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_411), .A2(n_367), .B1(n_379), .B2(n_217), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_417), .A2(n_370), .B(n_390), .Y(n_447) );
AOI22xp33_ASAP7_75t_SL g448 ( .A1(n_413), .A2(n_374), .B1(n_387), .B2(n_384), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_422), .B(n_374), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_431), .A2(n_374), .B1(n_388), .B2(n_370), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_416), .B(n_270), .Y(n_451) );
OAI22xp33_ASAP7_75t_L g452 ( .A1(n_415), .A2(n_388), .B1(n_387), .B2(n_349), .Y(n_452) );
INVx4_ASAP7_75t_L g453 ( .A(n_409), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_402), .Y(n_454) );
AOI22xp33_ASAP7_75t_SL g455 ( .A1(n_415), .A2(n_438), .B1(n_400), .B2(n_403), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_421), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_399), .A2(n_388), .B1(n_379), .B2(n_387), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g458 ( .A1(n_415), .A2(n_438), .B1(n_400), .B2(n_403), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_421), .Y(n_459) );
NOR2x1_ASAP7_75t_L g460 ( .A(n_415), .B(n_371), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_426), .B(n_395), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_402), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_434), .B(n_291), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_410), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_435), .A2(n_388), .B1(n_387), .B2(n_340), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_437), .A2(n_388), .B1(n_387), .B2(n_340), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_440), .A2(n_388), .B1(n_387), .B2(n_340), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_410), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_412), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_436), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_401), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_409), .Y(n_472) );
OAI21xp5_ASAP7_75t_SL g473 ( .A1(n_418), .A2(n_390), .B(n_367), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_412), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_431), .A2(n_374), .B1(n_390), .B2(n_372), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_401), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_408), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_426), .B(n_396), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_439), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_409), .Y(n_480) );
OAI22xp5_ASAP7_75t_SL g481 ( .A1(n_433), .A2(n_372), .B1(n_369), .B2(n_376), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_433), .A2(n_372), .B1(n_396), .B2(n_238), .Y(n_482) );
OR2x2_ASAP7_75t_SL g483 ( .A(n_441), .B(n_369), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_408), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_420), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_424), .A2(n_340), .B1(n_309), .B2(n_296), .Y(n_486) );
OAI222xp33_ASAP7_75t_L g487 ( .A1(n_436), .A2(n_386), .B1(n_382), .B2(n_378), .C1(n_376), .C2(n_218), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_409), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_420), .Y(n_489) );
AOI222xp33_ASAP7_75t_L g490 ( .A1(n_423), .A2(n_295), .B1(n_291), .B2(n_217), .C1(n_297), .C2(n_318), .Y(n_490) );
BUFx3_ASAP7_75t_L g491 ( .A(n_436), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_429), .A2(n_238), .B1(n_386), .B2(n_382), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_414), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_429), .A2(n_378), .B1(n_344), .B2(n_354), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_398), .Y(n_495) );
INVx3_ASAP7_75t_L g496 ( .A(n_414), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_425), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_441), .B(n_295), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_441), .B(n_295), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_439), .A2(n_340), .B1(n_309), .B2(n_296), .Y(n_500) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_414), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g502 ( .A1(n_405), .A2(n_354), .B1(n_356), .B2(n_338), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_425), .B(n_359), .Y(n_503) );
BUFx4f_ASAP7_75t_SL g504 ( .A(n_414), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_427), .B(n_245), .C(n_232), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_407), .A2(n_309), .B1(n_218), .B2(n_338), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_432), .A2(n_309), .B1(n_296), .B2(n_336), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_441), .A2(n_309), .B1(n_296), .B2(n_336), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_427), .A2(n_309), .B1(n_296), .B2(n_336), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_407), .A2(n_312), .B1(n_336), .B2(n_318), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_407), .B(n_393), .Y(n_511) );
AOI222xp33_ASAP7_75t_L g512 ( .A1(n_428), .A2(n_297), .B1(n_318), .B2(n_312), .C1(n_351), .C2(n_360), .Y(n_512) );
OAI221xp5_ASAP7_75t_L g513 ( .A1(n_442), .A2(n_341), .B1(n_280), .B2(n_358), .C(n_356), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_492), .A2(n_312), .B1(n_303), .B2(n_352), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_454), .B(n_430), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_482), .A2(n_303), .B1(n_352), .B2(n_296), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_490), .A2(n_448), .B1(n_450), .B2(n_481), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_481), .A2(n_303), .B1(n_352), .B2(n_280), .Y(n_518) );
OAI222xp33_ASAP7_75t_L g519 ( .A1(n_446), .A2(n_430), .B1(n_352), .B2(n_314), .C1(n_316), .C2(n_311), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_446), .A2(n_341), .B1(n_351), .B2(n_360), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_463), .A2(n_303), .B1(n_245), .B2(n_251), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_445), .A2(n_303), .B1(n_251), .B2(n_232), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_473), .A2(n_302), .B(n_311), .C(n_301), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_494), .A2(n_465), .B1(n_466), .B2(n_510), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_502), .A2(n_302), .B(n_301), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_452), .A2(n_303), .B1(n_360), .B2(n_363), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_512), .A2(n_303), .B1(n_363), .B2(n_366), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_444), .A2(n_303), .B1(n_394), .B2(n_393), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_486), .A2(n_316), .B1(n_314), .B2(n_302), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_467), .A2(n_303), .B1(n_366), .B2(n_363), .Y(n_530) );
OAI222xp33_ASAP7_75t_L g531 ( .A1(n_455), .A2(n_311), .B1(n_357), .B2(n_366), .C1(n_358), .C2(n_359), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_443), .Y(n_532) );
OAI222xp33_ASAP7_75t_L g533 ( .A1(n_458), .A2(n_357), .B1(n_359), .B2(n_368), .C1(n_287), .C2(n_350), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_444), .A2(n_303), .B1(n_393), .B2(n_394), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_451), .A2(n_303), .B1(n_350), .B2(n_368), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_498), .A2(n_350), .B1(n_393), .B2(n_394), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_499), .A2(n_394), .B1(n_393), .B2(n_305), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_479), .B(n_305), .Y(n_538) );
OAI22xp33_ASAP7_75t_L g539 ( .A1(n_504), .A2(n_276), .B1(n_394), .B2(n_393), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_475), .A2(n_394), .B1(n_393), .B2(n_305), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_487), .B(n_160), .C(n_159), .Y(n_541) );
INVxp67_ASAP7_75t_L g542 ( .A(n_456), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_454), .B(n_393), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_505), .A2(n_394), .B1(n_305), .B2(n_284), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_505), .A2(n_394), .B1(n_284), .B2(n_307), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_457), .A2(n_284), .B1(n_307), .B2(n_299), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_500), .A2(n_284), .B1(n_307), .B2(n_299), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_507), .A2(n_284), .B1(n_304), .B2(n_294), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_444), .A2(n_304), .B1(n_299), .B2(n_294), .Y(n_549) );
AOI222xp33_ASAP7_75t_L g550 ( .A1(n_444), .A2(n_259), .B1(n_258), .B2(n_257), .C1(n_287), .C2(n_306), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_508), .A2(n_304), .B1(n_294), .B2(n_243), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_447), .A2(n_287), .B1(n_355), .B2(n_348), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_506), .A2(n_276), .B1(n_241), .B2(n_243), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_491), .A2(n_241), .B1(n_333), .B2(n_259), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_462), .B(n_17), .Y(n_555) );
OAI222xp33_ASAP7_75t_L g556 ( .A1(n_453), .A2(n_258), .B1(n_332), .B2(n_321), .C1(n_331), .C2(n_160), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_462), .B(n_17), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_491), .A2(n_333), .B1(n_271), .B2(n_290), .Y(n_558) );
AOI221xp5_ASAP7_75t_SL g559 ( .A1(n_483), .A2(n_176), .B1(n_162), .B2(n_159), .C(n_160), .Y(n_559) );
AOI222xp33_ASAP7_75t_L g560 ( .A1(n_461), .A2(n_306), .B1(n_333), .B2(n_300), .C1(n_271), .C2(n_228), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_459), .A2(n_333), .B1(n_290), .B2(n_324), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_470), .A2(n_333), .B1(n_290), .B2(n_324), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_453), .A2(n_333), .B1(n_321), .B2(n_332), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_464), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_483), .A2(n_362), .B1(n_355), .B2(n_348), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_509), .A2(n_325), .B1(n_324), .B2(n_290), .Y(n_566) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_464), .A2(n_300), .B1(n_228), .B2(n_261), .C1(n_278), .C2(n_293), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_460), .A2(n_290), .B1(n_324), .B2(n_325), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_460), .A2(n_290), .B1(n_324), .B2(n_325), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_468), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_453), .A2(n_325), .B1(n_324), .B2(n_300), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_480), .A2(n_362), .B1(n_355), .B2(n_348), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_480), .A2(n_355), .B1(n_348), .B2(n_362), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_478), .A2(n_325), .B1(n_320), .B2(n_330), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_449), .A2(n_362), .B1(n_355), .B2(n_348), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_478), .A2(n_325), .B1(n_320), .B2(n_330), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_468), .A2(n_320), .B1(n_330), .B2(n_334), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_501), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_469), .A2(n_320), .B1(n_330), .B2(n_334), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_449), .A2(n_362), .B1(n_355), .B2(n_348), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_469), .B(n_159), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_480), .A2(n_362), .B1(n_355), .B2(n_348), .Y(n_582) );
INVx4_ASAP7_75t_L g583 ( .A(n_501), .Y(n_583) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_474), .A2(n_261), .B1(n_278), .B2(n_293), .C1(n_332), .C2(n_331), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_493), .A2(n_355), .B1(n_362), .B2(n_332), .Y(n_585) );
OAI221xp5_ASAP7_75t_L g586 ( .A1(n_495), .A2(n_163), .B1(n_162), .B2(n_160), .C(n_310), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_474), .B(n_18), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_485), .B(n_160), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_485), .B(n_489), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_489), .A2(n_330), .B1(n_320), .B2(n_334), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_472), .A2(n_330), .B1(n_320), .B2(n_334), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_472), .A2(n_330), .B1(n_320), .B2(n_334), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_488), .A2(n_330), .B1(n_334), .B2(n_355), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_488), .A2(n_162), .B1(n_163), .B2(n_310), .C(n_293), .Y(n_594) );
OAI21xp5_ASAP7_75t_SL g595 ( .A1(n_493), .A2(n_278), .B(n_331), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_493), .A2(n_330), .B1(n_362), .B2(n_315), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_501), .B(n_362), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_496), .A2(n_330), .B1(n_313), .B2(n_292), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_496), .A2(n_331), .B1(n_308), .B2(n_317), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_496), .A2(n_292), .B1(n_315), .B2(n_313), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_501), .A2(n_292), .B1(n_315), .B2(n_313), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_503), .B(n_19), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_443), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_511), .A2(n_317), .B1(n_308), .B2(n_327), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_471), .B(n_162), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_471), .B(n_163), .C(n_156), .Y(n_606) );
OAI22xp33_ASAP7_75t_L g607 ( .A1(n_476), .A2(n_230), .B1(n_244), .B2(n_256), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_511), .A2(n_317), .B1(n_308), .B2(n_327), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_542), .B(n_163), .C(n_176), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_515), .B(n_477), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_543), .B(n_477), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_565), .B(n_484), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_543), .B(n_497), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_517), .A2(n_176), .B(n_156), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_565), .B(n_166), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_524), .A2(n_176), .B1(n_156), .B2(n_164), .C(n_155), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_564), .B(n_19), .Y(n_617) );
NOR3xp33_ASAP7_75t_SL g618 ( .A(n_524), .B(n_256), .C(n_246), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_520), .A2(n_167), .B1(n_166), .B2(n_327), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_559), .B(n_176), .C(n_156), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_513), .A2(n_176), .B1(n_156), .B2(n_164), .C(n_155), .Y(n_621) );
OAI21xp5_ASAP7_75t_SL g622 ( .A1(n_595), .A2(n_176), .B(n_21), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_532), .B(n_155), .Y(n_623) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_559), .B(n_176), .C(n_156), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_532), .B(n_155), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_531), .B(n_20), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_570), .B(n_21), .Y(n_627) );
AOI211xp5_ASAP7_75t_L g628 ( .A1(n_595), .A2(n_155), .B(n_156), .C(n_164), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_570), .B(n_22), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_589), .B(n_22), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_555), .B(n_246), .C(n_326), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g632 ( .A(n_557), .B(n_155), .C(n_156), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_578), .B(n_23), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_520), .B(n_25), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_578), .B(n_25), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_587), .B(n_155), .C(n_164), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_603), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_583), .B(n_552), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_541), .B(n_155), .C(n_164), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_603), .B(n_26), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_516), .B(n_155), .C(n_164), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_518), .B(n_164), .C(n_166), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_540), .B(n_164), .Y(n_643) );
OAI221xp5_ASAP7_75t_SL g644 ( .A1(n_514), .A2(n_26), .B1(n_27), .B2(n_28), .C(n_29), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_549), .A2(n_166), .B1(n_167), .B2(n_164), .C(n_244), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_550), .A2(n_164), .B1(n_326), .B2(n_327), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_553), .A2(n_166), .B(n_167), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_581), .B(n_30), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_583), .B(n_31), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_588), .B(n_31), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_583), .B(n_32), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_525), .B(n_32), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_525), .B(n_33), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_563), .A2(n_167), .B1(n_326), .B2(n_327), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_536), .B(n_34), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_528), .B(n_167), .C(n_249), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_538), .B(n_35), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_605), .B(n_36), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_572), .B(n_167), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_534), .B(n_167), .C(n_249), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_605), .B(n_36), .Y(n_661) );
OAI221xp5_ASAP7_75t_SL g662 ( .A1(n_527), .A2(n_526), .B1(n_523), .B2(n_530), .C(n_550), .Y(n_662) );
OAI21xp33_ASAP7_75t_SL g663 ( .A1(n_597), .A2(n_37), .B(n_38), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_537), .B(n_38), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_575), .B(n_39), .Y(n_665) );
NAND4xp25_ASAP7_75t_L g666 ( .A(n_560), .B(n_281), .C(n_41), .D(n_42), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_602), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_575), .B(n_40), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_580), .B(n_41), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_580), .B(n_42), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_582), .B(n_43), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_529), .B(n_43), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_582), .B(n_167), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_563), .A2(n_326), .B1(n_327), .B2(n_167), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_584), .B(n_167), .C(n_274), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_574), .B(n_44), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_529), .B(n_44), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_584), .B(n_47), .Y(n_678) );
OA21x2_ASAP7_75t_L g679 ( .A1(n_533), .A2(n_274), .B(n_272), .Y(n_679) );
OAI22xp5_ASAP7_75t_SL g680 ( .A1(n_568), .A2(n_326), .B1(n_49), .B2(n_51), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_569), .A2(n_326), .B1(n_274), .B2(n_272), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_576), .B(n_48), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_521), .B(n_52), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_553), .B(n_54), .C(n_55), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_535), .A2(n_522), .B1(n_558), .B2(n_561), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_519), .A2(n_208), .B1(n_57), .B2(n_58), .C(n_59), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g687 ( .A1(n_546), .A2(n_56), .B1(n_60), .B2(n_61), .C(n_63), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_573), .B(n_65), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_544), .B(n_585), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_567), .B(n_68), .Y(n_690) );
OAI221xp5_ASAP7_75t_SL g691 ( .A1(n_571), .A2(n_70), .B1(n_71), .B2(n_72), .C(n_74), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_567), .B(n_83), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_586), .B(n_84), .C(n_85), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_577), .B(n_86), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_599), .B(n_89), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_545), .A2(n_90), .B1(n_91), .B2(n_93), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_599), .B(n_94), .Y(n_697) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_539), .A2(n_95), .B(n_96), .Y(n_698) );
AND2x2_ASAP7_75t_SL g699 ( .A(n_596), .B(n_97), .Y(n_699) );
NAND4xp25_ASAP7_75t_L g700 ( .A(n_554), .B(n_99), .C(n_101), .D(n_103), .Y(n_700) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_606), .B(n_104), .C(n_105), .Y(n_701) );
AOI22xp33_ASAP7_75t_SL g702 ( .A1(n_594), .A2(n_108), .B1(n_109), .B2(n_216), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_579), .B(n_208), .Y(n_703) );
INVxp67_ASAP7_75t_SL g704 ( .A(n_637), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_614), .A2(n_548), .B1(n_547), .B2(n_551), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_666), .B(n_556), .C(n_606), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_616), .B(n_593), .C(n_592), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_622), .B(n_591), .C(n_598), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g709 ( .A1(n_663), .A2(n_607), .B(n_562), .C(n_566), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_667), .B(n_600), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_611), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_630), .B(n_608), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g713 ( .A(n_618), .B(n_590), .C(n_601), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_657), .B(n_604), .Y(n_714) );
NOR2xp33_ASAP7_75t_SL g715 ( .A(n_699), .B(n_283), .Y(n_715) );
INVxp67_ASAP7_75t_L g716 ( .A(n_649), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_613), .B(n_283), .Y(n_717) );
INVxp67_ASAP7_75t_SL g718 ( .A(n_612), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_628), .B(n_283), .C(n_638), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_652), .B(n_283), .Y(n_720) );
NOR3xp33_ASAP7_75t_L g721 ( .A(n_644), .B(n_283), .C(n_700), .Y(n_721) );
AO21x2_ASAP7_75t_L g722 ( .A1(n_617), .A2(n_627), .B(n_629), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_653), .B(n_634), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_658), .B(n_661), .Y(n_724) );
INVx2_ASAP7_75t_SL g725 ( .A(n_649), .Y(n_725) );
OR2x2_ASAP7_75t_SL g726 ( .A(n_679), .B(n_675), .Y(n_726) );
NOR3xp33_ASAP7_75t_L g727 ( .A(n_691), .B(n_684), .C(n_651), .Y(n_727) );
NOR3xp33_ASAP7_75t_L g728 ( .A(n_672), .B(n_677), .C(n_621), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_689), .B(n_643), .Y(n_729) );
AO21x2_ASAP7_75t_L g730 ( .A1(n_623), .A2(n_625), .B(n_615), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_649), .B(n_615), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_689), .B(n_633), .Y(n_732) );
AOI22xp33_ASAP7_75t_SL g733 ( .A1(n_679), .A2(n_670), .B1(n_665), .B2(n_671), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_635), .B(n_640), .Y(n_734) );
NOR3xp33_ASAP7_75t_SL g735 ( .A(n_662), .B(n_680), .C(n_690), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_643), .B(n_625), .Y(n_736) );
NAND4xp75_ASAP7_75t_L g737 ( .A(n_665), .B(n_670), .C(n_679), .D(n_671), .Y(n_737) );
NAND4xp75_ASAP7_75t_L g738 ( .A(n_668), .B(n_669), .C(n_664), .D(n_692), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_685), .A2(n_631), .B1(n_646), .B2(n_664), .Y(n_739) );
NAND4xp75_ASAP7_75t_L g740 ( .A(n_686), .B(n_678), .C(n_650), .D(n_648), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_685), .A2(n_646), .B1(n_655), .B2(n_676), .Y(n_741) );
OA211x2_ASAP7_75t_L g742 ( .A1(n_673), .A2(n_659), .B(n_695), .C(n_647), .Y(n_742) );
AO21x2_ASAP7_75t_L g743 ( .A1(n_632), .A2(n_636), .B(n_698), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_688), .B(n_676), .Y(n_744) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_687), .B(n_642), .C(n_609), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_694), .B(n_697), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_694), .B(n_620), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_624), .B(n_619), .Y(n_748) );
INVxp67_ASAP7_75t_SL g749 ( .A(n_639), .Y(n_749) );
AO21x2_ASAP7_75t_L g750 ( .A1(n_693), .A2(n_641), .B(n_701), .Y(n_750) );
NOR3xp33_ASAP7_75t_L g751 ( .A(n_696), .B(n_656), .C(n_660), .Y(n_751) );
BUFx2_ASAP7_75t_L g752 ( .A(n_682), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_674), .B(n_703), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_654), .Y(n_754) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_702), .B(n_683), .C(n_645), .Y(n_755) );
AO21x2_ASAP7_75t_L g756 ( .A1(n_681), .A2(n_638), .B(n_627), .Y(n_756) );
NOR2x1_ASAP7_75t_L g757 ( .A(n_649), .B(n_622), .Y(n_757) );
NAND4xp75_ASAP7_75t_L g758 ( .A(n_699), .B(n_618), .C(n_651), .D(n_616), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g759 ( .A(n_616), .B(n_622), .C(n_618), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_637), .Y(n_760) );
OR2x2_ASAP7_75t_L g761 ( .A(n_637), .B(n_610), .Y(n_761) );
OR2x2_ASAP7_75t_L g762 ( .A(n_637), .B(n_610), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_638), .B(n_565), .Y(n_763) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_637), .Y(n_764) );
OA211x2_ASAP7_75t_L g765 ( .A1(n_638), .A2(n_626), .B(n_614), .C(n_615), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_667), .B(n_542), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_667), .B(n_610), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_735), .B(n_719), .C(n_757), .Y(n_768) );
XOR2x2_ASAP7_75t_L g769 ( .A(n_738), .B(n_740), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g770 ( .A(n_735), .B(n_728), .C(n_706), .Y(n_770) );
INVx2_ASAP7_75t_SL g771 ( .A(n_760), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_729), .B(n_732), .Y(n_772) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_760), .Y(n_773) );
INVx2_ASAP7_75t_L g774 ( .A(n_764), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_764), .Y(n_775) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_704), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_761), .B(n_762), .Y(n_777) );
NAND4xp75_ASAP7_75t_SL g778 ( .A(n_747), .B(n_765), .C(n_729), .D(n_723), .Y(n_778) );
XNOR2xp5_ASAP7_75t_L g779 ( .A(n_734), .B(n_741), .Y(n_779) );
XNOR2x2_ASAP7_75t_L g780 ( .A(n_737), .B(n_763), .Y(n_780) );
NAND4xp75_ASAP7_75t_SL g781 ( .A(n_747), .B(n_723), .C(n_715), .D(n_726), .Y(n_781) );
NAND4xp75_ASAP7_75t_SL g782 ( .A(n_712), .B(n_714), .C(n_746), .D(n_753), .Y(n_782) );
INVx5_ASAP7_75t_L g783 ( .A(n_731), .Y(n_783) );
NOR4xp25_ASAP7_75t_L g784 ( .A(n_766), .B(n_741), .C(n_763), .D(n_739), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_711), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_767), .B(n_766), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_742), .A2(n_727), .B1(n_754), .B2(n_751), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_718), .B(n_716), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_725), .B(n_724), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_730), .Y(n_790) );
BUFx2_ASAP7_75t_L g791 ( .A(n_725), .Y(n_791) );
OR2x2_ASAP7_75t_L g792 ( .A(n_730), .B(n_756), .Y(n_792) );
NAND4xp75_ASAP7_75t_SL g793 ( .A(n_712), .B(n_714), .C(n_746), .D(n_753), .Y(n_793) );
BUFx2_ASAP7_75t_L g794 ( .A(n_731), .Y(n_794) );
XNOR2x2_ASAP7_75t_L g795 ( .A(n_758), .B(n_759), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_739), .A2(n_733), .B1(n_731), .B2(n_710), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_722), .B(n_756), .Y(n_797) );
INVx3_ASAP7_75t_L g798 ( .A(n_736), .Y(n_798) );
OR2x2_ASAP7_75t_L g799 ( .A(n_722), .B(n_736), .Y(n_799) );
NAND4xp75_ASAP7_75t_SL g800 ( .A(n_744), .B(n_710), .C(n_717), .D(n_720), .Y(n_800) );
NOR4xp25_ASAP7_75t_L g801 ( .A(n_708), .B(n_748), .C(n_749), .D(n_755), .Y(n_801) );
OR2x2_ASAP7_75t_L g802 ( .A(n_717), .B(n_752), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_743), .Y(n_803) );
AND2x2_ASAP7_75t_L g804 ( .A(n_743), .B(n_720), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_707), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_709), .B(n_750), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_750), .B(n_745), .Y(n_807) );
XNOR2xp5_ASAP7_75t_L g808 ( .A(n_769), .B(n_705), .Y(n_808) );
XOR2x2_ASAP7_75t_L g809 ( .A(n_769), .B(n_721), .Y(n_809) );
XOR2x2_ASAP7_75t_L g810 ( .A(n_770), .B(n_713), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_776), .Y(n_811) );
XNOR2x1_ASAP7_75t_L g812 ( .A(n_795), .B(n_770), .Y(n_812) );
AND2x2_ASAP7_75t_SL g813 ( .A(n_784), .B(n_801), .Y(n_813) );
OR2x2_ASAP7_75t_L g814 ( .A(n_799), .B(n_777), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_802), .Y(n_815) );
INVxp67_ASAP7_75t_L g816 ( .A(n_797), .Y(n_816) );
XNOR2x2_ASAP7_75t_L g817 ( .A(n_795), .B(n_780), .Y(n_817) );
INVx2_ASAP7_75t_SL g818 ( .A(n_777), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_805), .B(n_806), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_805), .B(n_806), .Y(n_820) );
INVxp67_ASAP7_75t_L g821 ( .A(n_804), .Y(n_821) );
XNOR2x1_ASAP7_75t_L g822 ( .A(n_778), .B(n_779), .Y(n_822) );
AO22x2_ASAP7_75t_L g823 ( .A1(n_768), .A2(n_792), .B1(n_807), .B2(n_799), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_773), .Y(n_824) );
INVx1_ASAP7_75t_SL g825 ( .A(n_771), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_785), .Y(n_826) );
XNOR2xp5_ASAP7_75t_L g827 ( .A(n_782), .B(n_793), .Y(n_827) );
XNOR2x1_ASAP7_75t_L g828 ( .A(n_779), .B(n_780), .Y(n_828) );
INVx2_ASAP7_75t_SL g829 ( .A(n_783), .Y(n_829) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_828), .A2(n_768), .B1(n_796), .B2(n_787), .Y(n_830) );
AOI22x1_ASAP7_75t_L g831 ( .A1(n_827), .A2(n_807), .B1(n_792), .B2(n_801), .Y(n_831) );
INVxp67_ASAP7_75t_L g832 ( .A(n_817), .Y(n_832) );
OA22x2_ASAP7_75t_L g833 ( .A1(n_808), .A2(n_796), .B1(n_794), .B2(n_804), .Y(n_833) );
AOI22xp5_ASAP7_75t_SL g834 ( .A1(n_829), .A2(n_794), .B1(n_791), .B2(n_781), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_811), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_818), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_826), .Y(n_837) );
AO22x2_ASAP7_75t_L g838 ( .A1(n_812), .A2(n_803), .B1(n_800), .B2(n_790), .Y(n_838) );
OA22x2_ASAP7_75t_L g839 ( .A1(n_821), .A2(n_788), .B1(n_772), .B2(n_789), .Y(n_839) );
OA22x2_ASAP7_75t_L g840 ( .A1(n_821), .A2(n_788), .B1(n_789), .B2(n_798), .Y(n_840) );
INVx1_ASAP7_75t_SL g841 ( .A(n_825), .Y(n_841) );
OA22x2_ASAP7_75t_L g842 ( .A1(n_812), .A2(n_798), .B1(n_775), .B2(n_774), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_815), .Y(n_843) );
AO22x1_ASAP7_75t_L g844 ( .A1(n_819), .A2(n_783), .B1(n_798), .B2(n_786), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_837), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_835), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_836), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_841), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_843), .Y(n_849) );
INVx1_ASAP7_75t_SL g850 ( .A(n_834), .Y(n_850) );
NOR2x1_ASAP7_75t_L g851 ( .A(n_837), .B(n_822), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_832), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_848), .Y(n_853) );
INVxp67_ASAP7_75t_L g854 ( .A(n_852), .Y(n_854) );
OAI222xp33_ASAP7_75t_L g855 ( .A1(n_850), .A2(n_833), .B1(n_831), .B2(n_830), .C1(n_842), .C2(n_840), .Y(n_855) );
OA22x2_ASAP7_75t_L g856 ( .A1(n_847), .A2(n_813), .B1(n_831), .B2(n_809), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_845), .Y(n_857) );
AOI31xp33_ASAP7_75t_L g858 ( .A1(n_854), .A2(n_851), .A3(n_820), .B(n_819), .Y(n_858) );
AOI221xp5_ASAP7_75t_L g859 ( .A1(n_855), .A2(n_823), .B1(n_820), .B2(n_838), .C(n_846), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_853), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_860), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_858), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_861), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_861), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_863), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_864), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_865), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_866), .A2(n_856), .B1(n_862), .B2(n_810), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_868), .A2(n_856), .B1(n_859), .B2(n_813), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_869), .Y(n_870) );
AOI211xp5_ASAP7_75t_L g871 ( .A1(n_870), .A2(n_867), .B(n_857), .C(n_844), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_871), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_872), .A2(n_849), .B1(n_839), .B2(n_816), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_873), .Y(n_874) );
AOI221xp5_ASAP7_75t_L g875 ( .A1(n_874), .A2(n_823), .B1(n_816), .B2(n_845), .C(n_838), .Y(n_875) );
AOI211xp5_ASAP7_75t_L g876 ( .A1(n_875), .A2(n_825), .B(n_814), .C(n_824), .Y(n_876) );
endmodule