module real_jpeg_6395_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_525;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_0),
.A2(n_151),
.B1(n_154),
.B2(n_157),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_0),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_0),
.B(n_174),
.C(n_177),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_0),
.B(n_79),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_0),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_0),
.B(n_168),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_0),
.B(n_267),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_1),
.Y(n_193)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_1),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_1),
.Y(n_240)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_1),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_1),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_1),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_2),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_58),
.B1(n_93),
.B2(n_133),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_2),
.A2(n_93),
.B1(n_387),
.B2(n_389),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_2),
.A2(n_93),
.B1(n_252),
.B2(n_420),
.Y(n_419)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_3),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_3),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_3),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_4),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_5),
.A2(n_123),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_5),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_5),
.A2(n_182),
.B1(n_252),
.B2(n_255),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_5),
.A2(n_182),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_5),
.A2(n_61),
.B1(n_182),
.B2(n_415),
.Y(n_414)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_6),
.Y(n_336)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_8),
.A2(n_62),
.B1(n_227),
.B2(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_8),
.A2(n_62),
.B1(n_167),
.B2(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_8),
.A2(n_62),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_9),
.Y(n_176)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_11),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_11),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_12),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_12),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_12),
.A2(n_163),
.B1(n_195),
.B2(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_12),
.A2(n_163),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_12),
.A2(n_163),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_14),
.A2(n_160),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_14),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_14),
.A2(n_209),
.B1(n_224),
.B2(n_228),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_14),
.A2(n_46),
.B1(n_209),
.B2(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_14),
.A2(n_37),
.B1(n_53),
.B2(n_209),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_15),
.A2(n_54),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_15),
.A2(n_54),
.B1(n_395),
.B2(n_396),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_15),
.A2(n_54),
.B1(n_409),
.B2(n_410),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_16),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_16),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_16),
.A2(n_99),
.B1(n_105),
.B2(n_127),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_16),
.A2(n_37),
.B1(n_99),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_16),
.A2(n_99),
.B1(n_183),
.B2(n_391),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_17),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_17),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_17),
.A2(n_280),
.B1(n_374),
.B2(n_376),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_17),
.A2(n_280),
.B1(n_404),
.B2(n_407),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_L g459 ( 
.A1(n_17),
.A2(n_280),
.B1(n_333),
.B2(n_460),
.Y(n_459)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_535),
.B(n_538),
.Y(n_25)
);

AO21x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_140),
.B(n_534),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_137),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_28),
.B(n_137),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_131),
.C(n_134),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_29),
.A2(n_30),
.B1(n_530),
.B2(n_531),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_63),
.C(n_100),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_31),
.B(n_522),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_51),
.B1(n_55),
.B2(n_57),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_32),
.A2(n_55),
.B1(n_57),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_32),
.A2(n_55),
.B1(n_132),
.B2(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_32),
.A2(n_360),
.B(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_32),
.A2(n_55),
.B1(n_414),
.B2(n_434),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_32),
.A2(n_51),
.B1(n_55),
.B2(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_33),
.A2(n_340),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_33),
.B(n_361),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_33),
.A2(n_56),
.B(n_537),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_41),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_37),
.Y(n_362)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_46),
.B2(n_49),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_45),
.Y(n_264)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_45),
.Y(n_412)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_50),
.Y(n_338)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_52),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_55),
.B(n_157),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_55),
.A2(n_434),
.B(n_461),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_56),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_56),
.B(n_459),
.Y(n_458)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_58),
.Y(n_133)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_63),
.A2(n_100),
.B1(n_101),
.B2(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_63),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_89),
.B1(n_94),
.B2(n_95),
.Y(n_63)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_64),
.A2(n_94),
.B1(n_304),
.B2(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_64),
.A2(n_94),
.B1(n_403),
.B2(n_408),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_64),
.A2(n_89),
.B1(n_94),
.B2(n_511),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_79),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_74),
.B2(n_77),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_70),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_73),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_73),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_73),
.Y(n_332)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_73),
.Y(n_339)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_78),
.Y(n_306)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_78),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_79),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_79),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_79),
.A2(n_135),
.B1(n_308),
.B2(n_436),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_79),
.A2(n_135),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_82),
.Y(n_375)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_82),
.Y(n_395)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_83),
.Y(n_257)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_84),
.Y(n_400)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_87),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_91),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_92),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_94),
.B(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_94),
.A2(n_304),
.B(n_307),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_100),
.A2(n_101),
.B1(n_509),
.B2(n_510),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_100),
.B(n_506),
.C(n_509),
.Y(n_517)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_115),
.B(n_126),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_102),
.A2(n_150),
.B(n_158),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_102),
.A2(n_115),
.B1(n_207),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_102),
.A2(n_158),
.B(n_251),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_102),
.A2(n_115),
.B1(n_373),
.B2(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_103),
.B(n_159),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_103),
.A2(n_168),
.B1(n_394),
.B2(n_397),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_103),
.A2(n_168),
.B1(n_397),
.B2(n_419),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_103),
.A2(n_168),
.B1(n_419),
.B2(n_450),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_115),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_107),
.Y(n_254)
);

INVx6_ASAP7_75t_L g377 ( 
.A(n_107),
.Y(n_377)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_115),
.A2(n_207),
.B(n_210),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_115),
.A2(n_210),
.B(n_373),
.Y(n_372)
);

AOI22x1_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_121),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_123),
.B(n_217),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_124),
.Y(n_317)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_124),
.Y(n_388)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_126),
.Y(n_450)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_130),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_131),
.B(n_134),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_135),
.A2(n_260),
.B(n_268),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_135),
.B(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_135),
.A2(n_268),
.B(n_474),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_137),
.B(n_536),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_137),
.B(n_536),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_138),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_528),
.B(n_533),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_500),
.B(n_525),
.Y(n_141)
);

OAI311xp33_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_380),
.A3(n_476),
.B1(n_494),
.C1(n_499),
.Y(n_142)
);

AOI21x1_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_323),
.B(n_379),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_295),
.B(n_322),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_245),
.B(n_294),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_213),
.B(n_244),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_179),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_148),
.B(n_179),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_169),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_149),
.A2(n_169),
.B1(n_170),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_149),
.Y(n_242)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_157),
.A2(n_188),
.B(n_191),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_SL g260 ( 
.A1(n_157),
.A2(n_261),
.B(n_265),
.Y(n_260)
);

HAxp5_ASAP7_75t_SL g340 ( 
.A(n_157),
.B(n_341),
.CON(n_340),
.SN(n_340)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_168),
.Y(n_158)
);

INVx4_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_SL g421 ( 
.A(n_172),
.Y(n_421)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_204),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_180),
.B(n_205),
.C(n_212),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_188),
.B(n_191),
.Y(n_180)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_187),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_188),
.A2(n_346),
.B1(n_347),
.B2(n_350),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_188),
.A2(n_283),
.B1(n_386),
.B2(n_390),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_188),
.A2(n_231),
.B(n_390),
.Y(n_422)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_194),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_189),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_189),
.A2(n_278),
.B1(n_312),
.B2(n_318),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_189),
.A2(n_351),
.B1(n_429),
.B2(n_430),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_200),
.Y(n_313)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_202),
.Y(n_392)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx8_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_203),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_211),
.B2(n_212),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_235),
.B(n_243),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_221),
.B(n_234),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_219),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_233),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_233),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_231),
.B(n_232),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_229),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_232),
.A2(n_277),
.B(n_283),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_241),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_246),
.B(n_247),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_275),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_258),
.B2(n_259),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_258),
.C(n_275),
.Y(n_296)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_SL g292 ( 
.A(n_253),
.B(n_293),
.Y(n_292)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_254),
.Y(n_396)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_264),
.Y(n_409)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_264),
.Y(n_446)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI32xp33_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_286),
.A3(n_287),
.B1(n_290),
.B2(n_292),
.Y(n_285)
);

INVx8_ASAP7_75t_L g407 ( 
.A(n_267),
.Y(n_407)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx5_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_285),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_282),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_286),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_296),
.B(n_297),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_302),
.B2(n_321),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_301),
.C(n_321),
.Y(n_324)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_302),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_309),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_303),
.B(n_310),
.C(n_311),
.Y(n_353)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_312),
.Y(n_346)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx6_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_324),
.B(n_325),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_356),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_326)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_344),
.B2(n_345),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_329),
.B(n_344),
.Y(n_472)
);

OAI32xp33_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_333),
.A3(n_335),
.B1(n_337),
.B2(n_340),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_353),
.B(n_355),
.C(n_356),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_365),
.B2(n_378),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_357),
.B(n_366),
.C(n_372),
.Y(n_485)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_363),
.Y(n_460)
);

INVx8_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_365),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_372),
.Y(n_365)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_367),
.Y(n_474)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx8_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_462),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_SL g494 ( 
.A1(n_381),
.A2(n_462),
.B(n_495),
.C(n_498),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_437),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_382),
.B(n_437),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_416),
.C(n_424),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g475 ( 
.A(n_383),
.B(n_416),
.CI(n_424),
.CON(n_475),
.SN(n_475)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_401),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_384),
.B(n_402),
.C(n_413),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_393),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_385),
.B(n_393),
.Y(n_468)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_386),
.Y(n_429)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_394),
.Y(n_427)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_413),
.Y(n_401)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_403),
.Y(n_436)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx4_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_422),
.B2(n_423),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_422),
.Y(n_454)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_422),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_422),
.A2(n_423),
.B1(n_456),
.B2(n_457),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_422),
.A2(n_454),
.B(n_457),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_432),
.C(n_435),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_425),
.B(n_466),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_426),
.B(n_428),
.Y(n_484)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_432),
.A2(n_433),
.B1(n_435),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_435),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_438),
.B(n_441),
.C(n_452),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_452),
.B2(n_453),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_448),
.B(n_451),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_443),
.B(n_449),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_445),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

FAx1_ASAP7_75t_SL g502 ( 
.A(n_451),
.B(n_503),
.CI(n_504),
.CON(n_502),
.SN(n_502)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_451),
.B(n_503),
.C(n_504),
.Y(n_524)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_461),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_459),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_475),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_463),
.B(n_475),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_468),
.C(n_469),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_464),
.A2(n_465),
.B1(n_468),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_468),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_487),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_472),
.C(n_473),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_470),
.A2(n_471),
.B1(n_473),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_473),
.Y(n_482)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_475),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_489),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_478),
.A2(n_496),
.B(n_497),
.Y(n_495)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_486),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_486),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_483),
.C(n_485),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_492),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_483),
.A2(n_484),
.B1(n_485),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_485),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_491),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_514),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_513),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_502),
.B(n_513),
.Y(n_526)
);

BUFx24_ASAP7_75t_SL g542 ( 
.A(n_502),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_506),
.B1(n_508),
.B2(n_512),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_505),
.A2(n_506),
.B1(n_520),
.B2(n_521),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_516),
.C(n_520),
.Y(n_532)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_508),
.Y(n_512)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_514),
.A2(n_526),
.B(n_527),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_515),
.B(n_524),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_524),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_532),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_529),
.B(n_532),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_531),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g538 ( 
.A(n_539),
.Y(n_538)
);


endmodule