module fake_jpeg_4479_n_40 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_1),
.B(n_2),
.Y(n_19)
);

OAI22x1_ASAP7_75t_SL g24 ( 
.A1(n_19),
.A2(n_7),
.B1(n_8),
.B2(n_13),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_1),
.B(n_2),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_20),
.A2(n_9),
.B1(n_12),
.B2(n_4),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_12),
.B1(n_9),
.B2(n_13),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_18),
.C(n_19),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_26),
.C(n_24),
.Y(n_32)
);

OAI221xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_16),
.B1(n_7),
.B2(n_8),
.C(n_13),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_29),
.B(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_8),
.Y(n_31)
);

NOR3xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_35),
.C(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_29),
.B1(n_4),
.B2(n_3),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_25),
.C(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_37),
.B(n_38),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_25),
.Y(n_40)
);


endmodule