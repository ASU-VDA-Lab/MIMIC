module fake_jpeg_9882_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_219;
wire n_70;
wire n_121;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_23),
.C(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_32),
.B1(n_17),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_56),
.B1(n_31),
.B2(n_29),
.Y(n_88)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_61),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_17),
.B1(n_20),
.B2(n_25),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_57),
.A2(n_60),
.B1(n_64),
.B2(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_33),
.Y(n_86)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_21),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_35),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_17),
.B1(n_20),
.B2(n_25),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_35),
.A2(n_17),
.B1(n_20),
.B2(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_72),
.Y(n_95)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_73),
.B(n_84),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_1),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_43),
.B1(n_20),
.B2(n_29),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_93),
.B1(n_26),
.B2(n_19),
.Y(n_101)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_39),
.B1(n_55),
.B2(n_42),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_42),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_86),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_60),
.B1(n_51),
.B2(n_45),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_52),
.B1(n_49),
.B2(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_26),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_48),
.C(n_62),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_39),
.C(n_42),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_61),
.B(n_18),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_50),
.B(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_89),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_42),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_23),
.Y(n_92)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_43),
.B1(n_29),
.B2(n_18),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_98),
.A2(n_101),
.B1(n_104),
.B2(n_106),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_110),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_39),
.C(n_42),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_30),
.B1(n_24),
.B2(n_33),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_114),
.B1(n_91),
.B2(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_89),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_69),
.B1(n_87),
.B2(n_77),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_39),
.C(n_42),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_30),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_97),
.B1(n_100),
.B2(n_95),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_123),
.A2(n_128),
.B(n_129),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_124),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_126),
.A2(n_135),
.B1(n_138),
.B2(n_147),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_71),
.B1(n_91),
.B2(n_74),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_141),
.B(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_85),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_84),
.Y(n_132)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_72),
.B1(n_68),
.B2(n_88),
.Y(n_135)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_137),
.A2(n_144),
.B(n_113),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_74),
.B1(n_77),
.B2(n_70),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_103),
.B(n_86),
.Y(n_141)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_107),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_74),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_92),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_81),
.B1(n_87),
.B2(n_76),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_116),
.C(n_110),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_150),
.C(n_158),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_146),
.C(n_134),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_173),
.B1(n_135),
.B2(n_126),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_161),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_177),
.B(n_27),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_95),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_148),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_164),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_100),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_174),
.C(n_153),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_168),
.B(n_169),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_96),
.B(n_94),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_78),
.B(n_101),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_136),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_178),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_120),
.A2(n_104),
.B1(n_87),
.B2(n_78),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_93),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_1),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_144),
.B(n_139),
.Y(n_185)
);

AOI32xp33_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_39),
.A3(n_34),
.B1(n_27),
.B2(n_69),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_125),
.Y(n_178)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_182),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g182 ( 
.A(n_156),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_191),
.B1(n_199),
.B2(n_154),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_152),
.B(n_165),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_142),
.B(n_141),
.C(n_143),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_186),
.A2(n_27),
.B1(n_39),
.B2(n_21),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_1),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_188),
.A2(n_196),
.B(n_170),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_39),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_194),
.C(n_160),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_123),
.Y(n_193)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_1),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_2),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_202),
.Y(n_217)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_176),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_2),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_227),
.B1(n_200),
.B2(n_187),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_197),
.B(n_167),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_210),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_151),
.B1(n_172),
.B2(n_164),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_209),
.A2(n_193),
.B1(n_185),
.B2(n_188),
.Y(n_236)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_158),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_210),
.A2(n_220),
.B1(n_188),
.B2(n_189),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_168),
.B(n_163),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_215),
.C(n_184),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_160),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_219),
.B(n_226),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_196),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_121),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g225 ( 
.A(n_202),
.Y(n_225)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_234),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_183),
.B1(n_186),
.B2(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_231),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_213),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_184),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_243),
.B1(n_245),
.B2(n_211),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_217),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_242),
.Y(n_257)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_244),
.C(n_207),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_209),
.A2(n_196),
.B1(n_121),
.B2(n_190),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_241),
.B(n_206),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_21),
.C(n_4),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_238),
.C(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_208),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_258),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_256),
.B1(n_231),
.B2(n_227),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_230),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_216),
.C(n_211),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_234),
.C(n_244),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_216),
.B1(n_220),
.B2(n_225),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_235),
.B(n_218),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_205),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_259),
.B(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_260),
.Y(n_274)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_265),
.Y(n_276)
);

OAI221xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_229),
.B1(n_232),
.B2(n_240),
.C(n_10),
.Y(n_266)
);

OAI321xp33_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_6),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_240),
.C(n_7),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_269),
.B(n_21),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_6),
.C(n_7),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_271),
.Y(n_272)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_246),
.B1(n_252),
.B2(n_249),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_277),
.C(n_11),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_267),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_262),
.A2(n_254),
.B(n_248),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_16),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_268),
.A2(n_248),
.B(n_11),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_9),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_283),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_281),
.A2(n_270),
.B1(n_260),
.B2(n_12),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_9),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_285),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_14),
.C(n_15),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_13),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_287),
.Y(n_290)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_279),
.A3(n_272),
.B1(n_280),
.B2(n_274),
.C1(n_14),
.C2(n_15),
.Y(n_289)
);

OA21x2_ASAP7_75t_SL g295 ( 
.A1(n_289),
.A2(n_14),
.B(n_290),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_285),
.B(n_288),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_294),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_291),
.C(n_292),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_295),
.Y(n_298)
);


endmodule