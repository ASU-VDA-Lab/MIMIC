module fake_jpeg_20545_n_206 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_29),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_35),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_22),
.B1(n_20),
.B2(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_20),
.B1(n_12),
.B2(n_18),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_33),
.B1(n_26),
.B2(n_12),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_12),
.B1(n_18),
.B2(n_19),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_30),
.B1(n_31),
.B2(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_52),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_31),
.B1(n_25),
.B2(n_21),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_30),
.B(n_33),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_58),
.B(n_42),
.C(n_28),
.Y(n_73)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_43),
.B1(n_44),
.B2(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_16),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_15),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_37),
.Y(n_68)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_31),
.B1(n_42),
.B2(n_28),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_73),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_44),
.B1(n_41),
.B2(n_36),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_44),
.B1(n_41),
.B2(n_37),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_29),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_76),
.C(n_79),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_55),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_61),
.B1(n_57),
.B2(n_48),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_51),
.B1(n_55),
.B2(n_48),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_13),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_29),
.C(n_28),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_86),
.B1(n_77),
.B2(n_49),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_83),
.B(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_53),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_60),
.B(n_21),
.Y(n_117)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_47),
.B1(n_57),
.B2(n_49),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_71),
.B1(n_77),
.B2(n_59),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_62),
.B1(n_74),
.B2(n_72),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_110),
.B1(n_59),
.B2(n_42),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_102),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_74),
.B(n_66),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_107),
.B(n_13),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_96),
.B1(n_97),
.B2(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_95),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_16),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_19),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_113),
.B(n_111),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_80),
.C(n_85),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_122),
.C(n_137),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_129),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_120),
.A2(n_104),
.B1(n_124),
.B2(n_137),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_100),
.C(n_115),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_86),
.B1(n_82),
.B2(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_124),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_125),
.B(n_127),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_132),
.B1(n_105),
.B2(n_28),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_29),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_81),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_81),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_133),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_25),
.B1(n_21),
.B2(n_19),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_23),
.A3(n_27),
.B1(n_28),
.B2(n_25),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_23),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_98),
.C(n_113),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_17),
.B(n_23),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_142),
.B1(n_148),
.B2(n_0),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_104),
.B1(n_108),
.B2(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_27),
.C(n_17),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_126),
.C(n_122),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_132),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_27),
.A3(n_6),
.B1(n_7),
.B2(n_10),
.C1(n_9),
.C2(n_5),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_130),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_156),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_129),
.C(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_159),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_127),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_138),
.C(n_119),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_166),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_163),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_27),
.C(n_6),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_10),
.Y(n_166)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_141),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_145),
.C(n_27),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_153),
.B(n_144),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_139),
.B(n_142),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_139),
.C(n_153),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_182),
.C(n_183),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_144),
.B1(n_149),
.B2(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_171),
.A2(n_145),
.B(n_149),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_174),
.B(n_168),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_184),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_175),
.B(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_167),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_7),
.C(n_8),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_176),
.B(n_177),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_187),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_168),
.B(n_172),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_190),
.A2(n_169),
.B(n_1),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_2),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_169),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_197),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_198),
.C(n_3),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_0),
.B(n_2),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_3),
.B(n_4),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_3),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_196),
.A2(n_189),
.B(n_3),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_4),
.B(n_199),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_202),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_4),
.C(n_204),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_4),
.Y(n_206)
);


endmodule