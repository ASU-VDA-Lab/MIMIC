module fake_jpeg_2545_n_157 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_15),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_21),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_0),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_71),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_52),
.B1(n_54),
.B2(n_53),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_68),
.B1(n_60),
.B2(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_47),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_47),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_39),
.B1(n_51),
.B2(n_53),
.Y(n_68)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

OAI211xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_58),
.B(n_56),
.C(n_41),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_2),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_78),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_45),
.C(n_48),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_0),
.C(n_1),
.Y(n_96)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_84),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_70),
.B1(n_49),
.B2(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_4),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_59),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_38),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_90),
.B1(n_91),
.B2(n_97),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_71),
.B1(n_49),
.B2(n_46),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_46),
.B1(n_70),
.B2(n_40),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_40),
.B1(n_18),
.B2(n_24),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_25),
.B(n_33),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_101),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_7),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_108),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_85),
.B1(n_72),
.B2(n_79),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_105),
.B1(n_8),
.B2(n_9),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_99),
.B1(n_97),
.B2(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_5),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_5),
.B(n_6),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_116),
.B(n_13),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_115),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_7),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_34),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_11),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_125),
.B1(n_127),
.B2(n_132),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_32),
.B(n_30),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_128),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_130),
.B(n_107),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_27),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_116),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_14),
.B1(n_15),
.B2(n_28),
.Y(n_132)
);

INVxp33_ASAP7_75t_SL g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_135),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_136),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_125),
.A2(n_118),
.B1(n_129),
.B2(n_120),
.Y(n_139)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_141),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_138),
.B(n_128),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_147),
.A2(n_121),
.B(n_145),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_149),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_146),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_131),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_134),
.B(n_144),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_137),
.B(n_150),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_140),
.C(n_133),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_29),
.Y(n_157)
);


endmodule