module fake_jpeg_27368_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_6),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_17),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_31),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_16),
.A2(n_7),
.B(n_8),
.C(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

OA21x2_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_15),
.B(n_20),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_17),
.C(n_21),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_31),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_13),
.B1(n_20),
.B2(n_15),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_20),
.B1(n_13),
.B2(n_14),
.Y(n_50)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_56),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_51),
.B(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_14),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_13),
.B1(n_21),
.B2(n_19),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_63),
.B1(n_48),
.B2(n_25),
.Y(n_75)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_19),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_25),
.B1(n_18),
.B2(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_67),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_73),
.B(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_47),
.B1(n_45),
.B2(n_39),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_75),
.B1(n_45),
.B2(n_53),
.Y(n_88)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_39),
.B(n_42),
.C(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_79),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_58),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_39),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_24),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_12),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_52),
.B(n_57),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_88),
.B(n_79),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_52),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_86),
.C(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_90),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_99),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_70),
.B(n_71),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_69),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_75),
.B1(n_70),
.B2(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_103),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_68),
.C(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_88),
.Y(n_109)
);

OAI321xp33_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_69),
.A3(n_7),
.B1(n_2),
.B2(n_4),
.C(n_6),
.Y(n_102)
);

OA21x2_ASAP7_75t_SL g107 ( 
.A1(n_102),
.A2(n_82),
.B(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

XNOR2x1_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_96),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_92),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

AOI31xp67_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_97),
.A3(n_1),
.B(n_4),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_118),
.C(n_108),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_95),
.C(n_86),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_110),
.B(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_113),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_112),
.B1(n_105),
.B2(n_98),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_112),
.B(n_80),
.Y(n_122)
);

NAND4xp25_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_39),
.C(n_53),
.D(n_42),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_126),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_42),
.B1(n_4),
.B2(n_6),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_130),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_0),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_124),
.C(n_0),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

NAND2x1_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_128),
.Y(n_134)
);


endmodule