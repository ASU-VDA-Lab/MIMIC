module real_aes_11949_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1744;
wire n_1730;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1225;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_1712;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_1740;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1691;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1679;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_1735;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1647;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_394;
wire n_729;
wire n_1323;
wire n_1280;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g1269 ( .A1(n_0), .A2(n_719), .B1(n_734), .B2(n_1270), .C(n_1275), .Y(n_1269) );
AOI21xp33_ASAP7_75t_L g1302 ( .A1(n_0), .A2(n_567), .B(n_1303), .Y(n_1302) );
INVxp67_ASAP7_75t_L g811 ( .A(n_1), .Y(n_811) );
AOI221xp5_ASAP7_75t_L g852 ( .A1(n_1), .A2(n_189), .B1(n_838), .B2(n_853), .C(n_857), .Y(n_852) );
AOI221xp5_ASAP7_75t_L g558 ( .A1(n_2), .A2(n_61), .B1(n_559), .B2(n_561), .C(n_563), .Y(n_558) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_2), .A2(n_172), .B1(n_613), .B2(n_625), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g657 ( .A1(n_3), .A2(n_469), .B1(n_658), .B2(n_664), .C(n_670), .Y(n_657) );
INVx1_ASAP7_75t_L g688 ( .A(n_3), .Y(n_688) );
XNOR2x2_ASAP7_75t_L g1095 ( .A(n_4), .B(n_1096), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1228 ( .A1(n_5), .A2(n_72), .B1(n_1143), .B2(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1240 ( .A(n_5), .Y(n_1240) );
INVxp33_ASAP7_75t_L g1168 ( .A(n_6), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g1197 ( .A1(n_6), .A2(n_91), .B1(n_1198), .B2(n_1199), .C(n_1200), .Y(n_1197) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_7), .Y(n_1009) );
OAI221xp5_ASAP7_75t_L g786 ( .A1(n_8), .A2(n_242), .B1(n_787), .B2(n_788), .C(n_790), .Y(n_786) );
INVx1_ASAP7_75t_L g847 ( .A(n_8), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_9), .A2(n_103), .B1(n_606), .B2(n_649), .C(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g700 ( .A(n_9), .Y(n_700) );
INVx1_ASAP7_75t_L g1183 ( .A(n_10), .Y(n_1183) );
OAI221xp5_ASAP7_75t_L g1280 ( .A1(n_11), .A2(n_177), .B1(n_799), .B2(n_802), .C(n_804), .Y(n_1280) );
CKINVDCx5p33_ASAP7_75t_R g1308 ( .A(n_11), .Y(n_1308) );
AO22x1_ASAP7_75t_L g636 ( .A1(n_12), .A2(n_637), .B1(n_703), .B2(n_704), .Y(n_636) );
INVx1_ASAP7_75t_L g704 ( .A(n_12), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g1332 ( .A1(n_13), .A2(n_294), .B1(n_438), .B2(n_645), .C(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1340 ( .A(n_13), .Y(n_1340) );
INVx1_ASAP7_75t_L g896 ( .A(n_14), .Y(n_896) );
INVx1_ASAP7_75t_L g1444 ( .A(n_15), .Y(n_1444) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_16), .Y(n_826) );
INVx1_ASAP7_75t_L g1235 ( .A(n_17), .Y(n_1235) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_17), .A2(n_81), .B1(n_516), .B2(n_702), .Y(n_1258) );
INVx1_ASAP7_75t_L g1317 ( .A(n_18), .Y(n_1317) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_19), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_20), .A2(n_252), .B1(n_389), .B2(n_546), .Y(n_545) );
INVxp33_ASAP7_75t_SL g599 ( .A(n_20), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g1371 ( .A1(n_21), .A2(n_151), .B1(n_948), .B2(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1394 ( .A(n_21), .Y(n_1394) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_22), .A2(n_76), .B1(n_770), .B2(n_771), .C(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g777 ( .A(n_22), .Y(n_777) );
OAI221xp5_ASAP7_75t_L g796 ( .A1(n_23), .A2(n_111), .B1(n_797), .B2(n_800), .C(n_804), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_23), .A2(n_111), .B1(n_771), .B2(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g1223 ( .A(n_24), .Y(n_1223) );
OAI221xp5_ASAP7_75t_L g1243 ( .A1(n_24), .A2(n_469), .B1(n_488), .B2(n_1244), .C(n_1248), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_25), .A2(n_26), .B1(n_438), .B2(n_1101), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_25), .A2(n_266), .B1(n_512), .B2(n_516), .Y(n_1148) );
INVxp67_ASAP7_75t_SL g1146 ( .A(n_26), .Y(n_1146) );
AOI22xp5_ASAP7_75t_L g1415 ( .A1(n_27), .A2(n_125), .B1(n_1416), .B2(n_1424), .Y(n_1415) );
AOI221xp5_ASAP7_75t_L g1320 ( .A1(n_28), .A2(n_51), .B1(n_971), .B2(n_1321), .C(n_1322), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_28), .A2(n_270), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
CKINVDCx5p33_ASAP7_75t_R g1273 ( .A(n_29), .Y(n_1273) );
INVx1_ASAP7_75t_L g1324 ( .A(n_30), .Y(n_1324) );
AOI221xp5_ASAP7_75t_L g1342 ( .A1(n_30), .A2(n_51), .B1(n_1343), .B2(n_1344), .C(n_1346), .Y(n_1342) );
CKINVDCx5p33_ASAP7_75t_R g1734 ( .A(n_31), .Y(n_1734) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_32), .A2(n_89), .B1(n_855), .B2(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g975 ( .A(n_32), .Y(n_975) );
INVx1_ASAP7_75t_L g1121 ( .A(n_33), .Y(n_1121) );
AOI221xp5_ASAP7_75t_L g1127 ( .A1(n_33), .A2(n_169), .B1(n_561), .B2(n_1128), .C(n_1129), .Y(n_1127) );
OAI22xp5_ASAP7_75t_L g1282 ( .A1(n_34), .A2(n_73), .B1(n_1283), .B2(n_1284), .Y(n_1282) );
INVx1_ASAP7_75t_L g1300 ( .A(n_34), .Y(n_1300) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_35), .A2(n_57), .B1(n_928), .B2(n_946), .Y(n_945) );
AOI21xp33_ASAP7_75t_L g964 ( .A1(n_35), .A2(n_446), .B(n_720), .Y(n_964) );
INVxp33_ASAP7_75t_L g990 ( .A(n_36), .Y(n_990) );
AOI221xp5_ASAP7_75t_L g1014 ( .A1(n_36), .A2(n_88), .B1(n_371), .B2(n_944), .C(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1335 ( .A(n_37), .Y(n_1335) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_38), .A2(n_233), .B1(n_858), .B2(n_1022), .C(n_1025), .Y(n_1052) );
INVx1_ASAP7_75t_L g1081 ( .A(n_38), .Y(n_1081) );
AOI22xp33_ASAP7_75t_SL g997 ( .A1(n_39), .A2(n_162), .B1(n_998), .B2(n_999), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_39), .A2(n_162), .B1(n_1029), .B2(n_1031), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_40), .A2(n_48), .B1(n_645), .B2(n_646), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_40), .A2(n_103), .B1(n_516), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g1708 ( .A1(n_41), .A2(n_155), .B1(n_1343), .B2(n_1709), .Y(n_1708) );
AOI22xp33_ASAP7_75t_SL g1725 ( .A1(n_41), .A2(n_155), .B1(n_487), .B2(n_645), .Y(n_1725) );
INVx1_ASAP7_75t_L g318 ( .A(n_42), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g1434 ( .A1(n_43), .A2(n_119), .B1(n_1416), .B2(n_1424), .Y(n_1434) );
INVx1_ASAP7_75t_L g1156 ( .A(n_44), .Y(n_1156) );
INVx1_ASAP7_75t_L g383 ( .A(n_45), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_45), .A2(n_469), .B1(n_472), .B2(n_482), .C(n_488), .Y(n_468) );
INVx1_ASAP7_75t_L g1465 ( .A(n_46), .Y(n_1465) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_47), .Y(n_1203) );
INVx1_ASAP7_75t_L g696 ( .A(n_48), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_49), .A2(n_178), .B1(n_944), .B2(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1252 ( .A(n_49), .Y(n_1252) );
INVx1_ASAP7_75t_L g1125 ( .A(n_50), .Y(n_1125) );
INVx1_ASAP7_75t_L g436 ( .A(n_52), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_52), .A2(n_228), .B1(n_519), .B2(n_521), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_53), .A2(n_280), .B1(n_1002), .B2(n_1003), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1021 ( .A1(n_53), .A2(n_280), .B1(n_1022), .B2(n_1023), .C(n_1026), .Y(n_1021) );
INVx1_ASAP7_75t_L g1653 ( .A(n_54), .Y(n_1653) );
AOI22xp33_ASAP7_75t_L g1672 ( .A1(n_54), .A2(n_271), .B1(n_974), .B2(n_1673), .Y(n_1672) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_55), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_56), .A2(n_100), .B1(n_466), .B2(n_653), .Y(n_652) );
OAI22xp5_ASAP7_75t_SL g677 ( .A1(n_56), .A2(n_100), .B1(n_406), .B2(n_412), .Y(n_677) );
INVx1_ASAP7_75t_L g963 ( .A(n_57), .Y(n_963) );
INVx1_ASAP7_75t_L g924 ( .A(n_58), .Y(n_924) );
OAI221xp5_ASAP7_75t_L g932 ( .A1(n_58), .A2(n_268), .B1(n_933), .B2(n_934), .C(n_936), .Y(n_932) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_59), .A2(n_129), .B1(n_999), .B2(n_1002), .Y(n_1004) );
INVxp67_ASAP7_75t_SL g1012 ( .A(n_59), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_60), .A2(n_80), .B1(n_1428), .B2(n_1432), .Y(n_1427) );
AOI22xp33_ASAP7_75t_SL g618 ( .A1(n_61), .A2(n_156), .B1(n_619), .B2(n_621), .Y(n_618) );
INVxp33_ASAP7_75t_L g1155 ( .A(n_62), .Y(n_1155) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_62), .A2(n_115), .B1(n_1190), .B2(n_1192), .C(n_1193), .Y(n_1189) );
INVx1_ASAP7_75t_L g1316 ( .A(n_63), .Y(n_1316) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_64), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_65), .A2(n_170), .B1(n_446), .B2(n_450), .Y(n_1278) );
OAI22xp5_ASAP7_75t_L g1289 ( .A1(n_65), .A2(n_170), .B1(n_582), .B2(n_1290), .Y(n_1289) );
INVxp33_ASAP7_75t_L g1167 ( .A(n_66), .Y(n_1167) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_66), .A2(n_265), .B1(n_540), .B2(n_749), .Y(n_1201) );
OAI221xp5_ASAP7_75t_L g1161 ( .A1(n_67), .A2(n_224), .B1(n_878), .B2(n_1071), .C(n_1162), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_67), .A2(n_224), .B1(n_552), .B2(n_771), .Y(n_1188) );
OAI221xp5_ASAP7_75t_L g1112 ( .A1(n_68), .A2(n_469), .B1(n_488), .B2(n_1113), .C(n_1119), .Y(n_1112) );
AOI221xp5_ASAP7_75t_L g1132 ( .A1(n_68), .A2(n_229), .B1(n_860), .B2(n_1133), .C(n_1135), .Y(n_1132) );
INVx1_ASAP7_75t_L g675 ( .A(n_69), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g1451 ( .A1(n_70), .A2(n_197), .B1(n_1416), .B2(n_1424), .Y(n_1451) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_71), .Y(n_550) );
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_71), .A2(n_193), .B1(n_613), .B2(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g1242 ( .A(n_72), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_73), .A2(n_117), .B1(n_369), .B2(n_1298), .Y(n_1301) );
AO22x1_ASAP7_75t_SL g1490 ( .A1(n_74), .A2(n_126), .B1(n_1416), .B2(n_1424), .Y(n_1490) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_75), .A2(n_285), .B1(n_530), .B2(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g774 ( .A(n_75), .Y(n_774) );
INVx1_ASAP7_75t_L g778 ( .A(n_76), .Y(n_778) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_77), .A2(n_112), .B1(n_998), .B2(n_1003), .Y(n_1005) );
INVxp67_ASAP7_75t_L g1020 ( .A(n_77), .Y(n_1020) );
CKINVDCx5p33_ASAP7_75t_R g1047 ( .A(n_78), .Y(n_1047) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_79), .Y(n_824) );
AOI221xp5_ASAP7_75t_L g1236 ( .A1(n_81), .A2(n_305), .B1(n_649), .B2(n_1237), .C(n_1238), .Y(n_1236) );
AOI22xp5_ASAP7_75t_L g1452 ( .A1(n_82), .A2(n_216), .B1(n_1432), .B2(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1226 ( .A(n_83), .Y(n_1226) );
OAI211xp5_ASAP7_75t_L g1231 ( .A1(n_83), .A2(n_419), .B(n_1232), .C(n_1239), .Y(n_1231) );
OAI222xp33_ASAP7_75t_L g876 ( .A1(n_84), .A2(n_140), .B1(n_278), .B2(n_530), .C1(n_877), .C2(n_878), .Y(n_876) );
INVx1_ASAP7_75t_L g909 ( .A(n_84), .Y(n_909) );
OAI211xp5_ASAP7_75t_SL g1660 ( .A1(n_85), .A2(n_1288), .B(n_1661), .C(n_1664), .Y(n_1660) );
AOI22xp33_ASAP7_75t_L g1678 ( .A1(n_85), .A2(n_185), .B1(n_1675), .B2(n_1679), .Y(n_1678) );
AOI22xp33_ASAP7_75t_L g1227 ( .A1(n_86), .A2(n_218), .B1(n_839), .B2(n_950), .Y(n_1227) );
OAI22xp5_ASAP7_75t_L g1253 ( .A1(n_86), .A2(n_218), .B1(n_1254), .B2(n_1255), .Y(n_1253) );
AO22x2_ASAP7_75t_L g705 ( .A1(n_87), .A2(n_706), .B1(n_779), .B2(n_780), .Y(n_705) );
CKINVDCx14_ASAP7_75t_R g779 ( .A(n_87), .Y(n_779) );
INVxp33_ASAP7_75t_SL g994 ( .A(n_88), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_89), .A2(n_94), .B1(n_422), .B2(n_461), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g1456 ( .A1(n_90), .A2(n_110), .B1(n_1432), .B2(n_1453), .Y(n_1456) );
INVxp67_ASAP7_75t_L g1171 ( .A(n_91), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_92), .A2(n_106), .B1(n_749), .B2(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g968 ( .A(n_92), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g1379 ( .A1(n_93), .A2(n_304), .B1(n_1050), .B2(n_1380), .Y(n_1379) );
OAI221xp5_ASAP7_75t_L g1391 ( .A1(n_93), .A2(n_304), .B1(n_797), .B2(n_801), .C(n_1071), .Y(n_1391) );
OAI222xp33_ASAP7_75t_L g980 ( .A1(n_94), .A2(n_134), .B1(n_217), .B2(n_519), .C1(n_521), .C2(n_532), .Y(n_980) );
BUFx2_ASAP7_75t_L g350 ( .A(n_95), .Y(n_350) );
BUFx2_ASAP7_75t_L g377 ( .A(n_95), .Y(n_377) );
INVx1_ASAP7_75t_L g403 ( .A(n_95), .Y(n_403) );
OR2x2_ASAP7_75t_L g531 ( .A(n_95), .B(n_463), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g1274 ( .A1(n_96), .A2(n_138), .B1(n_446), .B2(n_450), .Y(n_1274) );
INVx1_ASAP7_75t_L g1296 ( .A(n_96), .Y(n_1296) );
INVx1_ASAP7_75t_L g365 ( .A(n_97), .Y(n_365) );
INVx1_ASAP7_75t_L g1467 ( .A(n_98), .Y(n_1467) );
INVx1_ASAP7_75t_L g663 ( .A(n_99), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_99), .A2(n_214), .B1(n_390), .B2(n_560), .Y(n_684) );
INVx1_ASAP7_75t_L g956 ( .A(n_101), .Y(n_956) );
OAI221xp5_ASAP7_75t_L g976 ( .A1(n_101), .A2(n_195), .B1(n_466), .B2(n_653), .C(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_102), .A2(n_274), .B1(n_1416), .B2(n_1424), .Y(n_1477) );
INVx1_ASAP7_75t_L g642 ( .A(n_104), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_104), .A2(n_251), .B1(n_388), .B2(n_390), .Y(n_690) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_105), .Y(n_503) );
INVx1_ASAP7_75t_L g966 ( .A(n_106), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g1435 ( .A1(n_107), .A2(n_248), .B1(n_1428), .B2(n_1432), .Y(n_1435) );
AO221x1_ASAP7_75t_L g1729 ( .A1(n_108), .A2(n_191), .B1(n_450), .B2(n_451), .C(n_979), .Y(n_1729) );
INVx1_ASAP7_75t_L g1739 ( .A(n_108), .Y(n_1739) );
AOI221xp5_ASAP7_75t_L g1370 ( .A1(n_109), .A2(n_188), .B1(n_915), .B2(n_916), .C(n_1025), .Y(n_1370) );
INVxp67_ASAP7_75t_SL g1398 ( .A(n_109), .Y(n_1398) );
INVxp33_ASAP7_75t_L g1033 ( .A(n_112), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1644 ( .A1(n_113), .A2(n_1645), .B1(n_1646), .B2(n_1647), .Y(n_1644) );
CKINVDCx5p33_ASAP7_75t_R g1645 ( .A(n_113), .Y(n_1645) );
INVx1_ASAP7_75t_L g1334 ( .A(n_114), .Y(n_1334) );
OAI221xp5_ASAP7_75t_L g1338 ( .A1(n_114), .A2(n_294), .B1(n_353), .B2(n_1130), .C(n_1339), .Y(n_1338) );
INVxp33_ASAP7_75t_L g1159 ( .A(n_115), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_116), .A2(n_131), .B1(n_387), .B2(n_389), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_116), .A2(n_131), .B1(n_491), .B2(n_496), .Y(n_490) );
OAI22xp33_ASAP7_75t_L g1285 ( .A1(n_117), .A2(n_136), .B1(n_530), .B2(n_743), .Y(n_1285) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_118), .A2(n_163), .B1(n_552), .B2(n_555), .Y(n_551) );
INVxp67_ASAP7_75t_SL g591 ( .A(n_118), .Y(n_591) );
INVx1_ASAP7_75t_L g1493 ( .A(n_120), .Y(n_1493) );
INVx1_ASAP7_75t_L g993 ( .A(n_121), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1710 ( .A1(n_122), .A2(n_259), .B1(n_751), .B2(n_1348), .Y(n_1710) );
AOI221xp5_ASAP7_75t_L g1726 ( .A1(n_122), .A2(n_259), .B1(n_606), .B2(n_649), .C(n_720), .Y(n_1726) );
INVx1_ASAP7_75t_L g791 ( .A(n_123), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g1375 ( .A1(n_124), .A2(n_154), .B1(n_698), .B2(n_764), .C(n_1025), .Y(n_1375) );
INVx1_ASAP7_75t_L g1389 ( .A(n_124), .Y(n_1389) );
INVx1_ASAP7_75t_L g1206 ( .A(n_125), .Y(n_1206) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_127), .Y(n_1058) );
XOR2x2_ASAP7_75t_L g340 ( .A(n_128), .B(n_341), .Y(n_340) );
INVxp33_ASAP7_75t_L g1034 ( .A(n_129), .Y(n_1034) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_130), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_132), .Y(n_1057) );
CKINVDCx5p33_ASAP7_75t_R g1663 ( .A(n_133), .Y(n_1663) );
AOI221xp5_ASAP7_75t_L g972 ( .A1(n_134), .A2(n_256), .B1(n_650), .B2(n_973), .C(n_974), .Y(n_972) );
INVxp67_ASAP7_75t_SL g987 ( .A(n_135), .Y(n_987) );
OAI22xp33_ASAP7_75t_L g1013 ( .A1(n_135), .A2(n_166), .B1(n_771), .B2(n_836), .Y(n_1013) );
INVx1_ASAP7_75t_L g1305 ( .A(n_136), .Y(n_1305) );
INVx1_ASAP7_75t_L g1369 ( .A(n_137), .Y(n_1369) );
INVx1_ASAP7_75t_L g1293 ( .A(n_138), .Y(n_1293) );
AOI21xp33_ASAP7_75t_L g1658 ( .A1(n_139), .A2(n_560), .B(n_858), .Y(n_1658) );
AOI22xp33_ASAP7_75t_L g1674 ( .A1(n_139), .A2(n_165), .B1(n_1675), .B2(n_1677), .Y(n_1674) );
INVx1_ASAP7_75t_L g921 ( .A(n_140), .Y(n_921) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_141), .Y(n_725) );
INVx1_ASAP7_75t_L g443 ( .A(n_142), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_142), .A2(n_209), .B1(n_512), .B2(n_516), .Y(n_511) );
OAI22xp33_ASAP7_75t_L g1668 ( .A1(n_143), .A2(n_185), .B1(n_582), .B2(n_585), .Y(n_1668) );
AOI22xp33_ASAP7_75t_L g1680 ( .A1(n_143), .A2(n_254), .B1(n_974), .B2(n_1681), .Y(n_1680) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_144), .Y(n_1054) );
CKINVDCx5p33_ASAP7_75t_R g1662 ( .A(n_145), .Y(n_1662) );
INVx1_ASAP7_75t_L g1116 ( .A(n_146), .Y(n_1116) );
INVx1_ASAP7_75t_L g1420 ( .A(n_147), .Y(n_1420) );
AOI221xp5_ASAP7_75t_L g1103 ( .A1(n_148), .A2(n_266), .B1(n_650), .B2(n_1104), .C(n_1106), .Y(n_1103) );
INVxp67_ASAP7_75t_SL g1147 ( .A(n_148), .Y(n_1147) );
INVx1_ASAP7_75t_L g714 ( .A(n_149), .Y(n_714) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_149), .A2(n_282), .B1(n_390), .B2(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g1158 ( .A(n_150), .Y(n_1158) );
INVx1_ASAP7_75t_L g1399 ( .A(n_151), .Y(n_1399) );
OAI22xp5_ASAP7_75t_L g1360 ( .A1(n_152), .A2(n_1361), .B1(n_1403), .B2(n_1404), .Y(n_1360) );
INVx1_ASAP7_75t_L g1404 ( .A(n_152), .Y(n_1404) );
AOI221xp5_ASAP7_75t_L g1461 ( .A1(n_153), .A2(n_232), .B1(n_1462), .B2(n_1463), .C(n_1464), .Y(n_1461) );
INVx1_ASAP7_75t_L g1387 ( .A(n_154), .Y(n_1387) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_156), .A2(n_172), .B1(n_565), .B2(n_568), .Y(n_564) );
INVx1_ASAP7_75t_L g360 ( .A(n_157), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_158), .A2(n_201), .B1(n_1377), .B2(n_1378), .Y(n_1376) );
INVx1_ASAP7_75t_L g1386 ( .A(n_158), .Y(n_1386) );
INVx1_ASAP7_75t_L g1421 ( .A(n_159), .Y(n_1421) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_159), .B(n_1419), .Y(n_1426) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_160), .A2(n_190), .B1(n_368), .B2(n_389), .Y(n_1045) );
INVx1_ASAP7_75t_L g1063 ( .A(n_160), .Y(n_1063) );
INVx1_ASAP7_75t_L g886 ( .A(n_161), .Y(n_886) );
INVxp67_ASAP7_75t_SL g595 ( .A(n_163), .Y(n_595) );
INVx2_ASAP7_75t_L g330 ( .A(n_164), .Y(n_330) );
INVx1_ASAP7_75t_L g1655 ( .A(n_165), .Y(n_1655) );
INVxp67_ASAP7_75t_SL g988 ( .A(n_166), .Y(n_988) );
INVxp67_ASAP7_75t_L g888 ( .A(n_167), .Y(n_888) );
OAI222xp33_ASAP7_75t_L g911 ( .A1(n_167), .A2(n_175), .B1(n_263), .B2(n_353), .C1(n_522), .C2(n_912), .Y(n_911) );
AO221x2_ASAP7_75t_L g1438 ( .A1(n_168), .A2(n_206), .B1(n_1428), .B2(n_1439), .C(n_1441), .Y(n_1438) );
AOI21xp33_ASAP7_75t_L g1122 ( .A1(n_169), .A2(n_720), .B(n_1104), .Y(n_1122) );
INVx1_ASAP7_75t_L g357 ( .A(n_171), .Y(n_357) );
BUFx3_ASAP7_75t_L g370 ( .A(n_171), .Y(n_370) );
XNOR2x2_ASAP7_75t_L g783 ( .A(n_173), .B(n_784), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g1732 ( .A(n_174), .Y(n_1732) );
INVxp67_ASAP7_75t_L g894 ( .A(n_175), .Y(n_894) );
INVxp67_ASAP7_75t_L g819 ( .A(n_176), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_176), .A2(n_246), .B1(n_860), .B2(n_861), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g1309 ( .A(n_177), .Y(n_1309) );
INVx1_ASAP7_75t_L g1249 ( .A(n_178), .Y(n_1249) );
INVx1_ASAP7_75t_L g709 ( .A(n_179), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g768 ( .A1(n_179), .A2(n_388), .B(n_563), .Y(n_768) );
INVx1_ASAP7_75t_L g1177 ( .A(n_180), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g1718 ( .A(n_181), .Y(n_1718) );
INVx1_ASAP7_75t_L g1325 ( .A(n_182), .Y(n_1325) );
INVx1_ASAP7_75t_L g1181 ( .A(n_183), .Y(n_1181) );
AOI22xp33_ASAP7_75t_SL g1715 ( .A1(n_184), .A2(n_311), .B1(n_693), .B2(n_1372), .Y(n_1715) );
INVx1_ASAP7_75t_L g1722 ( .A(n_184), .Y(n_1722) );
INVx1_ASAP7_75t_L g1118 ( .A(n_186), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_187), .A2(n_296), .B1(n_367), .B2(n_371), .Y(n_366) );
INVxp67_ASAP7_75t_SL g485 ( .A(n_187), .Y(n_485) );
INVxp67_ASAP7_75t_SL g1395 ( .A(n_188), .Y(n_1395) );
INVxp67_ASAP7_75t_L g815 ( .A(n_189), .Y(n_815) );
INVx1_ASAP7_75t_L g1067 ( .A(n_190), .Y(n_1067) );
INVx1_ASAP7_75t_L g1742 ( .A(n_191), .Y(n_1742) );
INVx1_ASAP7_75t_L g347 ( .A(n_192), .Y(n_347) );
INVx1_ASAP7_75t_L g401 ( .A(n_192), .Y(n_401) );
INVxp33_ASAP7_75t_L g583 ( .A(n_193), .Y(n_583) );
INVx1_ASAP7_75t_L g1366 ( .A(n_194), .Y(n_1366) );
INVx1_ASAP7_75t_L g954 ( .A(n_195), .Y(n_954) );
INVx1_ASAP7_75t_L g991 ( .A(n_196), .Y(n_991) );
XNOR2xp5_ASAP7_75t_L g873 ( .A(n_197), .B(n_874), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g1056 ( .A(n_198), .Y(n_1056) );
INVxp67_ASAP7_75t_L g881 ( .A(n_199), .Y(n_881) );
AOI221xp5_ASAP7_75t_L g914 ( .A1(n_199), .A2(n_286), .B1(n_751), .B2(n_915), .C(n_916), .Y(n_914) );
OAI21xp33_ASAP7_75t_L g1313 ( .A1(n_200), .A2(n_1314), .B(n_1336), .Y(n_1313) );
INVx1_ASAP7_75t_L g1357 ( .A(n_200), .Y(n_1357) );
INVx1_ASAP7_75t_L g1390 ( .A(n_201), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1711 ( .A1(n_202), .A2(n_292), .B1(n_1025), .B2(n_1712), .Y(n_1711) );
OAI221xp5_ASAP7_75t_L g1728 ( .A1(n_202), .A2(n_419), .B1(n_1729), .B2(n_1730), .C(n_1733), .Y(n_1728) );
INVxp67_ASAP7_75t_SL g575 ( .A(n_203), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g629 ( .A1(n_203), .A2(n_267), .B1(n_621), .B2(n_630), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g724 ( .A(n_204), .Y(n_724) );
OA22x2_ASAP7_75t_L g1039 ( .A1(n_205), .A2(n_1040), .B1(n_1091), .B2(n_1092), .Y(n_1039) );
INVx1_ASAP7_75t_L g1092 ( .A(n_205), .Y(n_1092) );
XOR2xp5_ASAP7_75t_L g1266 ( .A(n_207), .B(n_1267), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1455 ( .A1(n_207), .A2(n_258), .B1(n_1416), .B2(n_1424), .Y(n_1455) );
INVx1_ASAP7_75t_L g1150 ( .A(n_208), .Y(n_1150) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_209), .A2(n_228), .B1(n_445), .B2(n_449), .C(n_451), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g1478 ( .A1(n_210), .A2(n_273), .B1(n_1432), .B2(n_1453), .Y(n_1478) );
XNOR2xp5_ASAP7_75t_L g938 ( .A(n_211), .B(n_939), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g1666 ( .A1(n_212), .A2(n_260), .B1(n_388), .B2(n_390), .Y(n_1666) );
OAI22xp5_ASAP7_75t_L g1686 ( .A1(n_212), .A2(n_307), .B1(n_743), .B2(n_1284), .Y(n_1686) );
INVx1_ASAP7_75t_L g1331 ( .A(n_213), .Y(n_1331) );
AOI221xp5_ASAP7_75t_L g1351 ( .A1(n_213), .A2(n_272), .B1(n_748), .B2(n_1303), .C(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g661 ( .A(n_214), .Y(n_661) );
INVx1_ASAP7_75t_L g1234 ( .A(n_215), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_215), .A2(n_305), .B1(n_519), .B2(n_521), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_217), .A2(n_300), .B1(n_646), .B2(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g1184 ( .A(n_219), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_220), .A2(n_227), .B1(n_738), .B2(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g757 ( .A(n_220), .Y(n_757) );
OA332x1_ASAP7_75t_L g707 ( .A1(n_221), .A2(n_708), .A3(n_713), .B1(n_719), .B2(n_722), .B3(n_726), .C1(n_733), .C2(n_734), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_221), .A2(n_763), .B(n_764), .Y(n_762) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_222), .A2(n_237), .B1(n_537), .B2(n_540), .C(n_543), .Y(n_536) );
INVxp33_ASAP7_75t_SL g604 ( .A(n_222), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_223), .A2(n_283), .B1(n_466), .B2(n_653), .Y(n_1108) );
OAI221xp5_ASAP7_75t_L g1140 ( .A1(n_223), .A2(n_283), .B1(n_1141), .B2(n_1143), .C(n_1144), .Y(n_1140) );
INVx1_ASAP7_75t_L g1382 ( .A(n_225), .Y(n_1382) );
INVx1_ASAP7_75t_L g1494 ( .A(n_226), .Y(n_1494) );
AOI22xp33_ASAP7_75t_SL g761 ( .A1(n_227), .A2(n_285), .B1(n_388), .B2(n_390), .Y(n_761) );
OAI211xp5_ASAP7_75t_L g1098 ( .A1(n_229), .A2(n_419), .B(n_1099), .C(n_1109), .Y(n_1098) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_230), .Y(n_525) );
INVx1_ASAP7_75t_L g1110 ( .A(n_231), .Y(n_1110) );
INVx1_ASAP7_75t_L g1078 ( .A(n_233), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_234), .A2(n_236), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
OAI221xp5_ASAP7_75t_L g1069 ( .A1(n_234), .A2(n_236), .B1(n_801), .B2(n_1070), .C(n_1071), .Y(n_1069) );
INVx1_ASAP7_75t_L g907 ( .A(n_235), .Y(n_907) );
INVxp33_ASAP7_75t_L g608 ( .A(n_237), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_238), .Y(n_669) );
INVx1_ASAP7_75t_L g385 ( .A(n_239), .Y(n_385) );
OAI211xp5_ASAP7_75t_SL g418 ( .A1(n_239), .A2(n_419), .B(n_429), .C(n_455), .Y(n_418) );
INVx1_ASAP7_75t_L g1111 ( .A(n_240), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1044 ( .A1(n_241), .A2(n_253), .B1(n_928), .B2(n_929), .C(n_1025), .Y(n_1044) );
INVx1_ASAP7_75t_L g1064 ( .A(n_241), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_242), .A2(n_309), .B1(n_838), .B2(n_841), .C(n_844), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g1035 ( .A(n_243), .Y(n_1035) );
INVx1_ASAP7_75t_L g359 ( .A(n_244), .Y(n_359) );
BUFx3_ASAP7_75t_L g374 ( .A(n_244), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g1717 ( .A(n_245), .Y(n_1717) );
INVxp67_ASAP7_75t_L g808 ( .A(n_246), .Y(n_808) );
AOI21xp33_ASAP7_75t_L g1667 ( .A1(n_247), .A2(n_698), .B(n_764), .Y(n_1667) );
INVx1_ASAP7_75t_L g1684 ( .A(n_247), .Y(n_1684) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_249), .Y(n_326) );
AND2x2_ASAP7_75t_L g423 ( .A(n_249), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g454 ( .A(n_249), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_249), .B(n_297), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g1731 ( .A(n_250), .Y(n_1731) );
INVx1_ASAP7_75t_L g641 ( .A(n_251), .Y(n_641) );
INVxp33_ASAP7_75t_SL g611 ( .A(n_252), .Y(n_611) );
INVx1_ASAP7_75t_L g1066 ( .A(n_253), .Y(n_1066) );
OAI221xp5_ASAP7_75t_L g1651 ( .A1(n_254), .A2(n_1290), .B1(n_1652), .B2(n_1656), .C(n_1659), .Y(n_1651) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_255), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_256), .A2(n_300), .B1(n_512), .B2(n_516), .Y(n_981) );
INVx2_ASAP7_75t_L g348 ( .A(n_257), .Y(n_348) );
OR2x2_ASAP7_75t_L g515 ( .A(n_257), .B(n_401), .Y(n_515) );
INVx1_ASAP7_75t_L g1685 ( .A(n_260), .Y(n_1685) );
INVx1_ASAP7_75t_L g883 ( .A(n_261), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_262), .A2(n_269), .B1(n_493), .B2(n_1277), .Y(n_1276) );
OAI22xp5_ASAP7_75t_L g1287 ( .A1(n_262), .A2(n_269), .B1(n_585), .B2(n_1288), .Y(n_1287) );
INVxp67_ASAP7_75t_L g892 ( .A(n_263), .Y(n_892) );
INVx1_ASAP7_75t_L g1271 ( .A(n_264), .Y(n_1271) );
AOI21xp33_ASAP7_75t_L g1294 ( .A1(n_264), .A2(n_858), .B(n_915), .Y(n_1294) );
INVxp67_ASAP7_75t_L g1173 ( .A(n_265), .Y(n_1173) );
INVxp33_ASAP7_75t_SL g580 ( .A(n_267), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g925 ( .A1(n_268), .A2(n_281), .B1(n_926), .B2(n_928), .C(n_929), .Y(n_925) );
INVxp67_ASAP7_75t_SL g1323 ( .A(n_270), .Y(n_1323) );
INVx1_ASAP7_75t_L g1657 ( .A(n_271), .Y(n_1657) );
INVx1_ASAP7_75t_L g1330 ( .A(n_272), .Y(n_1330) );
AOI22xp5_ASAP7_75t_L g1692 ( .A1(n_273), .A2(n_1693), .B1(n_1698), .B2(n_1745), .Y(n_1692) );
AOI22x1_ASAP7_75t_L g1701 ( .A1(n_273), .A2(n_1702), .B1(n_1703), .B2(n_1744), .Y(n_1701) );
INVxp67_ASAP7_75t_SL g1744 ( .A(n_273), .Y(n_1744) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_275), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_276), .A2(n_303), .B1(n_405), .B2(n_412), .Y(n_404) );
INVx1_ASAP7_75t_L g464 ( .A(n_276), .Y(n_464) );
OAI221xp5_ASAP7_75t_SL g1328 ( .A1(n_277), .A2(n_301), .B1(n_432), .B2(n_1117), .C(n_1329), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g1353 ( .A1(n_277), .A2(n_301), .B1(n_560), .B2(n_570), .Y(n_1353) );
INVx1_ASAP7_75t_L g903 ( .A(n_278), .Y(n_903) );
CKINVDCx5p33_ASAP7_75t_R g731 ( .A(n_279), .Y(n_731) );
OAI332xp33_ASAP7_75t_L g879 ( .A1(n_281), .A2(n_719), .A3(n_740), .B1(n_880), .B2(n_884), .B3(n_887), .C1(n_893), .C2(n_897), .Y(n_879) );
INVx1_ASAP7_75t_L g710 ( .A(n_282), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g949 ( .A1(n_284), .A2(n_287), .B1(n_840), .B2(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g959 ( .A(n_284), .Y(n_959) );
INVx1_ASAP7_75t_L g885 ( .A(n_286), .Y(n_885) );
INVx1_ASAP7_75t_L g960 ( .A(n_287), .Y(n_960) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_288), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_288), .B(n_318), .Y(n_1423) );
AND3x2_ASAP7_75t_L g1431 ( .A(n_288), .B(n_318), .C(n_1420), .Y(n_1431) );
CKINVDCx5p33_ASAP7_75t_R g1209 ( .A(n_289), .Y(n_1209) );
INVx2_ASAP7_75t_L g331 ( .A(n_290), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_291), .A2(n_306), .B1(n_841), .B2(n_928), .Y(n_1053) );
INVx1_ASAP7_75t_L g1077 ( .A(n_291), .Y(n_1077) );
INVx1_ASAP7_75t_L g1727 ( .A(n_292), .Y(n_1727) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_293), .A2(n_419), .B(n_640), .C(n_643), .Y(n_639) );
INVx1_ASAP7_75t_L g689 ( .A(n_293), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g1218 ( .A(n_295), .Y(n_1218) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_296), .Y(n_483) );
INVx1_ASAP7_75t_L g333 ( .A(n_297), .Y(n_333) );
INVx2_ASAP7_75t_L g424 ( .A(n_297), .Y(n_424) );
OR2x2_ASAP7_75t_L g1649 ( .A(n_298), .B(n_529), .Y(n_1649) );
CKINVDCx5p33_ASAP7_75t_R g1214 ( .A(n_299), .Y(n_1214) );
INVx1_ASAP7_75t_L g1374 ( .A(n_302), .Y(n_1374) );
INVx1_ASAP7_75t_L g456 ( .A(n_303), .Y(n_456) );
INVx1_ASAP7_75t_L g1083 ( .A(n_306), .Y(n_1083) );
INVx1_ASAP7_75t_L g1665 ( .A(n_307), .Y(n_1665) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_308), .Y(n_715) );
INVxp33_ASAP7_75t_SL g793 ( .A(n_309), .Y(n_793) );
INVx1_ASAP7_75t_L g1365 ( .A(n_310), .Y(n_1365) );
INVx1_ASAP7_75t_L g1723 ( .A(n_311), .Y(n_1723) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_334), .B(n_1405), .Y(n_312) );
BUFx12f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_321), .Y(n_315) );
AND2x4_ASAP7_75t_L g1697 ( .A(n_316), .B(n_322), .Y(n_1697) );
NOR2xp33_ASAP7_75t_SL g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_SL g1691 ( .A(n_317), .Y(n_1691) );
NAND2xp5_ASAP7_75t_L g1750 ( .A(n_317), .B(n_319), .Y(n_1750) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_319), .B(n_1691), .Y(n_1690) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_327), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g481 ( .A(n_325), .B(n_333), .Y(n_481) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OR2x2_ASAP7_75t_L g720 ( .A(n_326), .B(n_721), .Y(n_720) );
OR2x6_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
INVx2_ASAP7_75t_SL g479 ( .A(n_328), .Y(n_479) );
OR2x2_ASAP7_75t_L g530 ( .A(n_328), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_SL g668 ( .A(n_328), .Y(n_668) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_328), .Y(n_723) );
INVx1_ASAP7_75t_L g810 ( .A(n_328), .Y(n_810) );
BUFx2_ASAP7_75t_L g1076 ( .A(n_328), .Y(n_1076) );
OAI22xp33_ASAP7_75t_L g1322 ( .A1(n_328), .A2(n_717), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
OAI22xp33_ASAP7_75t_L g1333 ( .A1(n_328), .A2(n_717), .B1(n_1334), .B2(n_1335), .Y(n_1333) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g427 ( .A(n_330), .Y(n_427) );
INVx2_ASAP7_75t_L g435 ( .A(n_330), .Y(n_435) );
AND2x4_ASAP7_75t_L g442 ( .A(n_330), .B(n_428), .Y(n_442) );
AND2x2_ASAP7_75t_L g448 ( .A(n_330), .B(n_331), .Y(n_448) );
INVx1_ASAP7_75t_L g477 ( .A(n_330), .Y(n_477) );
INVx2_ASAP7_75t_L g428 ( .A(n_331), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_331), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g459 ( .A(n_331), .Y(n_459) );
INVx1_ASAP7_75t_L g476 ( .A(n_331), .Y(n_476) );
INVx1_ASAP7_75t_L g495 ( .A(n_331), .Y(n_495) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_1262), .B2(n_1263), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
XNOR2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_781), .Y(n_336) );
XOR2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_634), .Y(n_337) );
AO22x1_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_523), .B2(n_633), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND4x1_ASAP7_75t_L g341 ( .A(n_342), .B(n_417), .C(n_502), .D(n_510), .Y(n_341) );
NOR3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_391), .C(n_404), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_351), .B1(n_375), .B2(n_380), .Y(n_343) );
INVx2_ASAP7_75t_L g1131 ( .A(n_344), .Y(n_1131) );
OR2x6_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
INVx1_ASAP7_75t_L g1027 ( .A(n_345), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1707 ( .A(n_345), .B(n_349), .Y(n_1707) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g563 ( .A(n_346), .Y(n_563) );
INVx1_ASAP7_75t_L g680 ( .A(n_346), .Y(n_680) );
INVx2_ASAP7_75t_SL g858 ( .A(n_346), .Y(n_858) );
BUFx3_ASAP7_75t_L g917 ( .A(n_346), .Y(n_917) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x4_ASAP7_75t_L g378 ( .A(n_347), .B(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_348), .Y(n_379) );
INVx2_ASAP7_75t_L g501 ( .A(n_349), .Y(n_501) );
AND2x4_ASAP7_75t_L g617 ( .A(n_349), .B(n_481), .Y(n_617) );
OR2x2_ASAP7_75t_L g679 ( .A(n_349), .B(n_680), .Y(n_679) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_349), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_349), .B(n_651), .Y(n_1279) );
AND2x4_ASAP7_75t_L g1319 ( .A(n_349), .B(n_481), .Y(n_1319) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g673 ( .A(n_350), .Y(n_673) );
OR2x6_ASAP7_75t_L g719 ( .A(n_350), .B(n_720), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_360), .B1(n_361), .B2(n_365), .C(n_366), .Y(n_351) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OAI221xp5_ASAP7_75t_SL g913 ( .A1(n_353), .A2(n_862), .B1(n_883), .B2(n_886), .C(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g382 ( .A(n_355), .Y(n_382) );
OR2x2_ASAP7_75t_L g582 ( .A(n_355), .B(n_515), .Y(n_582) );
INVx1_ASAP7_75t_L g687 ( .A(n_355), .Y(n_687) );
BUFx2_ASAP7_75t_L g1016 ( .A(n_355), .Y(n_1016) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
AND2x2_ASAP7_75t_L g364 ( .A(n_356), .B(n_358), .Y(n_364) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g373 ( .A(n_357), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g369 ( .A(n_359), .B(n_370), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g472 ( .A1(n_360), .A2(n_365), .B1(n_473), .B2(n_478), .C(n_480), .Y(n_472) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI211xp5_ASAP7_75t_L g765 ( .A1(n_362), .A2(n_715), .B(n_766), .C(n_768), .Y(n_765) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g384 ( .A(n_363), .Y(n_384) );
INVx2_ASAP7_75t_SL g683 ( .A(n_363), .Y(n_683) );
BUFx4f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g517 ( .A(n_364), .Y(n_517) );
INVx1_ASAP7_75t_L g760 ( .A(n_364), .Y(n_760) );
BUFx2_ASAP7_75t_L g846 ( .A(n_364), .Y(n_846) );
INVx1_ASAP7_75t_L g1194 ( .A(n_364), .Y(n_1194) );
INVx1_ASAP7_75t_L g1217 ( .A(n_364), .Y(n_1217) );
BUFx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g522 ( .A(n_368), .Y(n_522) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_368), .B(n_549), .Y(n_1046) );
BUFx4f_ASAP7_75t_L g1137 ( .A(n_368), .Y(n_1137) );
AOI22xp5_ASAP7_75t_L g1339 ( .A1(n_368), .A2(n_574), .B1(n_1335), .B2(n_1340), .Y(n_1339) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_369), .Y(n_388) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_369), .Y(n_560) );
INVx2_ASAP7_75t_SL g694 ( .A(n_369), .Y(n_694) );
BUFx3_ASAP7_75t_L g840 ( .A(n_369), .Y(n_840) );
BUFx6f_ASAP7_75t_L g915 ( .A(n_369), .Y(n_915) );
BUFx2_ASAP7_75t_L g1022 ( .A(n_369), .Y(n_1022) );
BUFx2_ASAP7_75t_L g1198 ( .A(n_369), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1377 ( .A(n_369), .Y(n_1377) );
AND2x2_ASAP7_75t_L g396 ( .A(n_370), .B(n_374), .Y(n_396) );
INVx2_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g1031 ( .A(n_372), .Y(n_1031) );
INVx1_ASAP7_75t_L g1192 ( .A(n_372), .Y(n_1192) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_373), .Y(n_390) );
INVx1_ASAP7_75t_L g513 ( .A(n_373), .Y(n_513) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_373), .Y(n_571) );
INVx2_ASAP7_75t_L g586 ( .A(n_373), .Y(n_586) );
INVx2_ASAP7_75t_L g410 ( .A(n_374), .Y(n_410) );
OAI22xp5_ASAP7_75t_SL g678 ( .A1(n_375), .A2(n_679), .B1(n_681), .B2(n_685), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_375), .A2(n_1212), .B1(n_1213), .B2(n_1222), .Y(n_1211) );
INVx4_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g1126 ( .A1(n_376), .A2(n_1127), .B1(n_1131), .B2(n_1132), .C(n_1140), .Y(n_1126) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AND2x4_ASAP7_75t_L g505 ( .A(n_377), .B(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g951 ( .A(n_377), .B(n_378), .Y(n_951) );
INVx2_ASAP7_75t_L g544 ( .A(n_378), .Y(n_544) );
INVx2_ASAP7_75t_SL g764 ( .A(n_378), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g844 ( .A1(n_378), .A2(n_791), .B1(n_845), .B2(n_847), .C(n_848), .Y(n_844) );
INVx1_ASAP7_75t_L g929 ( .A(n_378), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g1303 ( .A(n_378), .Y(n_1303) );
AND2x4_ASAP7_75t_L g399 ( .A(n_379), .B(n_400), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B1(n_384), .B2(n_385), .C(n_386), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g1652 ( .A1(n_381), .A2(n_1653), .B1(n_1654), .B2(n_1655), .Y(n_1652) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g520 ( .A(n_382), .Y(n_520) );
INVx2_ASAP7_75t_L g682 ( .A(n_382), .Y(n_682) );
INVx2_ASAP7_75t_L g848 ( .A(n_382), .Y(n_848) );
OAI211xp5_ASAP7_75t_L g1664 ( .A1(n_384), .A2(n_1665), .B(n_1666), .C(n_1667), .Y(n_1664) );
BUFx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g547 ( .A(n_388), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_388), .B(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g1654 ( .A(n_390), .Y(n_1654) );
NOR3xp33_ASAP7_75t_SL g1210 ( .A(n_391), .B(n_1211), .C(n_1228), .Y(n_1210) );
BUFx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NOR3xp33_ASAP7_75t_L g676 ( .A(n_392), .B(n_677), .C(n_678), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g952 ( .A1(n_392), .A2(n_953), .B1(n_954), .B2(n_955), .C(n_956), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g1716 ( .A1(n_392), .A2(n_953), .B1(n_955), .B2(n_1717), .C(n_1718), .Y(n_1716) );
AND2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_395), .Y(n_539) );
INVx2_ASAP7_75t_L g856 ( .A(n_395), .Y(n_856) );
BUFx6f_ASAP7_75t_L g1352 ( .A(n_395), .Y(n_1352) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_396), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_397), .B(n_946), .Y(n_1144) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_SL g411 ( .A(n_398), .Y(n_411) );
OR2x6_ASAP7_75t_L g412 ( .A(n_398), .B(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_398), .B(n_413), .Y(n_1143) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
AND2x2_ASAP7_75t_L g506 ( .A(n_399), .B(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g553 ( .A(n_399), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g556 ( .A(n_399), .B(n_414), .Y(n_556) );
INVx1_ASAP7_75t_L g578 ( .A(n_399), .Y(n_578) );
BUFx2_ASAP7_75t_L g754 ( .A(n_399), .Y(n_754) );
AND2x2_ASAP7_75t_L g772 ( .A(n_399), .B(n_414), .Y(n_772) );
AND2x4_ASAP7_75t_L g906 ( .A(n_399), .B(n_554), .Y(n_906) );
AND2x4_ASAP7_75t_L g908 ( .A(n_399), .B(n_414), .Y(n_908) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x6_ASAP7_75t_L g632 ( .A(n_402), .B(n_452), .Y(n_632) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OR2x2_ASAP7_75t_L g514 ( .A(n_403), .B(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g603 ( .A(n_403), .B(n_423), .Y(n_603) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g953 ( .A(n_406), .Y(n_953) );
INVx2_ASAP7_75t_L g1142 ( .A(n_406), .Y(n_1142) );
NAND2x1p5_ASAP7_75t_L g406 ( .A(n_407), .B(n_411), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g554 ( .A(n_408), .Y(n_554) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g507 ( .A(n_410), .B(n_416), .Y(n_507) );
INVx2_ASAP7_75t_L g955 ( .A(n_412), .Y(n_955) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g1307 ( .A1(n_414), .A2(n_554), .B1(n_1308), .B2(n_1309), .Y(n_1307) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI31xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_468), .A3(n_490), .B(n_500), .Y(n_417) );
INVx8_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI221xp5_ASAP7_75t_SL g969 ( .A1(n_420), .A2(n_970), .B1(n_972), .B2(n_975), .C(n_976), .Y(n_969) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_425), .Y(n_420) );
AND2x4_ASAP7_75t_L g497 ( .A(n_421), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g470 ( .A(n_423), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g492 ( .A(n_423), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g453 ( .A(n_424), .Y(n_453) );
INVx1_ASAP7_75t_L g721 ( .A(n_424), .Y(n_721) );
BUFx6f_ASAP7_75t_L g974 ( .A(n_425), .Y(n_974) );
BUFx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_426), .Y(n_450) );
BUFx2_ASAP7_75t_L g597 ( .A(n_426), .Y(n_597) );
BUFx3_ASAP7_75t_L g606 ( .A(n_426), .Y(n_606) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_426), .Y(n_623) );
AND2x4_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_436), .B1(n_437), .B2(n_443), .C(n_444), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
INVx2_ASAP7_75t_L g1172 ( .A(n_431), .Y(n_1172) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_432), .A2(n_966), .B1(n_967), .B2(n_968), .Y(n_965) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g818 ( .A(n_433), .Y(n_818) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g660 ( .A(n_434), .Y(n_660) );
INVx1_ASAP7_75t_L g730 ( .A(n_434), .Y(n_730) );
INVx1_ASAP7_75t_L g467 ( .A(n_435), .Y(n_467) );
AND2x4_ASAP7_75t_L g493 ( .A(n_435), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_440), .Y(n_712) );
AND2x2_ASAP7_75t_L g744 ( .A(n_440), .B(n_603), .Y(n_744) );
INVx1_ASAP7_75t_L g891 ( .A(n_440), .Y(n_891) );
INVx2_ASAP7_75t_L g1082 ( .A(n_440), .Y(n_1082) );
INVx2_ASAP7_75t_L g1087 ( .A(n_440), .Y(n_1087) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g602 ( .A(n_441), .Y(n_602) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_441), .Y(n_647) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g487 ( .A(n_442), .Y(n_487) );
INVx1_ASAP7_75t_L g499 ( .A(n_442), .Y(n_499) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_446), .B(n_460), .Y(n_509) );
AND2x2_ASAP7_75t_L g735 ( .A(n_446), .B(n_603), .Y(n_735) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g610 ( .A(n_447), .Y(n_610) );
INVx2_ASAP7_75t_L g979 ( .A(n_447), .Y(n_979) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_448), .Y(n_471) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_SL g1107 ( .A(n_450), .Y(n_1107) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g651 ( .A(n_452), .Y(n_651) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_464), .B2(n_465), .Y(n_455) );
HB1xp67_ASAP7_75t_L g1241 ( .A(n_457), .Y(n_1241) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
AND2x4_ASAP7_75t_L g589 ( .A(n_458), .B(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g655 ( .A(n_459), .Y(n_655) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OR2x6_ASAP7_75t_L g466 ( .A(n_461), .B(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g488 ( .A(n_461), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g656 ( .A(n_461), .Y(n_656) );
OR2x6_ASAP7_75t_L g670 ( .A(n_461), .B(n_489), .Y(n_670) );
INVx1_ASAP7_75t_L g1737 ( .A(n_461), .Y(n_1737) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_465), .A2(n_1240), .B1(n_1241), .B2(n_1242), .Y(n_1239) );
CKINVDCx11_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g803 ( .A(n_467), .Y(n_803) );
CKINVDCx6p67_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g1724 ( .A1(n_470), .A2(n_1725), .B1(n_1726), .B2(n_1727), .Y(n_1724) );
INVx3_ASAP7_75t_L g620 ( .A(n_471), .Y(n_620) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_471), .Y(n_649) );
BUFx2_ASAP7_75t_L g973 ( .A(n_471), .Y(n_973) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g489 ( .A(n_475), .Y(n_489) );
INVx3_ASAP7_75t_L g665 ( .A(n_475), .Y(n_665) );
INVx2_ASAP7_75t_L g1120 ( .A(n_475), .Y(n_1120) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_476), .B(n_477), .Y(n_718) );
INVx1_ASAP7_75t_L g594 ( .A(n_477), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_478), .A2(n_1089), .B1(n_1394), .B2(n_1395), .Y(n_1393) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OAI221xp5_ASAP7_75t_L g664 ( .A1(n_480), .A2(n_665), .B1(n_666), .B2(n_667), .C(n_669), .Y(n_664) );
BUFx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g1247 ( .A(n_481), .Y(n_1247) );
OAI22xp5_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_484), .B1(n_485), .B2(n_486), .Y(n_482) );
INVx2_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
BUFx3_ASAP7_75t_L g625 ( .A(n_487), .Y(n_625) );
INVx4_ASAP7_75t_L g628 ( .A(n_487), .Y(n_628) );
INVx2_ASAP7_75t_SL g732 ( .A(n_487), .Y(n_732) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_489), .A2(n_667), .B1(n_885), .B2(n_886), .Y(n_884) );
INVx1_ASAP7_75t_L g1090 ( .A(n_489), .Y(n_1090) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_492), .A2(n_497), .B1(n_641), .B2(n_642), .Y(n_640) );
AOI221x1_ASAP7_75t_L g958 ( .A1(n_492), .A2(n_497), .B1(n_959), .B2(n_960), .C(n_961), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_492), .A2(n_497), .B1(n_1110), .B2(n_1111), .Y(n_1109) );
INVx3_ASAP7_75t_L g1254 ( .A(n_492), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g1721 ( .A1(n_492), .A2(n_497), .B1(n_1722), .B2(n_1723), .Y(n_1721) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_493), .Y(n_613) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_493), .Y(n_645) );
BUFx6f_ASAP7_75t_L g971 ( .A(n_493), .Y(n_971) );
INVx1_ASAP7_75t_L g1102 ( .A(n_493), .Y(n_1102) );
INVx1_ASAP7_75t_L g1676 ( .A(n_493), .Y(n_1676) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx3_ASAP7_75t_L g1255 ( .A(n_497), .Y(n_1255) );
INVx1_ASAP7_75t_L g967 ( .A(n_498), .Y(n_967) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g1277 ( .A(n_499), .Y(n_1277) );
AOI31xp33_ASAP7_75t_L g534 ( .A1(n_500), .A2(n_535), .A3(n_557), .B(n_579), .Y(n_534) );
AOI31xp33_ASAP7_75t_SL g1336 ( .A1(n_500), .A2(n_1337), .A3(n_1341), .B(n_1350), .Y(n_1336) );
INVx1_ASAP7_75t_L g1669 ( .A(n_500), .Y(n_1669) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2xp67_ASAP7_75t_L g508 ( .A(n_501), .B(n_509), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g1041 ( .A1(n_501), .A2(n_1042), .B1(n_1058), .B2(n_1059), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_504), .B(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_504), .B(n_1125), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_504), .B(n_1209), .Y(n_1208) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_508), .Y(n_504) );
INVx2_ASAP7_75t_L g532 ( .A(n_505), .Y(n_532) );
AOI222xp33_ASAP7_75t_L g1738 ( .A1(n_505), .A2(n_697), .B1(n_1731), .B2(n_1734), .C1(n_1739), .C2(n_1740), .Y(n_1738) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_506), .B(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g902 ( .A(n_506), .Y(n_902) );
INVx6_ASAP7_75t_L g542 ( .A(n_507), .Y(n_542) );
INVx2_ASAP7_75t_L g699 ( .A(n_507), .Y(n_699) );
BUFx2_ASAP7_75t_L g1030 ( .A(n_507), .Y(n_1030) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_518), .Y(n_510) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
OR2x6_ASAP7_75t_L g702 ( .A(n_513), .B(n_514), .Y(n_702) );
INVx2_ASAP7_75t_L g950 ( .A(n_513), .Y(n_950) );
OR2x6_ASAP7_75t_L g516 ( .A(n_514), .B(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g519 ( .A(n_514), .B(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g521 ( .A(n_514), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g695 ( .A(n_514), .Y(n_695) );
INVx2_ASAP7_75t_L g549 ( .A(n_515), .Y(n_549) );
OR2x2_ASAP7_75t_L g585 ( .A(n_515), .B(n_586), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_515), .A2(n_747), .B(n_750), .C(n_752), .Y(n_746) );
CKINVDCx6p67_ASAP7_75t_R g1743 ( .A(n_516), .Y(n_1743) );
INVx1_ASAP7_75t_L g1225 ( .A(n_517), .Y(n_1225) );
OAI21xp33_ASAP7_75t_L g1292 ( .A1(n_517), .A2(n_1293), .B(n_1294), .Y(n_1292) );
INVx1_ASAP7_75t_L g633 ( .A(n_523), .Y(n_633) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
XNOR2x1_ASAP7_75t_SL g524 ( .A(n_525), .B(n_526), .Y(n_524) );
OAI22xp33_ASAP7_75t_L g1441 ( .A1(n_525), .A2(n_1442), .B1(n_1444), .B2(n_1445), .Y(n_1441) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_587), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_533), .B(n_534), .Y(n_527) );
INVx1_ASAP7_75t_L g869 ( .A(n_528), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g1185 ( .A1(n_528), .A2(n_775), .B1(n_1186), .B2(n_1203), .Y(n_1185) );
INVx5_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g1008 ( .A(n_529), .Y(n_1008) );
INVx2_ASAP7_75t_SL g1059 ( .A(n_529), .Y(n_1059) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
INVx2_ASAP7_75t_L g1326 ( .A(n_530), .Y(n_1326) );
INVx3_ASAP7_75t_L g590 ( .A(n_531), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_545), .B1(n_548), .B2(n_550), .C(n_551), .Y(n_535) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g562 ( .A(n_539), .Y(n_562) );
AND2x4_ASAP7_75t_L g576 ( .A(n_539), .B(n_577), .Y(n_576) );
BUFx6f_ASAP7_75t_L g1199 ( .A(n_539), .Y(n_1199) );
INVx4_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g948 ( .A(n_541), .Y(n_948) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g567 ( .A(n_542), .Y(n_567) );
INVx2_ASAP7_75t_L g748 ( .A(n_542), .Y(n_748) );
INVx1_ASAP7_75t_L g767 ( .A(n_542), .Y(n_767) );
INVx1_ASAP7_75t_L g928 ( .A(n_542), .Y(n_928) );
INVx2_ASAP7_75t_SL g1714 ( .A(n_542), .Y(n_1714) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_548), .Y(n_834) );
AOI211xp5_ASAP7_75t_L g1011 ( .A1(n_548), .A2(n_1012), .B(n_1013), .C(n_1014), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_548), .A2(n_581), .B1(n_1177), .B2(n_1183), .Y(n_1202) );
AND2x4_ASAP7_75t_L g573 ( .A(n_549), .B(n_574), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_549), .A2(n_573), .B1(n_753), .B2(n_896), .C(n_911), .Y(n_910) );
AOI222xp33_ASAP7_75t_L g1337 ( .A1(n_549), .A2(n_906), .B1(n_908), .B2(n_1316), .C1(n_1317), .C2(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_SL g770 ( .A(n_553), .Y(n_770) );
INVx2_ASAP7_75t_SL g836 ( .A(n_553), .Y(n_836) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_564), .B1(n_572), .B2(n_575), .C(n_576), .Y(n_557) );
BUFx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g1191 ( .A(n_560), .Y(n_1191) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx6f_ASAP7_75t_L g1348 ( .A(n_567), .Y(n_1348) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx6f_ASAP7_75t_L g749 ( .A(n_571), .Y(n_749) );
INVx1_ASAP7_75t_L g862 ( .A(n_571), .Y(n_862) );
INVx2_ASAP7_75t_L g912 ( .A(n_571), .Y(n_912) );
INVx1_ASAP7_75t_L g1130 ( .A(n_571), .Y(n_1130) );
HB1xp67_ASAP7_75t_L g1372 ( .A(n_571), .Y(n_1372) );
INVx1_ASAP7_75t_L g851 ( .A(n_572), .Y(n_851) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_572), .A2(n_576), .B1(n_1184), .B2(n_1197), .C(n_1201), .Y(n_1196) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_573), .Y(n_1019) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_573), .A2(n_753), .B1(n_1052), .B2(n_1053), .C(n_1054), .Y(n_1051) );
INVx2_ASAP7_75t_SL g1290 ( .A(n_573), .Y(n_1290) );
BUFx4f_ASAP7_75t_L g751 ( .A(n_574), .Y(n_751) );
AND2x4_ASAP7_75t_L g753 ( .A(n_574), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g927 ( .A(n_574), .Y(n_927) );
BUFx6f_ASAP7_75t_L g946 ( .A(n_574), .Y(n_946) );
INVx2_ASAP7_75t_SL g1345 ( .A(n_574), .Y(n_1345) );
INVx1_ASAP7_75t_L g864 ( .A(n_576), .Y(n_864) );
AOI221xp5_ASAP7_75t_L g1018 ( .A1(n_576), .A2(n_1019), .B1(n_1020), .B2(n_1021), .C(n_1028), .Y(n_1018) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B1(n_583), .B2(n_584), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_581), .A2(n_584), .B1(n_823), .B2(n_826), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_581), .A2(n_584), .B1(n_1033), .B2(n_1034), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_581), .A2(n_584), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
AOI22xp5_ASAP7_75t_L g1364 ( .A1(n_581), .A2(n_584), .B1(n_1365), .B2(n_1366), .Y(n_1364) );
INVx6_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI211xp5_ASAP7_75t_L g1187 ( .A1(n_584), .A2(n_1181), .B(n_1188), .C(n_1189), .Y(n_1187) );
INVx4_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g843 ( .A(n_586), .Y(n_843) );
INVx1_ASAP7_75t_L g1298 ( .A(n_586), .Y(n_1298) );
AND4x1_ASAP7_75t_L g587 ( .A(n_588), .B(n_598), .C(n_607), .D(n_614), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B1(n_592), .B2(n_595), .C(n_596), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g776 ( .A1(n_589), .A2(n_592), .B1(n_596), .B2(n_777), .C(n_778), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_589), .A2(n_596), .B(n_907), .Y(n_936) );
AOI221xp5_ASAP7_75t_L g986 ( .A1(n_589), .A2(n_592), .B1(n_596), .B2(n_987), .C(n_988), .Y(n_986) );
AOI221xp5_ASAP7_75t_L g1315 ( .A1(n_589), .A2(n_592), .B1(n_596), .B2(n_1316), .C(n_1317), .Y(n_1315) );
AOI221xp5_ASAP7_75t_L g1682 ( .A1(n_589), .A2(n_592), .B1(n_596), .B2(n_1662), .C(n_1663), .Y(n_1682) );
AND2x4_ASAP7_75t_L g592 ( .A(n_590), .B(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g596 ( .A(n_590), .B(n_597), .Y(n_596) );
NAND2x1_ASAP7_75t_SL g799 ( .A(n_590), .B(n_654), .Y(n_799) );
NAND2x1p5_ASAP7_75t_L g802 ( .A(n_590), .B(n_803), .Y(n_802) );
NAND2x1p5_ASAP7_75t_L g804 ( .A(n_590), .B(n_606), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g1736 ( .A1(n_593), .A2(n_654), .B1(n_1717), .B2(n_1718), .Y(n_1736) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g1003 ( .A(n_597), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_597), .A2(n_610), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B1(n_604), .B2(n_605), .Y(n_598) );
BUFx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx2_ASAP7_75t_L g795 ( .A(n_601), .Y(n_795) );
BUFx2_ASAP7_75t_L g935 ( .A(n_601), .Y(n_935) );
BUFx2_ASAP7_75t_L g995 ( .A(n_601), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_601), .A2(n_605), .B1(n_1063), .B2(n_1064), .Y(n_1062) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx1_ASAP7_75t_L g662 ( .A(n_602), .Y(n_662) );
BUFx3_ASAP7_75t_L g821 ( .A(n_602), .Y(n_821) );
INVx2_ASAP7_75t_L g1117 ( .A(n_602), .Y(n_1117) );
INVx1_ASAP7_75t_SL g1272 ( .A(n_602), .Y(n_1272) );
AND2x6_ASAP7_75t_L g605 ( .A(n_603), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g609 ( .A(n_603), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g612 ( .A(n_603), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g739 ( .A(n_603), .B(n_613), .Y(n_739) );
AND2x2_ASAP7_75t_L g741 ( .A(n_603), .B(n_623), .Y(n_741) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_603), .B(n_613), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_603), .B(n_613), .Y(n_1160) );
AOI22xp5_ASAP7_75t_L g1327 ( .A1(n_603), .A2(n_1279), .B1(n_1328), .B2(n_1332), .Y(n_1327) );
BUFx2_ASAP7_75t_L g789 ( .A(n_605), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_605), .A2(n_795), .B1(n_1155), .B2(n_1156), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1237 ( .A(n_606), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_611), .B2(n_612), .Y(n_607) );
BUFx2_ASAP7_75t_L g792 ( .A(n_609), .Y(n_792) );
INVx1_ASAP7_75t_L g933 ( .A(n_609), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_609), .A2(n_1066), .B1(n_1067), .B2(n_1068), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_609), .A2(n_1158), .B1(n_1159), .B2(n_1160), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_609), .A2(n_739), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
AOI221xp5_ASAP7_75t_L g1683 ( .A1(n_609), .A2(n_1160), .B1(n_1684), .B2(n_1685), .C(n_1686), .Y(n_1683) );
BUFx3_ASAP7_75t_L g630 ( .A(n_610), .Y(n_630) );
INVx1_ASAP7_75t_L g1105 ( .A(n_610), .Y(n_1105) );
BUFx2_ASAP7_75t_L g1673 ( .A(n_610), .Y(n_1673) );
INVx1_ASAP7_75t_L g787 ( .A(n_612), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_612), .A2(n_789), .B1(n_990), .B2(n_991), .Y(n_989) );
AOI33xp33_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_618), .A3(n_624), .B1(n_626), .B2(n_629), .B3(n_631), .Y(n_614) );
AOI33xp33_ASAP7_75t_L g996 ( .A1(n_615), .A2(n_997), .A3(n_1001), .B1(n_1004), .B2(n_1005), .B3(n_1006), .Y(n_996) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g1681 ( .A(n_620), .Y(n_1681) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
OAI22xp33_ASAP7_75t_L g880 ( .A1(n_628), .A2(n_881), .B1(n_882), .B2(n_883), .Y(n_880) );
OAI221xp5_ASAP7_75t_L g1232 ( .A1(n_628), .A2(n_1233), .B1(n_1234), .B2(n_1235), .C(n_1236), .Y(n_1232) );
INVx1_ASAP7_75t_L g733 ( .A(n_631), .Y(n_733) );
INVx2_ASAP7_75t_L g897 ( .A(n_631), .Y(n_897) );
INVx6_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx5_ASAP7_75t_L g830 ( .A(n_632), .Y(n_830) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
XNOR2x1_ASAP7_75t_L g635 ( .A(n_636), .B(n_705), .Y(n_635) );
INVx1_ASAP7_75t_L g703 ( .A(n_637), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g637 ( .A(n_638), .B(n_674), .C(n_676), .D(n_691), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_657), .B(n_671), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_648), .B(n_652), .Y(n_643) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_645), .Y(n_1002) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g1175 ( .A(n_647), .Y(n_1175) );
INVx2_ASAP7_75t_L g1321 ( .A(n_647), .Y(n_1321) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g1238 ( .A(n_651), .Y(n_1238) );
NAND2x1p5_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g708 ( .A1(n_659), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_708) );
BUFx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g890 ( .A(n_660), .Y(n_890) );
OAI21xp5_ASAP7_75t_SL g962 ( .A1(n_665), .A2(n_963), .B(n_964), .Y(n_962) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_666), .A2(n_669), .B1(n_682), .B2(n_683), .C(n_684), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_667), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g1166 ( .A1(n_667), .A2(n_1167), .B1(n_1168), .B2(n_1169), .Y(n_1166) );
OAI22xp33_ASAP7_75t_L g1182 ( .A1(n_667), .A2(n_1169), .B1(n_1183), .B2(n_1184), .Y(n_1182) );
OAI221xp5_ASAP7_75t_L g1244 ( .A1(n_667), .A2(n_1214), .B1(n_1218), .B2(n_1245), .C(n_1246), .Y(n_1244) );
INVx3_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g961 ( .A1(n_670), .A2(n_962), .B(n_965), .Y(n_961) );
INVx5_ASAP7_75t_L g866 ( .A(n_671), .Y(n_866) );
OAI21xp5_ASAP7_75t_L g1719 ( .A1(n_671), .A2(n_1720), .B(n_1728), .Y(n_1719) );
BUFx8_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
AOI31xp33_ASAP7_75t_L g1010 ( .A1(n_672), .A2(n_1011), .A3(n_1018), .B(n_1032), .Y(n_1010) );
INVx2_ASAP7_75t_L g1311 ( .A(n_672), .Y(n_1311) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx2_ASAP7_75t_L g775 ( .A(n_673), .Y(n_775) );
INVx3_ASAP7_75t_L g942 ( .A(n_679), .Y(n_942) );
OAI221xp5_ASAP7_75t_L g1193 ( .A1(n_682), .A2(n_1156), .B1(n_1158), .B2(n_1194), .C(n_1195), .Y(n_1193) );
OAI221xp5_ASAP7_75t_L g685 ( .A1(n_683), .A2(n_686), .B1(n_688), .B2(n_689), .C(n_690), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g1656 ( .A1(n_683), .A2(n_1657), .B(n_1658), .Y(n_1656) );
OAI22xp5_ASAP7_75t_L g1295 ( .A1(n_686), .A2(n_1273), .B1(n_1296), .B2(n_1297), .Y(n_1295) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_696), .B1(n_697), .B2(n_700), .C(n_701), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g1145 ( .A1(n_692), .A2(n_697), .B1(n_1146), .B2(n_1147), .C(n_1148), .Y(n_1145) );
AOI22xp5_ASAP7_75t_L g1741 ( .A1(n_692), .A2(n_1732), .B1(n_1742), .B2(n_1743), .Y(n_1741) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_693), .A2(n_725), .B1(n_727), .B2(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_SL g944 ( .A(n_694), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_694), .A2(n_1116), .B1(n_1118), .B2(n_1130), .Y(n_1129) );
INVx1_ASAP7_75t_L g1343 ( .A(n_694), .Y(n_1343) );
AND2x2_ASAP7_75t_L g697 ( .A(n_695), .B(n_698), .Y(n_697) );
BUFx2_ASAP7_75t_L g860 ( .A(n_698), .Y(n_860) );
A2O1A1Ixp33_ASAP7_75t_L g1304 ( .A1(n_698), .A2(n_1305), .B(n_1306), .C(n_1310), .Y(n_1304) );
INVx2_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g763 ( .A(n_699), .Y(n_763) );
CKINVDCx6p67_ASAP7_75t_R g1740 ( .A(n_702), .Y(n_1740) );
INVx1_ASAP7_75t_SL g780 ( .A(n_706), .Y(n_780) );
NAND4xp75_ASAP7_75t_L g706 ( .A(n_707), .B(n_736), .C(n_745), .D(n_776), .Y(n_706) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
BUFx3_ASAP7_75t_L g827 ( .A(n_716), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g1073 ( .A1(n_716), .A2(n_1074), .B1(n_1077), .B2(n_1078), .Y(n_1073) );
BUFx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_717), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
INVx2_ASAP7_75t_L g813 ( .A(n_717), .Y(n_813) );
BUFx3_ASAP7_75t_L g1169 ( .A(n_717), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1735 ( .A(n_717), .B(n_1736), .Y(n_1735) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_719), .Y(n_806) );
OAI33xp33_ASAP7_75t_L g1072 ( .A1(n_719), .A2(n_829), .A3(n_1073), .B1(n_1079), .B2(n_1084), .B3(n_1088), .Y(n_1072) );
INVx1_ASAP7_75t_L g1165 ( .A(n_719), .Y(n_1165) );
OAI33xp33_ASAP7_75t_L g1392 ( .A1(n_719), .A2(n_897), .A3(n_1393), .B1(n_1396), .B2(n_1400), .B3(n_1402), .Y(n_1392) );
OAI22xp33_ASAP7_75t_L g1402 ( .A1(n_723), .A2(n_1169), .B1(n_1365), .B2(n_1369), .Y(n_1402) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_724), .A2(n_731), .B1(n_748), .B2(n_749), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_731), .B2(n_732), .Y(n_726) );
BUFx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
BUFx2_ASAP7_75t_L g1080 ( .A(n_729), .Y(n_1080) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
HB1xp67_ASAP7_75t_L g1115 ( .A(n_730), .Y(n_1115) );
INVx1_ASAP7_75t_L g1180 ( .A(n_730), .Y(n_1180) );
INVx2_ASAP7_75t_L g1233 ( .A(n_730), .Y(n_1233) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NOR2x1_ASAP7_75t_L g736 ( .A(n_737), .B(n_742), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g877 ( .A(n_739), .Y(n_877) );
INVx1_ASAP7_75t_L g1283 ( .A(n_739), .Y(n_1283) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g1284 ( .A(n_741), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_741), .A2(n_744), .B1(n_1386), .B2(n_1387), .Y(n_1385) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OAI31xp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_755), .A3(n_769), .B(n_775), .Y(n_745) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_748), .Y(n_1128) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g1341 ( .A1(n_753), .A2(n_1342), .B(n_1347), .Y(n_1341) );
AOI221xp5_ASAP7_75t_L g1367 ( .A1(n_753), .A2(n_1368), .B1(n_1369), .B2(n_1370), .C(n_1371), .Y(n_1367) );
INVx1_ASAP7_75t_L g1659 ( .A(n_753), .Y(n_1659) );
BUFx3_ASAP7_75t_L g1310 ( .A(n_754), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_765), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B(n_761), .C(n_762), .Y(n_756) );
OAI221xp5_ASAP7_75t_L g1015 ( .A1(n_758), .A2(n_991), .B1(n_993), .B2(n_1016), .C(n_1017), .Y(n_1015) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp33_ASAP7_75t_L g1306 ( .A(n_760), .B(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1195 ( .A(n_764), .Y(n_1195) );
INVx3_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g931 ( .A(n_775), .Y(n_931) );
AOI21x1_ASAP7_75t_L g957 ( .A1(n_775), .A2(n_958), .B(n_969), .Y(n_957) );
AO22x2_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_1037), .B1(n_1260), .B2(n_1261), .Y(n_781) );
INVx1_ASAP7_75t_L g1260 ( .A(n_782), .Y(n_1260) );
XNOR2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_870), .Y(n_782) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_831), .Y(n_784) );
NOR3xp33_ASAP7_75t_SL g785 ( .A(n_786), .B(n_796), .C(n_805), .Y(n_785) );
INVxp67_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_792), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_992) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_SL g1162 ( .A(n_798), .Y(n_1162) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_799), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx4f_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
BUFx4f_ASAP7_75t_L g878 ( .A(n_802), .Y(n_878) );
BUFx3_ASAP7_75t_L g1071 ( .A(n_804), .Y(n_1071) );
OAI33xp33_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_807), .A3(n_814), .B1(n_822), .B2(n_825), .B3(n_829), .Y(n_805) );
OAI22xp5_ASAP7_75t_SL g807 ( .A1(n_808), .A2(n_809), .B1(n_811), .B2(n_812), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g822 ( .A1(n_809), .A2(n_816), .B1(n_823), .B2(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g895 ( .A(n_810), .Y(n_895) );
OAI22xp5_ASAP7_75t_SL g893 ( .A1(n_812), .A2(n_894), .B1(n_895), .B2(n_896), .Y(n_893) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g1245 ( .A(n_813), .Y(n_1245) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B1(n_819), .B2(n_820), .Y(n_814) );
BUFx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_L g882 ( .A(n_818), .Y(n_882) );
INVx2_ASAP7_75t_L g1397 ( .A(n_818), .Y(n_1397) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_820), .A2(n_826), .B1(n_827), .B2(n_828), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_820), .A2(n_1177), .B1(n_1178), .B2(n_1181), .Y(n_1176) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_821), .Y(n_1000) );
AOI211xp5_ASAP7_75t_L g833 ( .A1(n_824), .A2(n_834), .B(n_835), .C(n_837), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g849 ( .A1(n_828), .A2(n_850), .B1(n_852), .B2(n_859), .C(n_863), .Y(n_849) );
INVx1_ASAP7_75t_L g1006 ( .A(n_829), .Y(n_1006) );
OAI33xp33_ASAP7_75t_L g1163 ( .A1(n_829), .A2(n_1164), .A3(n_1166), .B1(n_1170), .B2(n_1176), .B3(n_1182), .Y(n_1163) );
CKINVDCx8_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
AOI22xp33_ASAP7_75t_SL g831 ( .A1(n_832), .A2(n_866), .B1(n_867), .B2(n_868), .Y(n_831) );
NAND3xp33_ASAP7_75t_L g832 ( .A(n_833), .B(n_849), .C(n_865), .Y(n_832) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
BUFx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx2_ASAP7_75t_SL g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g923 ( .A(n_842), .Y(n_923) );
INVx1_ASAP7_75t_L g1709 ( .A(n_842), .Y(n_1709) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_843), .Y(n_1221) );
INVx2_ASAP7_75t_SL g845 ( .A(n_846), .Y(n_845) );
OAI221xp5_ASAP7_75t_L g1213 ( .A1(n_848), .A2(n_1214), .B1(n_1215), .B2(n_1218), .C(n_1219), .Y(n_1213) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx3_ASAP7_75t_L g1025 ( .A(n_856), .Y(n_1025) );
BUFx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g1139 ( .A(n_862), .Y(n_1139) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_SL g1256 ( .A(n_866), .Y(n_1256) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_983), .B2(n_1036), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
AO22x2_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_937), .B1(n_938), .B2(n_982), .Y(n_872) );
INVx1_ASAP7_75t_L g982 ( .A(n_873), .Y(n_982) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_898), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_879), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .B1(n_891), .B2(n_892), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_889), .A2(n_1249), .B1(n_1250), .B2(n_1252), .Y(n_1248) );
INVx2_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g1251 ( .A(n_891), .Y(n_1251) );
AOI21xp5_ASAP7_75t_SL g898 ( .A1(n_899), .A2(n_930), .B(n_932), .Y(n_898) );
NAND4xp25_ASAP7_75t_SL g899 ( .A(n_900), .B(n_910), .C(n_913), .D(n_918), .Y(n_899) );
AOI222xp33_ASAP7_75t_SL g900 ( .A1(n_901), .A2(n_903), .B1(n_904), .B2(n_907), .C1(n_908), .C2(n_909), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g1350 ( .A1(n_901), .A2(n_1325), .B1(n_1351), .B2(n_1353), .Y(n_1350) );
INVx2_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
INVx4_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx2_ASAP7_75t_L g1049 ( .A(n_906), .Y(n_1049) );
INVx1_ASAP7_75t_SL g1380 ( .A(n_906), .Y(n_1380) );
AOI22xp5_ASAP7_75t_L g1661 ( .A1(n_906), .A2(n_908), .B1(n_1662), .B2(n_1663), .Y(n_1661) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_908), .Y(n_1050) );
BUFx3_ASAP7_75t_L g920 ( .A(n_915), .Y(n_920) );
INVx3_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g1200 ( .A(n_917), .Y(n_1200) );
INVxp67_ASAP7_75t_L g1346 ( .A(n_917), .Y(n_1346) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_919), .A2(n_921), .B1(n_922), .B2(n_924), .C(n_925), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx1_ASAP7_75t_L g1017 ( .A(n_929), .Y(n_1017) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
NOR4xp75_ASAP7_75t_L g939 ( .A(n_940), .B(n_957), .C(n_980), .D(n_981), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_941), .B(n_952), .Y(n_940) );
AOI33xp33_ASAP7_75t_L g941 ( .A1(n_942), .A2(n_943), .A3(n_945), .B1(n_947), .B2(n_949), .B3(n_951), .Y(n_941) );
INVx1_ASAP7_75t_L g1134 ( .A(n_946), .Y(n_1134) );
AOI33xp33_ASAP7_75t_L g1705 ( .A1(n_951), .A2(n_1706), .A3(n_1708), .B1(n_1710), .B2(n_1711), .B3(n_1715), .Y(n_1705) );
INVx2_ASAP7_75t_L g1229 ( .A(n_953), .Y(n_1229) );
INVx1_ASAP7_75t_L g1679 ( .A(n_967), .Y(n_1679) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
BUFx3_ASAP7_75t_L g998 ( .A(n_979), .Y(n_998) );
INVx2_ASAP7_75t_L g1036 ( .A(n_983), .Y(n_1036) );
XOR2x2_ASAP7_75t_L g983 ( .A(n_984), .B(n_1035), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_1007), .Y(n_984) );
AND4x1_ASAP7_75t_L g985 ( .A(n_986), .B(n_989), .C(n_992), .D(n_996), .Y(n_985) );
INVx1_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
AOI21xp5_ASAP7_75t_L g1007 ( .A1(n_1008), .A2(n_1009), .B(n_1010), .Y(n_1007) );
OAI221xp5_ASAP7_75t_L g1222 ( .A1(n_1016), .A2(n_1223), .B1(n_1224), .B2(n_1226), .C(n_1227), .Y(n_1222) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1037), .Y(n_1261) );
XNOR2xp5_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1093), .Y(n_1037) );
INVx3_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1040), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_1041), .B(n_1060), .Y(n_1040) );
NAND3xp33_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1051), .C(n_1055), .Y(n_1042) );
AOI221xp5_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1045), .B1(n_1046), .B2(n_1047), .C(n_1048), .Y(n_1043) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1046), .Y(n_1288) );
AOI221xp5_ASAP7_75t_L g1373 ( .A1(n_1046), .A2(n_1374), .B1(n_1375), .B2(n_1376), .C(n_1379), .Y(n_1373) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_1047), .A2(n_1057), .B1(n_1080), .B2(n_1085), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g1088 ( .A1(n_1054), .A2(n_1056), .B1(n_1074), .B2(n_1089), .Y(n_1088) );
AOI22xp5_ASAP7_75t_L g1362 ( .A1(n_1059), .A2(n_1363), .B1(n_1381), .B2(n_1382), .Y(n_1362) );
NOR3xp33_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1069), .C(n_1072), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1065), .Y(n_1061) );
INVx2_ASAP7_75t_SL g1074 ( .A(n_1075), .Y(n_1074) );
INVx2_ASAP7_75t_SL g1075 ( .A(n_1076), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1081), .B1(n_1082), .B2(n_1083), .Y(n_1079) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1677 ( .A(n_1087), .Y(n_1677) );
OAI22xp5_ASAP7_75t_L g1730 ( .A1(n_1087), .A2(n_1233), .B1(n_1731), .B2(n_1732), .Y(n_1730) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
XOR2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1204), .Y(n_1093) );
XNOR2xp5_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1149), .Y(n_1094) );
NAND4xp25_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1124), .C(n_1126), .D(n_1145), .Y(n_1096) );
OAI21xp5_ASAP7_75t_SL g1097 ( .A1(n_1098), .A2(n_1112), .B(n_1123), .Y(n_1097) );
AOI21xp5_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1103), .B(n_1108), .Y(n_1099) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_1110), .A2(n_1111), .B1(n_1136), .B2(n_1138), .Y(n_1135) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_1114), .A2(n_1116), .B1(n_1117), .B2(n_1118), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1400 ( .A1(n_1114), .A2(n_1366), .B1(n_1374), .B2(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_1117), .A2(n_1397), .B1(n_1398), .B2(n_1399), .Y(n_1396) );
OAI21xp5_ASAP7_75t_SL g1119 ( .A1(n_1120), .A2(n_1121), .B(n_1122), .Y(n_1119) );
CKINVDCx8_ASAP7_75t_R g1381 ( .A(n_1123), .Y(n_1381) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1130), .Y(n_1349) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1130), .Y(n_1378) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1131), .Y(n_1212) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
XNOR2x1_ASAP7_75t_SL g1149 ( .A(n_1150), .B(n_1151), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1185), .Y(n_1151) );
NOR3xp33_ASAP7_75t_SL g1152 ( .A(n_1153), .B(n_1161), .C(n_1163), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1157), .Y(n_1153) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_1171), .A2(n_1172), .B1(n_1173), .B2(n_1174), .Y(n_1170) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
OAI221xp5_ASAP7_75t_L g1270 ( .A1(n_1180), .A2(n_1271), .B1(n_1272), .B2(n_1273), .C(n_1274), .Y(n_1270) );
NAND3xp33_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1196), .C(n_1202), .Y(n_1186) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
OAI211xp5_ASAP7_75t_L g1299 ( .A1(n_1194), .A2(n_1300), .B(n_1301), .C(n_1302), .Y(n_1299) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
XNOR2xp5_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1207), .Y(n_1205) );
AND4x1_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1210), .C(n_1230), .D(n_1257), .Y(n_1207) );
INVx2_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
HB1xp67_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
OAI31xp33_ASAP7_75t_L g1230 ( .A1(n_1231), .A2(n_1243), .A3(n_1253), .B(n_1256), .Y(n_1230) );
INVx2_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx2_ASAP7_75t_SL g1250 ( .A(n_1251), .Y(n_1250) );
NOR2xp33_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1259), .Y(n_1257) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
XNOR2xp5_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1358), .Y(n_1263) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
XNOR2xp5_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1312), .Y(n_1265) );
NAND3xp33_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1281), .C(n_1286), .Y(n_1267) );
NOR2xp33_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1280), .Y(n_1268) );
NAND3xp33_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1278), .C(n_1279), .Y(n_1275) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1277), .Y(n_1401) );
AOI33xp33_ASAP7_75t_L g1671 ( .A1(n_1279), .A2(n_1319), .A3(n_1672), .B1(n_1674), .B2(n_1678), .B3(n_1680), .Y(n_1671) );
NOR2xp33_ASAP7_75t_SL g1281 ( .A(n_1282), .B(n_1285), .Y(n_1281) );
OAI31xp33_ASAP7_75t_SL g1286 ( .A1(n_1287), .A2(n_1289), .A3(n_1291), .B(n_1311), .Y(n_1286) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1290), .Y(n_1368) );
OAI211xp5_ASAP7_75t_SL g1291 ( .A1(n_1292), .A2(n_1295), .B(n_1299), .C(n_1304), .Y(n_1291) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
NAND2xp5_ASAP7_75t_SL g1312 ( .A(n_1313), .B(n_1354), .Y(n_1312) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1314), .Y(n_1356) );
NAND3xp33_ASAP7_75t_SL g1314 ( .A(n_1315), .B(n_1318), .C(n_1327), .Y(n_1314) );
AOI22xp5_ASAP7_75t_L g1318 ( .A1(n_1319), .A2(n_1320), .B1(n_1325), .B2(n_1326), .Y(n_1318) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1336), .Y(n_1355) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
NAND3xp33_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1356), .C(n_1357), .Y(n_1354) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
HB1xp67_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1361), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1383), .Y(n_1361) );
NAND3xp33_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1367), .C(n_1373), .Y(n_1363) );
NOR3xp33_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1391), .C(n_1392), .Y(n_1383) );
NAND2xp5_ASAP7_75t_SL g1384 ( .A(n_1385), .B(n_1388), .Y(n_1384) );
OAI221xp5_ASAP7_75t_L g1405 ( .A1(n_1406), .A2(n_1643), .B1(n_1644), .B2(n_1687), .C(n_1692), .Y(n_1405) );
AOI211xp5_ASAP7_75t_L g1406 ( .A1(n_1407), .A2(n_1554), .B(n_1596), .C(n_1622), .Y(n_1406) );
NAND5xp2_ASAP7_75t_L g1407 ( .A(n_1408), .B(n_1516), .C(n_1541), .D(n_1546), .E(n_1551), .Y(n_1407) );
AOI21xp5_ASAP7_75t_L g1408 ( .A1(n_1409), .A2(n_1487), .B(n_1495), .Y(n_1408) );
OAI211xp5_ASAP7_75t_L g1409 ( .A1(n_1410), .A2(n_1447), .B(n_1457), .C(n_1481), .Y(n_1409) );
INVxp67_ASAP7_75t_SL g1410 ( .A(n_1411), .Y(n_1410) );
NOR2xp33_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1436), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
AOI22xp5_ASAP7_75t_L g1577 ( .A1(n_1413), .A2(n_1472), .B1(n_1578), .B2(n_1579), .Y(n_1577) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1433), .Y(n_1413) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1414), .Y(n_1483) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1414), .B(n_1499), .Y(n_1505) );
NAND2xp5_ASAP7_75t_L g1539 ( .A(n_1414), .B(n_1437), .Y(n_1539) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1414), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1414), .B(n_1488), .Y(n_1584) );
AOI221xp5_ASAP7_75t_L g1585 ( .A1(n_1414), .A2(n_1558), .B1(n_1586), .B2(n_1589), .C(n_1593), .Y(n_1585) );
INVx1_ASAP7_75t_L g1604 ( .A(n_1414), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1415), .B(n_1427), .Y(n_1414) );
AND2x4_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1422), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
OR2x2_ASAP7_75t_L g1443 ( .A(n_1418), .B(n_1423), .Y(n_1443) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1421), .Y(n_1418) );
HB1xp67_ASAP7_75t_L g1748 ( .A(n_1419), .Y(n_1748) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1421), .Y(n_1430) );
AND2x4_ASAP7_75t_L g1424 ( .A(n_1422), .B(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1423), .B(n_1426), .Y(n_1446) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
BUFx3_ASAP7_75t_L g1462 ( .A(n_1428), .Y(n_1462) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1428), .Y(n_1492) );
AND2x4_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1431), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1429), .B(n_1431), .Y(n_1453) );
HB1xp67_ASAP7_75t_L g1749 ( .A(n_1429), .Y(n_1749) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
AND2x4_ASAP7_75t_L g1432 ( .A(n_1430), .B(n_1431), .Y(n_1432) );
INVx2_ASAP7_75t_L g1440 ( .A(n_1432), .Y(n_1440) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1433), .Y(n_1480) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1433), .Y(n_1499) );
BUFx6f_ASAP7_75t_L g1537 ( .A(n_1433), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1433), .B(n_1483), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1619 ( .A(n_1433), .B(n_1489), .Y(n_1619) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1435), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1436), .B(n_1515), .Y(n_1566) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1436), .Y(n_1574) );
NAND2xp5_ASAP7_75t_L g1597 ( .A(n_1436), .B(n_1526), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1642 ( .A(n_1436), .B(n_1498), .Y(n_1642) );
BUFx3_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx2_ASAP7_75t_SL g1471 ( .A(n_1437), .Y(n_1471) );
NOR2xp33_ASAP7_75t_L g1482 ( .A(n_1437), .B(n_1483), .Y(n_1482) );
BUFx2_ASAP7_75t_L g1523 ( .A(n_1437), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1534 ( .A(n_1437), .B(n_1454), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1557 ( .A(n_1437), .B(n_1558), .Y(n_1557) );
INVx2_ASAP7_75t_SL g1437 ( .A(n_1438), .Y(n_1437) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1438), .B(n_1503), .Y(n_1561) );
AND2x2_ASAP7_75t_L g1636 ( .A(n_1438), .B(n_1483), .Y(n_1636) );
INVx2_ASAP7_75t_L g1439 ( .A(n_1440), .Y(n_1439) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1440), .Y(n_1463) );
OAI22xp5_ASAP7_75t_SL g1491 ( .A1(n_1440), .A2(n_1492), .B1(n_1493), .B2(n_1494), .Y(n_1491) );
BUFx3_ASAP7_75t_L g1466 ( .A(n_1442), .Y(n_1466) );
BUFx6f_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
HB1xp67_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1446), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1447), .B(n_1518), .Y(n_1517) );
NOR2xp33_ASAP7_75t_L g1593 ( .A(n_1447), .B(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
AOI221xp5_ASAP7_75t_L g1556 ( .A1(n_1448), .A2(n_1505), .B1(n_1531), .B2(n_1557), .C(n_1559), .Y(n_1556) );
A2O1A1Ixp33_ASAP7_75t_SL g1573 ( .A1(n_1448), .A2(n_1512), .B(n_1574), .C(n_1575), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1449), .B(n_1454), .Y(n_1448) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1449), .Y(n_1507) );
OR2x2_ASAP7_75t_L g1580 ( .A(n_1449), .B(n_1454), .Y(n_1580) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1450), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1450), .B(n_1475), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_1450), .B(n_1476), .Y(n_1527) );
INVxp67_ASAP7_75t_SL g1533 ( .A(n_1450), .Y(n_1533) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_1450), .B(n_1454), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1451), .B(n_1452), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1454), .B(n_1473), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1454), .B(n_1485), .Y(n_1484) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_1454), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1454), .B(n_1532), .Y(n_1549) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1454), .B(n_1527), .Y(n_1553) );
NOR2xp33_ASAP7_75t_L g1564 ( .A(n_1454), .B(n_1474), .Y(n_1564) );
NOR2xp33_ASAP7_75t_L g1571 ( .A(n_1454), .B(n_1507), .Y(n_1571) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1454), .B(n_1510), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1454), .B(n_1474), .Y(n_1613) );
HB1xp67_ASAP7_75t_L g1625 ( .A(n_1454), .Y(n_1625) );
AND2x4_ASAP7_75t_SL g1454 ( .A(n_1455), .B(n_1456), .Y(n_1454) );
OAI21xp5_ASAP7_75t_SL g1457 ( .A1(n_1458), .A2(n_1470), .B(n_1479), .Y(n_1457) );
OAI221xp5_ASAP7_75t_L g1576 ( .A1(n_1458), .A2(n_1489), .B1(n_1577), .B2(n_1581), .C(n_1583), .Y(n_1576) );
INVx2_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1459), .B(n_1480), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1487 ( .A(n_1459), .B(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1462), .Y(n_1643) );
OAI22xp33_ASAP7_75t_L g1464 ( .A1(n_1465), .A2(n_1466), .B1(n_1467), .B2(n_1468), .Y(n_1464) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
OAI31xp33_ASAP7_75t_L g1598 ( .A1(n_1470), .A2(n_1542), .A3(n_1599), .B(n_1601), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1471), .B(n_1472), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1509 ( .A(n_1471), .B(n_1510), .Y(n_1509) );
HB1xp67_ASAP7_75t_L g1514 ( .A(n_1471), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1471), .B(n_1564), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1471), .B(n_1498), .Y(n_1595) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1475), .B(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1532 ( .A(n_1476), .B(n_1533), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1478), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1480), .B(n_1489), .Y(n_1520) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1480), .Y(n_1535) );
OAI32xp33_ASAP7_75t_L g1559 ( .A1(n_1480), .A2(n_1510), .A3(n_1537), .B1(n_1560), .B2(n_1562), .Y(n_1559) );
OR2x2_ASAP7_75t_L g1605 ( .A(n_1480), .B(n_1489), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1609 ( .A(n_1480), .B(n_1488), .Y(n_1609) );
NAND2xp5_ASAP7_75t_L g1481 ( .A(n_1482), .B(n_1484), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1483), .B(n_1499), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1483), .B(n_1488), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1515 ( .A(n_1485), .B(n_1503), .Y(n_1515) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1485), .Y(n_1629) );
NAND2xp5_ASAP7_75t_SL g1497 ( .A(n_1488), .B(n_1498), .Y(n_1497) );
AOI32xp33_ASAP7_75t_L g1500 ( .A1(n_1488), .A2(n_1489), .A3(n_1501), .B1(n_1506), .B2(n_1508), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1488), .B(n_1545), .Y(n_1632) );
CKINVDCx6p67_ASAP7_75t_R g1488 ( .A(n_1489), .Y(n_1488) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1489), .B(n_1505), .Y(n_1550) );
CKINVDCx5p33_ASAP7_75t_R g1555 ( .A(n_1489), .Y(n_1555) );
NAND2xp5_ASAP7_75t_L g1635 ( .A(n_1489), .B(n_1636), .Y(n_1635) );
OR2x6_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1491), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g1495 ( .A1(n_1496), .A2(n_1500), .B1(n_1511), .B2(n_1513), .Y(n_1495) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1498), .Y(n_1528) );
AOI211xp5_ASAP7_75t_L g1565 ( .A1(n_1498), .A2(n_1566), .B(n_1567), .C(n_1576), .Y(n_1565) );
INVxp67_ASAP7_75t_SL g1501 ( .A(n_1502), .Y(n_1501) );
NAND2xp5_ASAP7_75t_L g1502 ( .A(n_1503), .B(n_1504), .Y(n_1502) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_1503), .B(n_1510), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1503), .B(n_1527), .Y(n_1526) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1503), .B(n_1532), .Y(n_1542) );
OR2x2_ASAP7_75t_L g1592 ( .A(n_1503), .B(n_1509), .Y(n_1592) );
OR2x2_ASAP7_75t_L g1630 ( .A(n_1503), .B(n_1587), .Y(n_1630) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
OAI21xp5_ASAP7_75t_SL g1541 ( .A1(n_1510), .A2(n_1542), .B(n_1543), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1611 ( .A(n_1510), .B(n_1534), .Y(n_1611) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_1514), .B(n_1515), .Y(n_1513) );
AOI311xp33_ASAP7_75t_L g1516 ( .A1(n_1517), .A2(n_1520), .A3(n_1521), .B(n_1524), .C(n_1529), .Y(n_1516) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
NAND2xp5_ASAP7_75t_L g1551 ( .A(n_1520), .B(n_1552), .Y(n_1551) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1520), .Y(n_1614) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1522), .B(n_1553), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1522), .B(n_1571), .Y(n_1570) );
INVx2_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
NAND2xp5_ASAP7_75t_L g1544 ( .A(n_1523), .B(n_1545), .Y(n_1544) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_1523), .B(n_1527), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1578 ( .A(n_1523), .B(n_1535), .Y(n_1578) );
OR2x2_ASAP7_75t_L g1587 ( .A(n_1523), .B(n_1588), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1591 ( .A(n_1523), .B(n_1571), .Y(n_1591) );
OR2x2_ASAP7_75t_L g1600 ( .A(n_1523), .B(n_1540), .Y(n_1600) );
NOR2xp33_ASAP7_75t_L g1524 ( .A(n_1525), .B(n_1528), .Y(n_1524) );
OAI22xp5_ASAP7_75t_L g1640 ( .A1(n_1525), .A2(n_1537), .B1(n_1641), .B2(n_1642), .Y(n_1640) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
OAI21xp33_ASAP7_75t_L g1569 ( .A1(n_1526), .A2(n_1570), .B(n_1572), .Y(n_1569) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1527), .Y(n_1628) );
OAI21xp33_ASAP7_75t_SL g1529 ( .A1(n_1530), .A2(n_1535), .B(n_1536), .Y(n_1529) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
NAND2xp67_ASAP7_75t_L g1621 ( .A(n_1531), .B(n_1558), .Y(n_1621) );
NAND2xp5_ASAP7_75t_L g1641 ( .A(n_1531), .B(n_1603), .Y(n_1641) );
AND2x2_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1534), .Y(n_1531) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1532), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1616 ( .A(n_1532), .B(n_1561), .Y(n_1616) );
NAND2xp5_ASAP7_75t_L g1536 ( .A(n_1537), .B(n_1538), .Y(n_1536) );
CKINVDCx14_ASAP7_75t_R g1590 ( .A(n_1537), .Y(n_1590) );
NOR2xp33_ASAP7_75t_SL g1620 ( .A(n_1538), .B(n_1582), .Y(n_1620) );
NOR2xp33_ASAP7_75t_L g1538 ( .A(n_1539), .B(n_1540), .Y(n_1538) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1542), .Y(n_1638) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1545), .Y(n_1568) );
INVxp67_ASAP7_75t_SL g1546 ( .A(n_1547), .Y(n_1546) );
NOR2xp33_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1550), .Y(n_1547) );
OAI211xp5_ASAP7_75t_L g1567 ( .A1(n_1548), .A2(n_1568), .B(n_1569), .C(n_1573), .Y(n_1567) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1550), .Y(n_1572) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1553), .Y(n_1639) );
OAI211xp5_ASAP7_75t_L g1554 ( .A1(n_1555), .A2(n_1556), .B(n_1565), .C(n_1585), .Y(n_1554) );
AOI221xp5_ASAP7_75t_L g1606 ( .A1(n_1555), .A2(n_1558), .B1(n_1607), .B2(n_1615), .C(n_1617), .Y(n_1606) );
OAI22xp33_ASAP7_75t_SL g1617 ( .A1(n_1555), .A2(n_1618), .B1(n_1620), .B2(n_1621), .Y(n_1617) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
CKINVDCx5p33_ASAP7_75t_R g1583 ( .A(n_1584), .Y(n_1583) );
INVx1_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
OAI21xp33_ASAP7_75t_L g1589 ( .A1(n_1590), .A2(n_1591), .B(n_1592), .Y(n_1589) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
O2A1O1Ixp33_ASAP7_75t_L g1633 ( .A1(n_1595), .A2(n_1634), .B(n_1637), .C(n_1640), .Y(n_1633) );
A2O1A1Ixp33_ASAP7_75t_L g1596 ( .A1(n_1597), .A2(n_1598), .B(n_1605), .C(n_1606), .Y(n_1596) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1602), .Y(n_1601) );
INVx1_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1603), .B(n_1616), .Y(n_1615) );
INVx3_ASAP7_75t_L g1603 ( .A(n_1604), .Y(n_1603) );
OAI22xp5_ASAP7_75t_L g1607 ( .A1(n_1608), .A2(n_1610), .B1(n_1612), .B2(n_1614), .Y(n_1607) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1609), .Y(n_1608) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
A2O1A1Ixp33_ASAP7_75t_L g1622 ( .A1(n_1623), .A2(n_1630), .B(n_1631), .C(n_1633), .Y(n_1622) );
INVxp67_ASAP7_75t_SL g1623 ( .A(n_1624), .Y(n_1623) );
NOR2xp33_ASAP7_75t_L g1624 ( .A(n_1625), .B(n_1626), .Y(n_1624) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_1628), .B(n_1629), .Y(n_1627) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
INVxp67_ASAP7_75t_SL g1634 ( .A(n_1635), .Y(n_1634) );
NAND2xp5_ASAP7_75t_L g1637 ( .A(n_1638), .B(n_1639), .Y(n_1637) );
INVx2_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
BUFx2_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
NAND4xp75_ASAP7_75t_L g1648 ( .A(n_1649), .B(n_1650), .C(n_1670), .D(n_1683), .Y(n_1648) );
OAI31xp33_ASAP7_75t_L g1650 ( .A1(n_1651), .A2(n_1660), .A3(n_1668), .B(n_1669), .Y(n_1650) );
AND2x2_ASAP7_75t_SL g1670 ( .A(n_1671), .B(n_1682), .Y(n_1670) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
A2O1A1Ixp33_ASAP7_75t_L g1733 ( .A1(n_1681), .A2(n_1734), .B(n_1735), .C(n_1737), .Y(n_1733) );
CKINVDCx14_ASAP7_75t_R g1687 ( .A(n_1688), .Y(n_1687) );
INVx2_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
CKINVDCx5p33_ASAP7_75t_R g1689 ( .A(n_1690), .Y(n_1689) );
A2O1A1Ixp33_ASAP7_75t_L g1746 ( .A1(n_1691), .A2(n_1747), .B(n_1749), .C(n_1750), .Y(n_1746) );
CKINVDCx5p33_ASAP7_75t_R g1693 ( .A(n_1694), .Y(n_1693) );
INVx2_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
INVx1_ASAP7_75t_L g1699 ( .A(n_1700), .Y(n_1699) );
INVx2_ASAP7_75t_SL g1700 ( .A(n_1701), .Y(n_1700) );
INVx2_ASAP7_75t_L g1702 ( .A(n_1703), .Y(n_1702) );
NAND4xp75_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1719), .C(n_1738), .D(n_1741), .Y(n_1703) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1705), .B(n_1716), .Y(n_1704) );
INVx1_ASAP7_75t_SL g1706 ( .A(n_1707), .Y(n_1706) );
INVx2_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
NAND2xp5_ASAP7_75t_L g1720 ( .A(n_1721), .B(n_1724), .Y(n_1720) );
HB1xp67_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
endmodule