module fake_jpeg_29162_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

HAxp5_ASAP7_75t_SL g29 ( 
.A(n_14),
.B(n_0),
.CON(n_29),
.SN(n_29)
);

AND2x4_ASAP7_75t_SL g44 ( 
.A(n_29),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_32),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_18),
.B(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_22),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_13),
.B1(n_16),
.B2(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_23),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_19),
.B1(n_27),
.B2(n_20),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_44),
.B(n_49),
.C(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_23),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_35),
.C(n_27),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_20),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_63),
.B(n_53),
.Y(n_75)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_56),
.Y(n_77)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_66),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_45),
.C(n_40),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_19),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_26),
.B(n_25),
.C(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_18),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_28),
.B1(n_38),
.B2(n_31),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_58),
.B1(n_64),
.B2(n_57),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_82),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_76),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_19),
.B1(n_31),
.B2(n_25),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_31),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_90),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_56),
.C(n_52),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_93),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_67),
.B1(n_68),
.B2(n_0),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_76),
.B(n_1),
.Y(n_100)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_98),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_73),
.B(n_77),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_72),
.C(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_95),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_77),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_86),
.C(n_84),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_86),
.B1(n_87),
.B2(n_84),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_97),
.C(n_103),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_101),
.C(n_79),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_104),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_116),
.B(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_117),
.B(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_120),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_110),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_114),
.C(n_106),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_124),
.B(n_125),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_79),
.Y(n_125)
);

AOI21x1_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_7),
.B(n_8),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_12),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_126),
.B(n_12),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_129),
.B(n_71),
.CI(n_128),
.CON(n_130),
.SN(n_130)
);


endmodule