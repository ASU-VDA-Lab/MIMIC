module fake_jpeg_27587_n_197 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_197);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_30),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_6),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_14),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_39),
.B1(n_16),
.B2(n_18),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_16),
.B1(n_13),
.B2(n_19),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_48),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_20),
.B1(n_22),
.B2(n_16),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_28),
.A2(n_19),
.B1(n_21),
.B2(n_18),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_17),
.B1(n_25),
.B2(n_22),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_13),
.C(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_54),
.Y(n_74)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_57),
.Y(n_75)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_65),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_59),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_45),
.B1(n_51),
.B2(n_41),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_81),
.B1(n_84),
.B2(n_91),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_45),
.B(n_38),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_83),
.B(n_20),
.Y(n_101)
);

AND2x6_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_44),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_10),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_0),
.B(n_1),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_54),
.B1(n_50),
.B2(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_71),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_48),
.C(n_38),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_61),
.B1(n_37),
.B2(n_42),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_100),
.Y(n_116)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_97),
.Y(n_114)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_101),
.B(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_34),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_29),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_77),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_29),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_108),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_14),
.B1(n_27),
.B2(n_29),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_110),
.B(n_100),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_72),
.B1(n_80),
.B2(n_73),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_129),
.B1(n_106),
.B2(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_122),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_79),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_127),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_88),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_125),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_126),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_83),
.B(n_81),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_14),
.B(n_112),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_81),
.B1(n_89),
.B2(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_10),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_142),
.B1(n_124),
.B2(n_145),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_137),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_134),
.B(n_136),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_93),
.C(n_99),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_93),
.C(n_94),
.Y(n_137)
);

AOI321xp33_ASAP7_75t_L g157 ( 
.A1(n_138),
.A2(n_139),
.A3(n_146),
.B1(n_126),
.B2(n_130),
.C(n_118),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_98),
.B(n_106),
.C(n_112),
.D(n_96),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_145),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_92),
.B(n_89),
.Y(n_141)
);

AOI21x1_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_113),
.B(n_124),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_123),
.C(n_129),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_135),
.B(n_29),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_153),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_147),
.B(n_125),
.Y(n_153)
);

AO221x1_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_111),
.B1(n_97),
.B2(n_112),
.C(n_119),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_155),
.A2(n_157),
.B(n_158),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_122),
.B1(n_118),
.B2(n_116),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_165),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_136),
.C(n_137),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_148),
.A2(n_146),
.B(n_135),
.Y(n_164)
);

OAI21x1_ASAP7_75t_SL g175 ( 
.A1(n_164),
.A2(n_27),
.B(n_7),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_131),
.C(n_144),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_138),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_151),
.B(n_1),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_152),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_159),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_171),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_169),
.A2(n_150),
.B1(n_149),
.B2(n_156),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_175),
.B(n_11),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_2),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_176),
.Y(n_181)
);

NAND4xp25_ASAP7_75t_SL g176 ( 
.A(n_164),
.B(n_0),
.C(n_2),
.D(n_3),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_9),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_163),
.C(n_167),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_183),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_12),
.B(n_3),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_166),
.C(n_11),
.Y(n_183)
);

AOI31xp33_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_176),
.A3(n_171),
.B(n_173),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_11),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_179),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_187),
.B(n_189),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_181),
.C(n_183),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_184),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_3),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_193),
.B(n_191),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_4),
.B1(n_194),
.B2(n_188),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_4),
.Y(n_197)
);


endmodule