module fake_netlist_6_3927_n_782 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_782);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_782;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_153;
wire n_758;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_772;
wire n_656;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_683;
wire n_420;
wire n_620;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_164;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g148 ( 
.A(n_21),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_73),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_71),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_66),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_3),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_3),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_69),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_0),
.Y(n_157)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_102),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_34),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_52),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_59),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_20),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_64),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_4),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_83),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_62),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_24),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_85),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_126),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_37),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_33),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_57),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_72),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_100),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_94),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_81),
.Y(n_188)
);

BUFx2_ASAP7_75t_SL g189 ( 
.A(n_90),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_47),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_2),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_106),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_16),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_130),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_137),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_45),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_99),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_14),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_30),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_103),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_136),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_80),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_0),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_154),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_155),
.B(n_1),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_162),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_5),
.Y(n_215)
);

AND2x4_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_22),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_169),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_5),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_186),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_172),
.B(n_23),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_192),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_158),
.B(n_6),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_7),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

BUFx8_ASAP7_75t_SL g238 ( 
.A(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_185),
.Y(n_240)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_7),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

AND2x6_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_25),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_159),
.B(n_8),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_238),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_209),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_209),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_217),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_217),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_211),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_189),
.B(n_202),
.Y(n_263)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_176),
.B(n_197),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_R g265 ( 
.A(n_235),
.B(n_199),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_231),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_245),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_245),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_220),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_247),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_225),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_R g274 ( 
.A(n_235),
.B(n_199),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_225),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_225),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_225),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_233),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_205),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_233),
.Y(n_281)
);

BUFx6f_ASAP7_75t_SL g282 ( 
.A(n_216),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_235),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_241),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_241),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_220),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_241),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_220),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_241),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_210),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_210),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_213),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_210),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_216),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_216),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_268),
.B(n_227),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_227),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_212),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

BUFx6f_ASAP7_75t_SL g304 ( 
.A(n_251),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_270),
.B(n_227),
.Y(n_305)
);

AOI221xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_236),
.B1(n_234),
.B2(n_242),
.C(n_215),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_279),
.Y(n_307)
);

NAND2x1_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_244),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_280),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_205),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_286),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_283),
.B(n_246),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_274),
.B(n_222),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_218),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_222),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_222),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_273),
.B(n_161),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g321 ( 
.A(n_269),
.B(n_218),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_275),
.B(n_163),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_249),
.Y(n_325)
);

AND2x6_ASAP7_75t_SL g326 ( 
.A(n_267),
.B(n_207),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_262),
.B(n_239),
.C(n_226),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_290),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_243),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_249),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_206),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_277),
.B(n_164),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_264),
.B(n_166),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_252),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_249),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_289),
.B(n_243),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_291),
.B(n_243),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_263),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_282),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_282),
.B(n_230),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_253),
.B(n_230),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_255),
.B(n_221),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_259),
.B(n_221),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_261),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_281),
.B(n_151),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

NAND3xp33_ASAP7_75t_L g352 ( 
.A(n_248),
.B(n_214),
.C(n_206),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_250),
.B(n_221),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_286),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_254),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_292),
.B(n_221),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_268),
.B(n_230),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_254),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_292),
.B(n_228),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_268),
.B(n_167),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_268),
.B(n_230),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_249),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_333),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_244),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_321),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_307),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_307),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_192),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_316),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_309),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_303),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_170),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_346),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_302),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_244),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_347),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_310),
.B(n_345),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_306),
.A2(n_196),
.B1(n_150),
.B2(n_203),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_305),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_361),
.B(n_345),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_349),
.A2(n_150),
.B1(n_203),
.B2(n_175),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_244),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_174),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_297),
.B(n_177),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_244),
.Y(n_394)
);

O2A1O1Ixp5_ASAP7_75t_L g395 ( 
.A1(n_341),
.A2(n_229),
.B(n_244),
.C(n_228),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_330),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_298),
.B(n_179),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

AND2x4_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_181),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_362),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_299),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_335),
.A2(n_228),
.B1(n_232),
.B2(n_230),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_183),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_301),
.B(n_228),
.Y(n_405)
);

AOI21xp33_ASAP7_75t_L g406 ( 
.A1(n_299),
.A2(n_229),
.B(n_228),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_315),
.B(n_300),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

NOR2x1p5_ASAP7_75t_L g409 ( 
.A(n_348),
.B(n_352),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_344),
.B(n_187),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_312),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_322),
.Y(n_413)
);

NAND2x1p5_ASAP7_75t_L g414 ( 
.A(n_308),
.B(n_232),
.Y(n_414)
);

A2O1A1Ixp33_ASAP7_75t_L g415 ( 
.A1(n_344),
.A2(n_193),
.B(n_190),
.C(n_188),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_335),
.A2(n_237),
.B1(n_232),
.B2(n_10),
.Y(n_416)
);

NOR3xp33_ASAP7_75t_SL g417 ( 
.A(n_313),
.B(n_8),
.C(n_9),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_354),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_350),
.A2(n_304),
.B1(n_351),
.B2(n_331),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_315),
.B(n_232),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_313),
.A2(n_237),
.B1(n_232),
.B2(n_11),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_300),
.B(n_237),
.Y(n_424)
);

NOR2x2_ASAP7_75t_L g425 ( 
.A(n_326),
.B(n_9),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_325),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_325),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_328),
.Y(n_429)
);

INVx5_ASAP7_75t_L g430 ( 
.A(n_332),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_320),
.B(n_237),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_300),
.B(n_237),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_388),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_339),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_390),
.A2(n_404),
.B(n_372),
.C(n_402),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_375),
.B(n_378),
.Y(n_436)
);

AOI21x1_ASAP7_75t_L g437 ( 
.A1(n_420),
.A2(n_318),
.B(n_319),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_423),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_402),
.A2(n_340),
.B1(n_323),
.B2(n_334),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_395),
.A2(n_338),
.B(n_334),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_376),
.A2(n_323),
.B1(n_320),
.B2(n_300),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_364),
.B(n_342),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_373),
.Y(n_444)
);

AOI21xp33_ASAP7_75t_L g445 ( 
.A1(n_383),
.A2(n_10),
.B(n_11),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_407),
.A2(n_300),
.B(n_304),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_384),
.B(n_380),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_386),
.B(n_300),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_407),
.A2(n_86),
.B(n_147),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_SL g450 ( 
.A1(n_365),
.A2(n_377),
.B(n_389),
.C(n_394),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_366),
.B(n_12),
.Y(n_451)
);

NAND2x1p5_ASAP7_75t_L g452 ( 
.A(n_401),
.B(n_26),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_411),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_400),
.B(n_12),
.Y(n_454)
);

NOR3xp33_ASAP7_75t_SL g455 ( 
.A(n_387),
.B(n_13),
.C(n_14),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_383),
.B(n_13),
.Y(n_456)
);

AOI21x1_ASAP7_75t_L g457 ( 
.A1(n_420),
.A2(n_88),
.B(n_145),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_369),
.B(n_15),
.Y(n_458)
);

A2O1A1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_365),
.A2(n_377),
.B(n_389),
.C(n_363),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_400),
.B(n_15),
.Y(n_460)
);

INVx8_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

O2A1O1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_415),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_463)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_409),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_405),
.A2(n_91),
.B(n_140),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_368),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_419),
.B(n_27),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_410),
.B(n_374),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_385),
.B(n_17),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_422),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_391),
.B(n_19),
.Y(n_472)
);

OR2x6_ASAP7_75t_L g473 ( 
.A(n_379),
.B(n_28),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_370),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_393),
.B(n_29),
.Y(n_475)
);

BUFx12f_ASAP7_75t_L g476 ( 
.A(n_411),
.Y(n_476)
);

O2A1O1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_406),
.A2(n_31),
.B(n_32),
.C(n_35),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_401),
.A2(n_36),
.B(n_38),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_432),
.A2(n_39),
.B(n_40),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_R g480 ( 
.A(n_392),
.B(n_41),
.Y(n_480)
);

A2O1A1Ixp33_ASAP7_75t_L g481 ( 
.A1(n_396),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_397),
.B(n_46),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_431),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_399),
.B(n_51),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_408),
.B(n_53),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_412),
.B(n_54),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_398),
.B(n_55),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_418),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_371),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_416),
.A2(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_413),
.A2(n_61),
.B1(n_65),
.B2(n_67),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_476),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_444),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_462),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_443),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_457),
.A2(n_432),
.B(n_424),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_459),
.A2(n_424),
.B(n_414),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_446),
.A2(n_414),
.B(n_429),
.Y(n_498)
);

NAND2x1p5_ASAP7_75t_L g499 ( 
.A(n_485),
.B(n_421),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_437),
.A2(n_428),
.B(n_427),
.Y(n_500)
);

AO21x2_ASAP7_75t_L g501 ( 
.A1(n_450),
.A2(n_435),
.B(n_448),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_449),
.A2(n_426),
.B(n_403),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_438),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_461),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_461),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_441),
.A2(n_430),
.B(n_421),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_441),
.A2(n_430),
.B(n_421),
.Y(n_507)
);

AO21x2_ASAP7_75t_L g508 ( 
.A1(n_482),
.A2(n_406),
.B(n_417),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_467),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_464),
.B(n_430),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_474),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_452),
.A2(n_430),
.B(n_74),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_433),
.Y(n_513)
);

AOI22x1_ASAP7_75t_L g514 ( 
.A1(n_489),
.A2(n_425),
.B1(n_75),
.B2(n_76),
.Y(n_514)
);

AOI22x1_ASAP7_75t_L g515 ( 
.A1(n_439),
.A2(n_68),
.B1(n_77),
.B2(n_78),
.Y(n_515)
);

INVx8_ASAP7_75t_L g516 ( 
.A(n_461),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_466),
.Y(n_517)
);

INVx6_ASAP7_75t_L g518 ( 
.A(n_485),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_434),
.A2(n_79),
.B(n_82),
.Y(n_519)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_469),
.A2(n_84),
.B(n_87),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_452),
.A2(n_92),
.B(n_93),
.Y(n_521)
);

CKINVDCx6p67_ASAP7_75t_R g522 ( 
.A(n_473),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_473),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_473),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g525 ( 
.A(n_456),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_436),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_486),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

NAND2x1p5_ASAP7_75t_L g530 ( 
.A(n_486),
.B(n_95),
.Y(n_530)
);

INVx8_ASAP7_75t_L g531 ( 
.A(n_458),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_480),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_436),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_470),
.A2(n_96),
.B(n_97),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g535 ( 
.A1(n_440),
.A2(n_101),
.B(n_104),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_472),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_453),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_484),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_442),
.A2(n_105),
.B(n_107),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_478),
.A2(n_108),
.B(n_109),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_455),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_495),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_525),
.A2(n_468),
.B1(n_451),
.B2(n_445),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g544 ( 
.A1(n_532),
.A2(n_454),
.B1(n_460),
.B2(n_471),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_492),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_493),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_SL g547 ( 
.A1(n_525),
.A2(n_471),
.B1(n_490),
.B2(n_487),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_494),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_500),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_518),
.A2(n_447),
.B1(n_490),
.B2(n_475),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_517),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_528),
.B(n_481),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_516),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_500),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_503),
.Y(n_555)
);

OA21x2_ASAP7_75t_L g556 ( 
.A1(n_496),
.A2(n_465),
.B(n_479),
.Y(n_556)
);

OAI21x1_ASAP7_75t_SL g557 ( 
.A1(n_539),
.A2(n_463),
.B(n_477),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_506),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_506),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_509),
.Y(n_560)
);

BUFx2_ASAP7_75t_R g561 ( 
.A(n_492),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_SL g562 ( 
.A1(n_523),
.A2(n_445),
.B1(n_483),
.B2(n_491),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_507),
.A2(n_498),
.B(n_496),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_507),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_513),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_518),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_517),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_498),
.A2(n_497),
.B(n_512),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_524),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_516),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_533),
.Y(n_571)
);

NAND2x1_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_113),
.Y(n_572)
);

OA21x2_ASAP7_75t_L g573 ( 
.A1(n_502),
.A2(n_114),
.B(n_115),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_533),
.B(n_526),
.Y(n_574)
);

INVx8_ASAP7_75t_L g575 ( 
.A(n_516),
.Y(n_575)
);

AOI21x1_ASAP7_75t_L g576 ( 
.A1(n_502),
.A2(n_116),
.B(n_117),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_511),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_533),
.Y(n_578)
);

CKINVDCx11_ASAP7_75t_R g579 ( 
.A(n_524),
.Y(n_579)
);

AO21x2_ASAP7_75t_L g580 ( 
.A1(n_501),
.A2(n_119),
.B(n_120),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_536),
.A2(n_518),
.B1(n_528),
.B2(n_531),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_526),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_SL g583 ( 
.A(n_547),
.B(n_543),
.C(n_562),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_542),
.B(n_536),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_567),
.B(n_529),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_548),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_551),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_SL g588 ( 
.A(n_569),
.B(n_541),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_567),
.B(n_522),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_546),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_546),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_544),
.B(n_531),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_555),
.B(n_522),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_571),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_555),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_582),
.B(n_565),
.Y(n_596)
);

OAI211xp5_ASAP7_75t_L g597 ( 
.A1(n_550),
.A2(n_514),
.B(n_519),
.C(n_541),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_569),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_582),
.B(n_508),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_560),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_574),
.B(n_523),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_577),
.B(n_508),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_570),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_577),
.B(n_531),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_552),
.A2(n_531),
.B1(n_538),
.B2(n_530),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_510),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_R g607 ( 
.A(n_552),
.B(n_534),
.Y(n_607)
);

BUFx8_ASAP7_75t_L g608 ( 
.A(n_570),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_545),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_570),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_575),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_561),
.Y(n_612)
);

NAND2xp33_ASAP7_75t_SL g613 ( 
.A(n_570),
.B(n_504),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_R g614 ( 
.A(n_552),
.B(n_534),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_R g615 ( 
.A(n_545),
.B(n_516),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_579),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_578),
.A2(n_499),
.B1(n_530),
.B2(n_537),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_578),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_572),
.Y(n_619)
);

BUFx4f_ASAP7_75t_L g620 ( 
.A(n_570),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_572),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_553),
.A2(n_499),
.B1(n_510),
.B2(n_505),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_R g623 ( 
.A(n_575),
.B(n_505),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_553),
.B(n_510),
.Y(n_624)
);

OA21x2_ASAP7_75t_L g625 ( 
.A1(n_568),
.A2(n_540),
.B(n_512),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_SL g626 ( 
.A1(n_557),
.A2(n_535),
.B1(n_515),
.B2(n_534),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_553),
.A2(n_527),
.B1(n_504),
.B2(n_520),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_549),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_557),
.A2(n_535),
.B1(n_566),
.B2(n_580),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_628),
.B(n_535),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_599),
.B(n_501),
.Y(n_631)
);

NOR4xp25_ASAP7_75t_SL g632 ( 
.A(n_607),
.B(n_580),
.C(n_576),
.D(n_521),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_591),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_602),
.B(n_501),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_590),
.B(n_580),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_594),
.B(n_554),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_600),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_584),
.B(n_521),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_594),
.B(n_554),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_586),
.B(n_549),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_595),
.Y(n_641)
);

NAND4xp25_ASAP7_75t_L g642 ( 
.A(n_601),
.B(n_564),
.C(n_559),
.D(n_558),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_625),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_619),
.B(n_564),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_625),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_621),
.B(n_559),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_618),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_596),
.B(n_573),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_601),
.B(n_558),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_583),
.B(n_568),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_583),
.B(n_563),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_592),
.A2(n_540),
.B1(n_575),
.B2(n_556),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_608),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_606),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_605),
.B(n_563),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_604),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_593),
.B(n_556),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_585),
.B(n_576),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_609),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_629),
.B(n_556),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_587),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_629),
.B(n_556),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_627),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_617),
.B(n_575),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_624),
.B(n_121),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_656),
.B(n_589),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_637),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_SL g668 ( 
.A1(n_654),
.A2(n_597),
.B1(n_615),
.B2(n_623),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_633),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_633),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_641),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_641),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_657),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_640),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_634),
.B(n_626),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_634),
.B(n_626),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_656),
.B(n_597),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_656),
.B(n_603),
.Y(n_678)
);

AND2x4_ASAP7_75t_SL g679 ( 
.A(n_649),
.B(n_603),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_640),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_631),
.B(n_603),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_631),
.B(n_603),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_654),
.B(n_610),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_636),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_643),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_636),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_657),
.B(n_588),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_639),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_649),
.B(n_610),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_637),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_675),
.B(n_660),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_689),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_675),
.B(n_660),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_676),
.B(n_662),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_676),
.B(n_662),
.Y(n_695)
);

NAND4xp25_ASAP7_75t_L g696 ( 
.A(n_677),
.B(n_666),
.C(n_659),
.D(n_668),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_681),
.B(n_655),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_673),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_667),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_681),
.B(n_655),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_690),
.B(n_659),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_673),
.B(n_650),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_671),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_671),
.Y(n_704)
);

BUFx2_ASAP7_75t_L g705 ( 
.A(n_682),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_669),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_692),
.B(n_687),
.Y(n_707)
);

OAI22xp33_ASAP7_75t_L g708 ( 
.A1(n_696),
.A2(n_650),
.B1(n_614),
.B2(n_607),
.Y(n_708)
);

OAI322xp33_ASAP7_75t_L g709 ( 
.A1(n_702),
.A2(n_688),
.A3(n_680),
.B1(n_674),
.B2(n_670),
.C1(n_672),
.C2(n_684),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_699),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_SL g711 ( 
.A1(n_691),
.A2(n_653),
.B1(n_683),
.B2(n_651),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_698),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_698),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_703),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_705),
.B(n_682),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_702),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_691),
.A2(n_642),
.B1(n_655),
.B2(n_613),
.Y(n_717)
);

OAI222xp33_ASAP7_75t_L g718 ( 
.A1(n_693),
.A2(n_687),
.B1(n_651),
.B2(n_683),
.C1(n_638),
.C2(n_686),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_708),
.A2(n_701),
.B(n_699),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_708),
.A2(n_694),
.B1(n_693),
.B2(n_695),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_714),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_714),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_717),
.A2(n_695),
.B1(n_694),
.B2(n_655),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_722),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_719),
.A2(n_718),
.B(n_709),
.Y(n_725)
);

O2A1O1Ixp5_ASAP7_75t_L g726 ( 
.A1(n_721),
.A2(n_707),
.B(n_710),
.C(n_713),
.Y(n_726)
);

AOI222xp33_ASAP7_75t_L g727 ( 
.A1(n_720),
.A2(n_661),
.B1(n_716),
.B2(n_712),
.C1(n_706),
.C2(n_705),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_724),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_726),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_725),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_728),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_SL g732 ( 
.A(n_730),
.B(n_727),
.C(n_723),
.Y(n_732)
);

AOI31xp33_ASAP7_75t_L g733 ( 
.A1(n_732),
.A2(n_612),
.A3(n_729),
.B(n_616),
.Y(n_733)
);

OAI211xp5_ASAP7_75t_L g734 ( 
.A1(n_731),
.A2(n_711),
.B(n_615),
.C(n_653),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_731),
.B(n_716),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_734),
.A2(n_653),
.B1(n_598),
.B2(n_678),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_735),
.Y(n_737)
);

NOR2x1_ASAP7_75t_L g738 ( 
.A(n_733),
.B(n_598),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_735),
.B(n_715),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_734),
.A2(n_700),
.B1(n_697),
.B2(n_665),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_735),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_738),
.A2(n_704),
.B1(n_620),
.B2(n_697),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_737),
.B(n_700),
.Y(n_743)
);

AND3x2_ASAP7_75t_L g744 ( 
.A(n_741),
.B(n_665),
.C(n_623),
.Y(n_744)
);

AOI221xp5_ASAP7_75t_L g745 ( 
.A1(n_739),
.A2(n_663),
.B1(n_652),
.B2(n_658),
.C(n_622),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_736),
.A2(n_614),
.B1(n_658),
.B2(n_679),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_740),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_744),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_747),
.B(n_679),
.Y(n_749)
);

XNOR2xp5_ASAP7_75t_L g750 ( 
.A(n_742),
.B(n_611),
.Y(n_750)
);

NAND4xp25_ASAP7_75t_L g751 ( 
.A(n_743),
.B(n_746),
.C(n_745),
.D(n_611),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_747),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_743),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_747),
.A2(n_620),
.B1(n_608),
.B2(n_610),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_748),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_753),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_752),
.Y(n_757)
);

OA22x2_ASAP7_75t_L g758 ( 
.A1(n_754),
.A2(n_663),
.B1(n_685),
.B2(n_688),
.Y(n_758)
);

OA22x2_ASAP7_75t_L g759 ( 
.A1(n_750),
.A2(n_663),
.B1(n_685),
.B2(n_647),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_749),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_751),
.A2(n_610),
.B1(n_630),
.B2(n_648),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_752),
.B(n_122),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_752),
.B(n_123),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_760),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_755),
.A2(n_664),
.B1(n_647),
.B2(n_643),
.Y(n_765)
);

AOI211xp5_ASAP7_75t_L g766 ( 
.A1(n_757),
.A2(n_664),
.B(n_630),
.C(n_648),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_759),
.Y(n_767)
);

XNOR2xp5_ASAP7_75t_L g768 ( 
.A(n_762),
.B(n_124),
.Y(n_768)
);

OAI31xp33_ASAP7_75t_L g769 ( 
.A1(n_756),
.A2(n_630),
.A3(n_635),
.B(n_646),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_763),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_758),
.Y(n_771)
);

OAI21x1_ASAP7_75t_L g772 ( 
.A1(n_764),
.A2(n_761),
.B(n_647),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_771),
.A2(n_632),
.B1(n_630),
.B2(n_645),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_SL g774 ( 
.A(n_767),
.B(n_125),
.C(n_127),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_768),
.A2(n_643),
.B1(n_645),
.B2(n_646),
.Y(n_775)
);

OAI21x1_ASAP7_75t_SL g776 ( 
.A1(n_770),
.A2(n_128),
.B(n_129),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_776),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_774),
.A2(n_770),
.B1(n_765),
.B2(n_766),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_777),
.A2(n_775),
.B1(n_773),
.B2(n_772),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_SL g780 ( 
.A1(n_779),
.A2(n_778),
.B1(n_769),
.B2(n_635),
.Y(n_780)
);

AOI221xp5_ASAP7_75t_L g781 ( 
.A1(n_780),
.A2(n_644),
.B1(n_646),
.B2(n_133),
.C(n_135),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_781),
.A2(n_646),
.B1(n_644),
.B2(n_645),
.Y(n_782)
);


endmodule