module fake_jpeg_5368_n_96 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_62;
wire n_43;
wire n_82;

INVx6_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_0),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_62),
.B(n_50),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_1),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_51),
.B1(n_39),
.B2(n_45),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_67),
.B1(n_55),
.B2(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_1),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_56),
.B1(n_51),
.B2(n_54),
.Y(n_67)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_72),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_47),
.B1(n_46),
.B2(n_64),
.Y(n_74)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_73),
.B(n_3),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_63),
.C(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_44),
.B1(n_40),
.B2(n_6),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_71),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_8),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_75),
.B1(n_10),
.B2(n_13),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_80),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_86),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_83),
.B1(n_81),
.B2(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_9),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_18),
.B(n_22),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_23),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_92),
.B(n_25),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_26),
.B(n_29),
.C(n_30),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_31),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_33),
.Y(n_96)
);


endmodule